module wa( IZZ,
 IAA, 
 IAB, 
 IAC, 
 IAD, 
 IAE, 
 IAF, 
 IAG, 
 IAH, 
 IAI, 
 IAJ, 
 IAK, 
 IAL, 
 IAM, 
 IAN, 
 IAO, 
 IAP, 
 IBA, 
 IBB, 
 IBC, 
 IBD, 
 IBE, 
 IBF, 
 IBG, 
 IBH, 
 IBI, 
 IBJ, 
 IBK, 
 IBL, 
 IBM, 
 IBN, 
 IBO, 
 IBP, 
 ICA, 
 ICB, 
 ICC, 
 ICD, 
 ICE, 
 ICF, 
 ICG, 
 ICH, 
 ICI, 
 ICJ, 
 ICK, 
 ICL, 
 ICM, 
 ICN, 
 ICO, 
 ICP, 
 IDA, 
 IDB, 
 IDC, 
 IDD, 
 IDE, 
 IDF, 
 IDG, 
 IDH, 
 IDI, 
 IDJ, 
 IDK, 
 IDL, 
 IDM, 
 IDN, 
 IDO, 
 IDP, 
 IEA, 
 IEB, 
 IEC, 
 IED, 
 IEE, 
 IEF, 
 IEG, 
 IEH, 
 IEI, 
 IEJ, 
 IEK, 
 IEL, 
 IEM, 
 IEN, 
 IEO, 
 IEP, 
 IFA, 
 IFB, 
 IFC, 
 IFD, 
 IFE, 
 IFFF , 
 IFG, 
 IFH, 
 IFI, 
 IFJ, 
 IFK, 
 IFL, 
 IFM, 
 IFN, 
 IFO, 
 IFP, 
 IGA, 
 IGB, 
 IGC, 
 IGD, 
 IGE, 
 IGF, 
 IGG, 
 IGH, 
 IGI, 
 IGJ, 
 IGK, 
 IGL, 
 IGM, 
 IGN, 
 IGO, 
 IGP, 
 IHA, 
 IHB, 
 IIA, 
 IIB, 
 IJA, 
 IJB, 
 IJC, 
 IJD, 
 OAA, 
 OAB, 
 OAC, 
 OAD, 
 OAE, 
 OAF, 
 OAG, 
 OAH, 
 OAI, 
 OAJ, 
 OAK, 
 OAL, 
 OAM, 
 OAN, 
 OAO, 
 OAP, 
 OBA, 
 OBB, 
 OBC, 
 OBD, 
 OBE, 
 OBF, 
 OBG, 
 OBH, 
 OBI, 
 OBJ, 
 OBK, 
 OBL, 
 OBM, 
 OBN, 
 OBO, 
 OBP, 
 OCA, 
 OCB, 
 OCC, 
 OCD, 
 OCE, 
 OCF, 
 OCG, 
 OCH, 
 OCI, 
 OCJ, 
 OCK, 
 OCL, 
 OCM, 
 OCN, 
 OCO, 
 OCP, 
 ODA, 
 ODB, 
 ODC, 
 ODD, 
 ODE, 
 ODF, 
 ODG, 
 ODH, 
 ODI, 
 ODJ, 
 ODK, 
 ODL, 
 ODM, 
 ODN, 
 ODO, 
 ODP, 
 OEA, 
 OEB, 
 OEC, 
 OED, 
 OEE, 
 OEF, 
 OEG, 
 OEH, 
 OEI, 
 OEJ, 
 OEK, 
 OEL, 
 OEM, 
 OEN, 
 OEO, 
 OEP, 
 OFA, 
 OFB, 
 OFC, 
 OFD, 
 OFE, 
 OFF, 
 OFG, 
 OFH, 
 OFI, 
 OFJ, 
 OFK, 
 OFL, 
 OFM, 
 OFN, 
 OFO, 
OFP ); 
    
 input IZZ; 
 input IAA; 
 input IAB; 
 input IAC; 
 input IAD; 
 input IAE; 
 input IAF; 
 input IAG; 
 input IAH; 
 input IAI; 
 input IAJ; 
 input IAK; 
 input IAL; 
 input IAM; 
 input IAN; 
 input IAO; 
 input IAP; 
 input IBA; 
 input IBB; 
 input IBC; 
 input IBD; 
 input IBE; 
 input IBF; 
 input IBG; 
 input IBH; 
 input IBI; 
 input IBJ; 
 input IBK; 
 input IBL; 
 input IBM; 
 input IBN; 
 input IBO; 
 input IBP; 
 input ICA; 
 input ICB; 
 input ICC; 
 input ICD; 
 input ICE; 
 input ICF; 
 input ICG; 
 input ICH; 
 input ICI; 
 input ICJ; 
 input ICK; 
 input ICL; 
 input ICM; 
 input ICN; 
 input ICO; 
 input ICP; 
 input IDA; 
 input IDB; 
 input IDC; 
 input IDD; 
 input IDE; 
 input IDF; 
 input IDG; 
 input IDH; 
 input IDI; 
 input IDJ; 
 input IDK; 
 input IDL; 
 input IDM; 
 input IDN; 
 input IDO; 
 input IDP; 
 input IEA; 
 input IEB; 
 input IEC; 
 input IED; 
 input IEE; 
 input IEF; 
 input IEG; 
 input IEH; 
 input IEI; 
 input IEJ; 
 input IEK; 
 input IEL; 
 input IEM; 
 input IEN; 
 input IEO; 
 input IEP; 
 input IFA; 
 input IFB; 
 input IFC; 
 input IFD; 
 input IFE; 
 input IFFF ; 
 input IFG; 
 input IFH; 
 input IFI; 
 input IFJ; 
 input IFK; 
 input IFL; 
 input IFM; 
 input IFN; 
 input IFO; 
 input IFP; 
 input IGA; 
 input IGB; 
 input IGC; 
 input IGD; 
 input IGE; 
 input IGF; 
 input IGG; 
 input IGH; 
 input IGI; 
 input IGJ; 
 input IGK; 
 input IGL; 
 input IGM; 
 input IGN; 
 input IGO; 
 input IGP; 
 input IHA; 
 input IHB; 
 input IIA; 
 input IIB; 
 input IJA; 
 input IJB; 
 input IJC; 
 input IJD; 
 output OAA; 
 output OAB; 
 output OAC; 
 output OAD; 
 output OAE; 
 output OAF; 
 output OAG; 
 output OAH; 
 output OAI; 
 output OAJ; 
 output OAK; 
 output OAL; 
 output OAM; 
 output OAN; 
 output OAO; 
 output OAP; 
 output OBA; 
 output OBB; 
 output OBC; 
 output OBD; 
 output OBE; 
 output OBF; 
 output OBG; 
 output OBH; 
 output OBI; 
 output OBJ; 
 output OBK; 
 output OBL; 
 output OBM; 
 output OBN; 
 output OBO; 
 output OBP; 
 output OCA; 
 output OCB; 
 output OCC; 
 output OCD; 
 output OCE; 
 output OCF; 
 output OCG; 
 output OCH; 
 output OCI; 
 output OCJ; 
 output OCK; 
 output OCL; 
 output OCM; 
 output OCN; 
 output OCO; 
 output OCP; 
 output ODA; 
 output ODB; 
 output ODC; 
 output ODD; 
 output ODE; 
 output ODF; 
 output ODG; 
 output ODH; 
 output ODI; 
 output ODJ; 
 output ODK; 
 output ODL; 
 output ODM; 
 output ODN; 
 output ODO; 
 output ODP; 
 output OEA; 
 output OEB; 
 output OEC; 
 output OED; 
 output OEE; 
 output OEF; 
 output OEG; 
 output OEH; 
 output OEI; 
 output OEJ; 
 output OEK; 
 output OEL; 
 output OEM; 
 output OEN; 
 output OEO; 
 output OEP; 
 output OFA; 
 output OFB; 
 output OFC; 
 output OFD; 
 output OFE; 
 output OFF; 
 output OFG; 
 output OFH; 
 output OFI; 
 output OFJ; 
 output OFK; 
 output OFL; 
 output OFM; 
 output OFN; 
 output OFO; 
 output OFP; 
  
  
reg  AAA ;
reg  AAB ;
reg  AAC ;
reg  AAD ;
reg  AAE ;
reg  AAF ;
reg  AAG ;
reg  AAH ;
reg  AAI ;
reg  AAJ ;
reg  AAK ;
reg  AAL ;
reg  ABA ;
reg  ABB ;
reg  ABC ;
reg  ABD ;
reg  ABE ;
reg  ABF ;
reg  ABG ;
reg  ABH ;
reg  ABI ;
reg  ABJ ;
reg  ABK ;
reg  ABL ;
reg  ACA ;
reg  ACB ;
reg  ACC ;
reg  ACD ;
reg  ACE ;
reg  ACF ;
reg  ACG ;
reg  ACH ;
reg  ACI ;
reg  ACJ ;
reg  ACK ;
reg  ACL ;
reg  ADA ;
reg  ADB ;
reg  ADC ;
reg  ADD ;
reg  ADE ;
reg  ADF ;
reg  ADG ;
reg  ADH ;
reg  ADI ;
reg  ADJ ;
reg  ADK ;
reg  ADL ;
reg  AEA ;
reg  AEB ;
reg  AEC ;
reg  AED ;
reg  AEE ;
reg  AEF ;
reg  AEG ;
reg  AEH ;
reg  AEI ;
reg  AEJ ;
reg  AEK ;
reg  AEL ;
reg  AFA ;
reg  AFB ;
reg  AFC ;
reg  AFD ;
reg  AFE ;
reg  AFF ;
reg  AFG ;
reg  AFH ;
reg  AFI ;
reg  AFJ ;
reg  AFK ;
reg  AFL ;
reg  AGA ;
reg  AGB ;
reg  AGC ;
reg  AGD ;
reg  AGE ;
reg  AGF ;
reg  AGG ;
reg  AGH ;
reg  AGI ;
reg  AGJ ;
reg  AGK ;
reg  AGL ;
reg  AHA ;
reg  AHB ;
reg  AHC ;
reg  AHD ;
reg  AHE ;
reg  AHF ;
reg  AHG ;
reg  AHH ;
reg  AHI ;
reg  AHJ ;
reg  AHK ;
reg  AHL ;
reg  BAA ;
reg  BAB ;
reg  BAC ;
reg  BAD ;
reg  BAE ;
reg  BAF ;
reg  BAG ;
reg  BAH ;
reg  BAI ;
reg  BAJ ;
reg  BAK ;
reg  BAL ;
reg  BAM ;
reg  BAN ;
reg  BAO ;
reg  BAP ;
reg  BBA ;
reg  BBB ;
reg  BBC ;
reg  BBD ;
reg  BBE ;
reg  BBF ;
reg  BBG ;
reg  BBH ;
reg  BBI ;
reg  BBJ ;
reg  BBK ;
reg  BBL ;
reg  BBM ;
reg  BBN ;
reg  BBO ;
reg  BBP ;
reg  BCA ;
reg  BCB ;
reg  BCC ;
reg  BCD ;
reg  BCE ;
reg  BCF ;
reg  BCG ;
reg  BCH ;
reg  BCI ;
reg  BCJ ;
reg  BCK ;
reg  BCL ;
reg  BCM ;
reg  BCN ;
reg  BCO ;
reg  BCP ;
reg  BDA ;
reg  BDB ;
reg  BDC ;
reg  BDD ;
reg  BDE ;
reg  BDF ;
reg  BDG ;
reg  BDH ;
reg  BDI ;
reg  BDJ ;
reg  BDK ;
reg  BDL ;
reg  BDM ;
reg  BDN ;
reg  BDO ;
reg  BDP ;
reg  BEA ;
reg  BEB ;
reg  BEC ;
reg  BED ;
reg  BEE ;
reg  BEF ;
reg  BEG ;
reg  BEH ;
reg  BEI ;
reg  BEJ ;
reg  BEK ;
reg  BEL ;
reg  BEM ;
reg  BEN ;
reg  BEO ;
reg  BEP ;
reg  BFA ;
reg  BFB ;
reg  BFC ;
reg  BFD ;
reg  BFE ;
reg  BFF ;
reg  BFG ;
reg  BFH ;
reg  BFI ;
reg  BFJ ;
reg  BFK ;
reg  BFL ;
reg  BFM ;
reg  BFN ;
reg  BFO ;
reg  BFP ;
reg  BGA ;
reg  BGB ;
reg  BGC ;
reg  BGD ;
reg  BGE ;
reg  BGF ;
reg  BGG ;
reg  BGH ;
reg  BGI ;
reg  BGJ ;
reg  BGK ;
reg  BGL ;
reg  BGM ;
reg  BGN ;
reg  BGO ;
reg  BGP ;
reg  BHA ;
reg  BHB ;
reg  BHC ;
reg  BHD ;
reg  BHE ;
reg  BHF ;
reg  BHG ;
reg  BHH ;
reg  BHI ;
reg  BHJ ;
reg  BHK ;
reg  BHL ;
reg  BHM ;
reg  BHN ;
reg  BHO ;
reg  BHP ;
reg  FAA ;
reg  FAB ;
reg  FAC ;
reg  FAD ;
reg  FAE ;
reg  FAF ;
reg  FAG ;
reg  FAH ;
reg  FAI ;
reg  FAJ ;
reg  FAK ;
reg  FAL ;
reg  FBA ;
reg  FBB ;
reg  FBC ;
reg  FBD ;
reg  FBE ;
reg  FBF ;
reg  FBG ;
reg  FBH ;
reg  FBI ;
reg  FBJ ;
reg  FBK ;
reg  FBL ;
reg  GAA ;
reg  GAB ;
reg  GAC ;
reg  GAD ;
reg  GAE ;
reg  GAF ;
reg  GAG ;
reg  GAH ;
reg  GAI ;
reg  GAJ ;
reg  GAK ;
reg  GAL ;
reg  JMA ;
reg  JMB ;
reg  JMC ;
reg  JMD ;
reg  JME ;
reg  JMF ;
reg  JMG ;
reg  JMH ;
reg  KAA ;
reg  KAB ;
reg  KAC ;
reg  KAD ;
reg  KAE ;
reg  KAF ;
reg  KAG ;
reg  KAH ;
reg  KAI ;
reg  KAJ ;
reg  KAK ;
reg  KAL ;
reg  KAM ;
reg  KAN ;
reg  KAO ;
reg  KAP ;
reg  MAA ;
reg  MAB ;
reg  MAC ;
reg  MAD ;
reg  MAE ;
reg  MAF ;
reg  MAG ;
reg  MAH ;
reg  MAI ;
reg  MAJ ;
reg  MAK ;
reg  MAL ;
reg  MAM ;
reg  MAN ;
reg  MAO ;
reg  MAP ;
reg  MAQ ;
reg  MAR ;
reg  MAS ;
reg  MAT ;
reg  MAU ;
reg  MAV ;
reg  MAW ;
reg  MAX ;
reg  NAA ;
reg  NAB ;
reg  NAC ;
reg  NAD ;
reg  NAE ;
reg  NAF ;
reg  NAG ;
reg  NAH ;
reg  NAI ;
reg  NAJ ;
reg  NAK ;
reg  NAL ;
reg  NAM ;
reg  NAN ;
reg  NAO ;
reg  NAP ;
reg  NBA ;
reg  NBB ;
reg  NBC ;
reg  NBD ;
reg  NBE ;
reg  NBF ;
reg  NBG ;
reg  NBH ;
reg  NBI ;
reg  NBJ ;
reg  NBK ;
reg  NBL ;
reg  NBM ;
reg  NBN ;
reg  NBO ;
reg  NBP ;
reg  NCA ;
reg  NCB ;
reg  NCC ;
reg  NCD ;
reg  NCE ;
reg  NCF ;
reg  NCG ;
reg  NCH ;
reg  nci ;
reg  ncj ;
reg  nck ;
reg  ncl ;
reg  ncm ;
reg  ncn ;
reg  nco ;
reg  ncp ;
reg  NDA ;
reg  NDB ;
reg  NDC ;
reg  NDD ;
reg  NDE ;
reg  NDF ;
reg  NDG ;
reg  NDH ;
reg  ndi ;
reg  ndj ;
reg  ndk ;
reg  ndl ;
reg  ndm ;
reg  ndn ;
reg  ndo ;
reg  ndp ;
reg  OAA ;
reg  OAB ;
reg  OAC ;
reg  OAD ;
reg  OAE ;
reg  OAF ;
reg  OAG ;
reg  OAH ;
reg  OAI ;
reg  OAJ ;
reg  OAK ;
reg  OAL ;
reg  OAM ;
reg  OAN ;
reg  OAO ;
reg  OAP ;
reg  OBA ;
reg  OBB ;
reg  OBC ;
reg  OBD ;
reg  OBE ;
reg  OBF ;
reg  OBG ;
reg  OBH ;
reg  OBI ;
reg  OBJ ;
reg  OBK ;
reg  OBL ;
reg  OBM ;
reg  OBN ;
reg  OBO ;
reg  OBP ;
reg  OCA ;
reg  OCB ;
reg  OCC ;
reg  OCD ;
reg  OCE ;
reg  OCF ;
reg  OCG ;
reg  OCH ;
reg  OCI ;
reg  OCJ ;
reg  OCK ;
reg  OCL ;
reg  OCM ;
reg  OCN ;
reg  OCO ;
reg  OCP ;
reg  ODA ;
reg  ODB ;
reg  ODC ;
reg  ODD ;
reg  ODE ;
reg  ODF ;
reg  ODG ;
reg  ODH ;
reg  ODI ;
reg  ODJ ;
reg  ODK ;
reg  ODL ;
reg  ODM ;
reg  ODN ;
reg  ODO ;
reg  ODP ;
reg  OEA ;
reg  OEB ;
reg  OEC ;
reg  OED ;
reg  OEE ;
reg  OEF ;
reg  OEG ;
reg  OEH ;
reg  OEI ;
reg  OEJ ;
reg  OEK ;
reg  OEL ;
reg  OEM ;
reg  OEN ;
reg  OEO ;
reg  OEP ;
reg  OFA ;
reg  OFB ;
reg  OFC ;
reg  OFD ;
reg  OFE ;
reg  OFF ;
reg  OFG ;
reg  OFH ;
reg  OFI ;
reg  OFJ ;
reg  OFK ;
reg  OFL ;
reg  OFM ;
reg  OFN ;
reg  OFO ;
reg  OFP ;
reg  OHA ;
reg  OHB ;
reg  OHC ;
reg  OHD ;
reg  OHE ;
reg  OHF ;
reg  OHG ;
reg  OHH ;
reg  PAA ;
reg  PAB ;
reg  PAC ;
reg  PAD ;
reg  PBA ;
reg  PBB ;
reg  PBC ;
reg  PBD ;
reg  PCA ;
reg  PCB ;
reg  PCC ;
reg  PCD ;
reg  PCE ;
reg  PCF ;
reg  PCG ;
reg  PCH ;
reg  PDA ;
reg  PDB ;
reg  PDC ;
reg  PDD ;
reg  PEA ;
reg  PEB ;
reg  PEC ;
reg  PED ;
reg  QAA ;
reg  QAB ;
reg  QAC ;
reg  QBB ;
reg  QBC ;
reg  QBD ;
reg  QDA ;
reg  QDB ;
reg  QDC ;
reg  QFA ;
reg  TEA ;
reg  TEB ;
reg  TEC ;
reg  TED ;
reg  TEE ;
reg  TEF ;
reg  TEG ;
reg  TEH ;
reg  TEI ;
reg  TEJ ;
reg  tek ;
reg  tel ;
reg  tem ;
reg  ten ;
reg  teo ;
reg  tep ;
reg  teq ;
reg  ter ;
reg  TFA ;
reg  TFB ;
reg  TFC ;
reg  TFD ;
reg  TFE ;
reg  TFF ;
reg  TFG ;
reg  TFH ;
reg  TFI ;
reg  TFJ ;
reg  tfk ;
reg  tfl ;
reg  tfm ;
reg  tfn ;
reg  tfo ;
reg  tfp ;
reg  tfq ;
reg  tfr ;
reg  TGA ;
reg  TGB ;
reg  TGC ;
reg  TGD ;
reg  TGE ;
reg  TGF ;
reg  TGG ;
reg  TGH ;
reg  TGI ;
reg  TGJ ;
reg  tgk ;
reg  tgl ;
reg  tgm ;
reg  tgn ;
reg  tgo ;
reg  tgp ;
reg  tgq ;
reg  tgr ;
reg  THA ;
reg  THB ;
reg  THC ;
reg  THD ;
reg  THE ;
reg  THF ;
reg  THG ;
reg  THH ;
reg  THI ;
reg  THJ ;
reg  thk ;
reg  thl ;
reg  thm ;
reg  thn ;
reg  tho ;
reg  thp ;
reg  thq ;
reg  thr ;
reg  TMA ;
reg  TMB ;
reg  TMC ;
reg  TMD ;
reg  TME ;
reg  TMF ;
reg  TMG ;
reg  TMH ;
reg  TUA ;
reg  TUB ;
reg  TUC ;
reg  TUD ;
reg  TUE ;
reg  TUF ;
reg  TUG ;
reg  TUH ;
reg  TUI ;
reg  TUJ ;
reg  tuk ;
reg  tul ;
reg  tum ;
reg  tun ;
reg  tuo ;
reg  tup ;
reg  tuq ;
reg  tur ;
reg  TVA ;
reg  TVB ;
reg  TVC ;
reg  TVD ;
reg  TVE ;
reg  TVF ;
reg  TVG ;
reg  TVH ;
reg  TVI ;
reg  TVJ ;
reg  tvk ;
reg  tvl ;
reg  tvm ;
reg  tvn ;
reg  tvo ;
reg  tvp ;
reg  tvq ;
reg  tvr ;
reg  TWA ;
reg  TWB ;
reg  TWC ;
reg  TWD ;
reg  TWE ;
reg  TWF ;
reg  TWG ;
reg  TWH ;
reg  TWI ;
reg  TWJ ;
reg  twk ;
reg  twl ;
reg  twm ;
reg  twn ;
reg  two ;
reg  twp ;
reg  twq ;
reg  twr ;
reg  TXA ;
reg  TXB ;
reg  TXC ;
reg  TXD ;
reg  TXE ;
reg  TXF ;
reg  TXG ;
reg  TXH ;
reg  TXI ;
reg  TXJ ;
reg  txk ;
reg  txl ;
reg  txm ;
reg  txn ;
reg  txo ;
reg  txp ;
reg  txq ;
reg  txr ;
reg  WAA ;
reg  WAB ;
reg  WAC ;
reg  WAD ;
reg  WAE ;
reg  WAF ;
reg  WAG ;
reg  WAH ;
reg  wai ;
reg  waj ;
reg  wak ;
reg  wal ;
reg  wam ;
reg  wan ;
reg  wao ;
reg  wap ;
reg  WBA ;
reg  WBB ;
reg  WBC ;
reg  WBD ;
reg  WBE ;
reg  WBF ;
reg  WBG ;
reg  WBH ;
reg  wbi ;
reg  wbj ;
reg  wbk ;
reg  wbl ;
reg  wbm ;
reg  wbn ;
reg  wbo ;
reg  wbp ;
reg  WCA ;
reg  WCB ;
reg  WCC ;
reg  WCD ;
reg  WCE ;
reg  WCF ;
reg  WCG ;
reg  WCH ;
reg  wci ;
reg  wcj ;
reg  wck ;
reg  wcl ;
reg  wcm ;
reg  wcn ;
reg  wco ;
reg  wcp ;
reg  WDA ;
reg  WDB ;
reg  WDC ;
reg  WDD ;
reg  WDE ;
reg  WDF ;
reg  WDG ;
reg  WDH ;
reg  wdi ;
reg  wdj ;
reg  wdk ;
reg  wdl ;
reg  wdm ;
reg  wdn ;
reg  wdo ;
reg  wdp ;
wire  aaa ;
wire  aab ;
wire  aac ;
wire  aad ;
wire  aae ;
wire  aaf ;
wire  aag ;
wire  aah ;
wire  aai ;
wire  aaj ;
wire  aak ;
wire  aal ;
wire  aba ;
wire  abb ;
wire  abc ;
wire  abd ;
wire  abe ;
wire  abf ;
wire  abg ;
wire  abh ;
wire  abi ;
wire  abj ;
wire  abk ;
wire  abl ;
wire  aca ;
wire  acb ;
wire  acc ;
wire  acd ;
wire  ace ;
wire  acf ;
wire  acg ;
wire  ach ;
wire  aci ;
wire  acj ;
wire  ack ;
wire  acl ;
wire  ada ;
wire  adb ;
wire  adc ;
wire  add ;
wire  ade ;
wire  adf ;
wire  adg ;
wire  adh ;
wire  adi ;
wire  adj ;
wire  adk ;
wire  adl ;
wire  aea ;
wire  aeb ;
wire  aec ;
wire  aed ;
wire  aee ;
wire  aef ;
wire  aeg ;
wire  aeh ;
wire  aei ;
wire  aej ;
wire  aek ;
wire  ael ;
wire  afa ;
wire  afb ;
wire  afc ;
wire  afd ;
wire  afe ;
wire  aff ;
wire  afg ;
wire  afh ;
wire  afi ;
wire  afj ;
wire  afk ;
wire  afl ;
wire  aga ;
wire  agb ;
wire  agc ;
wire  agd ;
wire  age ;
wire  agf ;
wire  agg ;
wire  agh ;
wire  agi ;
wire  agj ;
wire  agk ;
wire  agl ;
wire  aha ;
wire  ahb ;
wire  ahc ;
wire  ahd ;
wire  ahe ;
wire  ahf ;
wire  ahg ;
wire  ahh ;
wire  ahi ;
wire  ahj ;
wire  ahk ;
wire  ahl ;
wire  baa ;
wire  bab ;
wire  bac ;
wire  bad ;
wire  bae ;
wire  baf ;
wire  bag ;
wire  bah ;
wire  bai ;
wire  baj ;
wire  bak ;
wire  bal ;
wire  bam ;
wire  ban ;
wire  bao ;
wire  bap ;
wire  bba ;
wire  bbb ;
wire  bbc ;
wire  bbd ;
wire  bbe ;
wire  bbf ;
wire  bbg ;
wire  bbh ;
wire  bbi ;
wire  bbj ;
wire  bbk ;
wire  bbl ;
wire  bbm ;
wire  bbn ;
wire  bbo ;
wire  bbp ;
wire  bca ;
wire  bcb ;
wire  bcc ;
wire  bcd ;
wire  bce ;
wire  bcf ;
wire  bcg ;
wire  bch ;
wire  bci ;
wire  bcj ;
wire  bck ;
wire  bcl ;
wire  bcm ;
wire  bcn ;
wire  bco ;
wire  bcp ;
wire  bda ;
wire  bdb ;
wire  bdc ;
wire  bdd ;
wire  bde ;
wire  bdf ;
wire  bdg ;
wire  bdh ;
wire  bdi ;
wire  bdj ;
wire  bdk ;
wire  bdl ;
wire  bdm ;
wire  bdn ;
wire  bdo ;
wire  bdp ;
wire  bea ;
wire  beb ;
wire  bec ;
wire  bed ;
wire  bee ;
wire  bef ;
wire  beg ;
wire  beh ;
wire  bei ;
wire  bej ;
wire  bek ;
wire  bel ;
wire  bem ;
wire  ben ;
wire  beo ;
wire  bep ;
wire  bfa ;
wire  bfb ;
wire  bfc ;
wire  bfd ;
wire  bfe ;
wire  bff ;
wire  bfg ;
wire  bfh ;
wire  bfi ;
wire  bfj ;
wire  bfk ;
wire  bfl ;
wire  bfm ;
wire  bfn ;
wire  bfo ;
wire  bfp ;
wire  bga ;
wire  bgb ;
wire  bgc ;
wire  bgd ;
wire  bge ;
wire  bgf ;
wire  bgg ;
wire  bgh ;
wire  bgi ;
wire  bgj ;
wire  bgk ;
wire  bgl ;
wire  bgm ;
wire  bgn ;
wire  bgo ;
wire  bgp ;
wire  bha ;
wire  bhb ;
wire  bhc ;
wire  bhd ;
wire  bhe ;
wire  bhf ;
wire  bhg ;
wire  bhh ;
wire  bhi ;
wire  bhj ;
wire  bhk ;
wire  bhl ;
wire  bhm ;
wire  bhn ;
wire  bho ;
wire  bhp ;
wire  faa ;
wire  fab ;
wire  fac ;
wire  fad ;
wire  fae ;
wire  faf ;
wire  fag ;
wire  fah ;
wire  fai ;
wire  faj ;
wire  fak ;
wire  fal ;
wire  fao ;
wire  FAO ;
wire  fap ;
wire  FAP ;
wire  faq ;
wire  FAQ ;
wire  fba ;
wire  fbb ;
wire  fbc ;
wire  fbd ;
wire  fbe ;
wire  fbf ;
wire  fbg ;
wire  fbh ;
wire  fbi ;
wire  fbj ;
wire  fbk ;
wire  fbl ;
wire  fbo ;
wire  FBO ;
wire  fbp ;
wire  FBP ;
wire  gaa ;
wire  gab ;
wire  gac ;
wire  gad ;
wire  gae ;
wire  gaf ;
wire  gag ;
wire  gah ;
wire  gai ;
wire  gaj ;
wire  gak ;
wire  gal ;
wire  iaa ;
wire  iab ;
wire  iac ;
wire  iad ;
wire  iae ;
wire  iaf ;
wire  iag ;
wire  iah ;
wire  iai ;
wire  iaj ;
wire  iak ;
wire  ial ;
wire  iam ;
wire  ian ;
wire  iao ;
wire  iap ;
wire  iba ;
wire  ibb ;
wire  ibc ;
wire  ibd ;
wire  ibe ;
wire  ibf ;
wire  ibg ;
wire  ibh ;
wire  ibi ;
wire  ibj ;
wire  ibk ;
wire  ibl ;
wire  ibm ;
wire  ibn ;
wire  ibo ;
wire  ibp ;
wire  ica ;
wire  icb ;
wire  icc ;
wire  icd ;
wire  ice ;
wire  icf ;
wire  icg ;
wire  ich ;
wire  ici ;
wire  icj ;
wire  ick ;
wire  icl ;
wire  icm ;
wire  icn ;
wire  ico ;
wire  icp ;
wire  ida ;
wire  idb ;
wire  idc ;
wire  idd ;
wire  ide ;
wire  idf ;
wire  idg ;
wire  idh ;
wire  idi ;
wire  idj ;
wire  idk ;
wire  idl ;
wire  idm ;
wire  idn ;
wire  ido ;
wire  idp ;
wire  iea ;
wire  ieb ;
wire  iec ;
wire  ied ;
wire  iee ;
wire  ief ;
wire  ieg ;
wire  ieh ;
wire  iei ;
wire  iej ;
wire  iek ;
wire  iel ;
wire  iem ;
wire  ien ;
wire  ieo ;
wire  iep ;
wire  ifa ;
wire  ifb ;
wire  ifc ;
wire  ifd ;
wire  ife ;
wire  ifff  ;
wire  ifg ;
wire  ifh ;
wire  ifi ;
wire  ifj ;
wire  ifk ;
wire  ifl ;
wire  ifm ;
wire  ifn ;
wire  ifo ;
wire  ifp ;
wire  iga ;
wire  igb ;
wire  igc ;
wire  igd ;
wire  ige ;
wire  igf ;
wire  igg ;
wire  igh ;
wire  igi ;
wire  igj ;
wire  igk ;
wire  igl ;
wire  igm ;
wire  ign ;
wire  igo ;
wire  igp ;
wire  iha ;
wire  ihb ;
wire  iia ;
wire  iib ;
wire  ija ;
wire  ijb ;
wire  ijc ;
wire  ijd ;
wire  jca ;
wire  JCA ;
wire  jcb ;
wire  JCB ;
wire  jcc ;
wire  JCC ;
wire  jcd ;
wire  JCD ;
wire  jda ;
wire  JDA ;
wire  jdb ;
wire  JDB ;
wire  jdc ;
wire  JDC ;
wire  jdd ;
wire  JDD ;
wire  jea ;
wire  JEA ;
wire  jeb ;
wire  JEB ;
wire  jec ;
wire  JEC ;
wire  jed ;
wire  JED ;
wire  jma ;
wire  jmb ;
wire  jmc ;
wire  jmd ;
wire  jme ;
wire  jmf ;
wire  jmg ;
wire  jmh ;
wire  kaa ;
wire  kab ;
wire  kac ;
wire  kad ;
wire  kae ;
wire  kaf ;
wire  kag ;
wire  kah ;
wire  kai ;
wire  kaj ;
wire  kak ;
wire  kal ;
wire  kam ;
wire  kan ;
wire  kao ;
wire  kap ;
wire  maa ;
wire  mab ;
wire  mac ;
wire  mad ;
wire  mae ;
wire  maf ;
wire  mag ;
wire  mah ;
wire  mai ;
wire  maj ;
wire  mak ;
wire  mal ;
wire  mam ;
wire  man ;
wire  mao ;
wire  map ;
wire  maq ;
wire  mar ;
wire  mas ;
wire  mat ;
wire  mau ;
wire  mav ;
wire  maw ;
wire  max ;
wire  naa ;
wire  nab ;
wire  nac ;
wire  nad ;
wire  nae ;
wire  naf ;
wire  nag ;
wire  nah ;
wire  nai ;
wire  naj ;
wire  nak ;
wire  nal ;
wire  nam ;
wire  nan ;
wire  nao ;
wire  nap ;
wire  nba ;
wire  nbb ;
wire  nbc ;
wire  nbd ;
wire  nbe ;
wire  nbf ;
wire  nbg ;
wire  nbh ;
wire  nbi ;
wire  nbj ;
wire  nbk ;
wire  nbl ;
wire  nbm ;
wire  nbn ;
wire  nbo ;
wire  nbp ;
wire  nca ;
wire  ncb ;
wire  ncc ;
wire  ncd ;
wire  nce ;
wire  ncf ;
wire  ncg ;
wire  nch ;
wire  NCI ;
wire  NCJ ;
wire  NCK ;
wire  NCL ;
wire  NCM ;
wire  NCN ;
wire  NCO ;
wire  NCP ;
wire  nda ;
wire  ndb ;
wire  ndc ;
wire  ndd ;
wire  nde ;
wire  ndf ;
wire  ndg ;
wire  ndh ;
wire  NDI ;
wire  NDJ ;
wire  NDK ;
wire  NDL ;
wire  NDM ;
wire  NDN ;
wire  NDO ;
wire  NDP ;
wire  oaa ;
wire  oab ;
wire  oac ;
wire  oad ;
wire  oae ;
wire  oaf ;
wire  oag ;
wire  oah ;
wire  oai ;
wire  oaj ;
wire  oak ;
wire  oal ;
wire  oam ;
wire  oan ;
wire  oao ;
wire  oap ;
wire  oba ;
wire  obb ;
wire  obc ;
wire  obd ;
wire  obe ;
wire  obf ;
wire  obg ;
wire  obh ;
wire  obi ;
wire  obj ;
wire  obk ;
wire  obl ;
wire  obm ;
wire  obn ;
wire  obo ;
wire  obp ;
wire  oca ;
wire  ocb ;
wire  occ ;
wire  ocd ;
wire  oce ;
wire  ocf ;
wire  ocg ;
wire  och ;
wire  oci ;
wire  ocj ;
wire  ock ;
wire  ocl ;
wire  ocm ;
wire  ocn ;
wire  oco ;
wire  ocp ;
wire  oda ;
wire  odb ;
wire  odc ;
wire  odd ;
wire  ode ;
wire  odf ;
wire  odg ;
wire  odh ;
wire  odi ;
wire  odj ;
wire  odk ;
wire  odl ;
wire  odm ;
wire  odn ;
wire  odo ;
wire  odp ;
wire  oea ;
wire  oeb ;
wire  oec ;
wire  oed ;
wire  oee ;
wire  oef ;
wire  oeg ;
wire  oeh ;
wire  oei ;
wire  oej ;
wire  oek ;
wire  oel ;
wire  oem ;
wire  oen ;
wire  oeo ;
wire  oep ;
wire  ofa ;
wire  ofb ;
wire  ofc ;
wire  ofd ;
wire  ofe ;
wire  off ;
wire  ofg ;
wire  ofh ;
wire  ofi ;
wire  ofj ;
wire  ofk ;
wire  ofl ;
wire  ofm ;
wire  ofn ;
wire  ofo ;
wire  ofp ;
wire  oha ;
wire  ohb ;
wire  ohc ;
wire  ohd ;
wire  ohe ;
wire  ohf ;
wire  ohg ;
wire  ohh ;
wire  paa ;
wire  pab ;
wire  pac ;
wire  pad ;
wire  pba ;
wire  pbb ;
wire  pbc ;
wire  pbd ;
wire  pca ;
wire  pcb ;
wire  pcc ;
wire  pcd ;
wire  pce ;
wire  pcf ;
wire  pcg ;
wire  pch ;
wire  pda ;
wire  pdb ;
wire  pdc ;
wire  pdd ;
wire  pea ;
wire  peb ;
wire  pec ;
wire  ped ;
wire  qaa ;
wire  qab ;
wire  qac ;
wire  qbb ;
wire  qbc ;
wire  qbd ;
wire  qda ;
wire  qdb ;
wire  qdc ;
wire  qfa ;
wire  taa ;
wire  TAA ;
wire  tab ;
wire  TAB ;
wire  tac ;
wire  TAC ;
wire  tad ;
wire  TAD ;
wire  tba ;
wire  TBA ;
wire  tbb ;
wire  TBB ;
wire  tbc ;
wire  TBC ;
wire  tbd ;
wire  TBD ;
wire  tca ;
wire  TCA ;
wire  tcb ;
wire  TCB ;
wire  tcc ;
wire  TCC ;
wire  tcd ;
wire  TCD ;
wire  tda ;
wire  TDA ;
wire  tdb ;
wire  TDB ;
wire  tdc ;
wire  TDC ;
wire  tdd ;
wire  TDD ;
wire  tea ;
wire  teb ;
wire  tec ;
wire  ted ;
wire  tee ;
wire  tef ;
wire  teg ;
wire  teh ;
wire  tei ;
wire  tej ;
wire  TEK ;
wire  TEL ;
wire  TEM ;
wire  TEN ;
wire  TEO ;
wire  TEP ;
wire  TEQ ;
wire  TER ;
wire  tfa ;
wire  tfb ;
wire  tfc ;
wire  tfd ;
wire  tfe ;
wire  tff ;
wire  tfg ;
wire  tfh ;
wire  tfi ;
wire  tfj ;
wire  TFK ;
wire  TFL ;
wire  TFM ;
wire  TFN ;
wire  TFO ;
wire  TFP ;
wire  TFQ ;
wire  TFR ;
wire  tga ;
wire  tgb ;
wire  tgc ;
wire  tgd ;
wire  tge ;
wire  tgf ;
wire  tgg ;
wire  tgh ;
wire  tgi ;
wire  tgj ;
wire  TGK ;
wire  TGL ;
wire  TGM ;
wire  TGN ;
wire  TGO ;
wire  TGP ;
wire  TGQ ;
wire  TGR ;
wire  tha ;
wire  thb ;
wire  thc ;
wire  thd ;
wire  the ;
wire  thf ;
wire  thg ;
wire  thh ;
wire  thi ;
wire  thj ;
wire  THK ;
wire  THL ;
wire  THM ;
wire  THN ;
wire  THO ;
wire  THP ;
wire  THQ ;
wire  THR ;
wire  tla ;
wire  TLA ;
wire  tma ;
wire  tmb ;
wire  tmc ;
wire  tmd ;
wire  tme ;
wire  tmf ;
wire  tmg ;
wire  tmh ;
wire  tna ;
wire  TNA ;
wire  tnb ;
wire  TNB ;
wire  tnc ;
wire  TNC ;
wire  tnd ;
wire  TND ;
wire  tne ;
wire  TNE ;
wire  tnf ;
wire  TNF ;
wire  tng ;
wire  TNG ;
wire  tnh ;
wire  TNH ;
wire  toa ;
wire  TOA ;
wire  tob ;
wire  TOB ;
wire  toc ;
wire  TOC ;
wire  tod ;
wire  TOD ;
wire  toe ;
wire  TOE ;
wire  tof ;
wire  TOF ;
wire  tog ;
wire  TOG ;
wire  toh ;
wire  TOH ;
wire  tua ;
wire  tub ;
wire  tuc ;
wire  tud ;
wire  tue ;
wire  tuf ;
wire  tug ;
wire  tuh ;
wire  tui ;
wire  tuj ;
wire  TUK ;
wire  TUL ;
wire  TUM ;
wire  TUN ;
wire  TUO ;
wire  TUP ;
wire  TUQ ;
wire  TUR ;
wire  tva ;
wire  tvb ;
wire  tvc ;
wire  tvd ;
wire  tve ;
wire  tvf ;
wire  tvg ;
wire  tvh ;
wire  tvi ;
wire  tvj ;
wire  TVK ;
wire  TVL ;
wire  TVM ;
wire  TVN ;
wire  TVO ;
wire  TVP ;
wire  TVQ ;
wire  TVR ;
wire  twa ;
wire  twb ;
wire  twc ;
wire  twd ;
wire  twe ;
wire  twf ;
wire  twg ;
wire  twh ;
wire  twi ;
wire  twj ;
wire  TWK ;
wire  TWL ;
wire  TWM ;
wire  TWN ;
wire  TWO ;
wire  TWP ;
wire  TWQ ;
wire  TWR ;
wire  txa ;
wire  txb ;
wire  txc ;
wire  txd ;
wire  txe ;
wire  txf ;
wire  txg ;
wire  txh ;
wire  txi ;
wire  txj ;
wire  TXK ;
wire  TXL ;
wire  TXM ;
wire  TXN ;
wire  TXO ;
wire  TXP ;
wire  TXQ ;
wire  TXR ;
wire  waa ;
wire  wab ;
wire  wac ;
wire  wad ;
wire  wae ;
wire  waf ;
wire  wag ;
wire  wah ;
wire  WAI ;
wire  WAJ ;
wire  WAK ;
wire  WAL ;
wire  WAM ;
wire  WAN ;
wire  WAO ;
wire  WAP ;
wire  wba ;
wire  wbb ;
wire  wbc ;
wire  wbd ;
wire  wbe ;
wire  wbf ;
wire  wbg ;
wire  wbh ;
wire  WBI ;
wire  WBJ ;
wire  WBK ;
wire  WBL ;
wire  WBM ;
wire  WBN ;
wire  WBO ;
wire  WBP ;
wire  wca ;
wire  wcb ;
wire  wcc ;
wire  wcd ;
wire  wce ;
wire  wcf ;
wire  wcg ;
wire  wch ;
wire  WCI ;
wire  WCJ ;
wire  WCK ;
wire  WCL ;
wire  WCM ;
wire  WCN ;
wire  WCO ;
wire  WCP ;
wire  wda ;
wire  wdb ;
wire  wdc ;
wire  wdd ;
wire  wde ;
wire  wdf ;
wire  wdg ;
wire  wdh ;
wire  WDI ;
wire  WDJ ;
wire  WDK ;
wire  WDL ;
wire  WDM ;
wire  WDN ;
wire  WDO ;
wire  WDP ;
wire  ZZI ;
wire  ZZO ;
   
wire SAA;
wire SAB;
wire SAC;
wire SAD;
wire SAE;
wire SAF;
wire SAG;
wire SAH;
wire SAI;
wire SAJ;
wire SAK;
wire SAL;
wire SAM;
wire SAN;
wire SAO;
wire SAP;
wire SBA;
wire SBB;
wire SBC;
wire SBD;
wire SBE;
wire SBF;
wire SBG;
wire SBH;
wire SBI;
wire SBJ;
wire SBK;
wire SBL;
wire SBM;
wire SBN;
wire SBO;
wire SBP;
wire SCA;
wire SCB;
wire SCC;
wire SCD;
wire SCE;
wire SCF;
wire SCG;
wire SCH;
wire SCI;
wire SCJ;
wire SCK;
wire SCL;
wire SCM;
wire SCN;
wire SCO;
wire SCP;
wire SDA;
wire SDB;
wire SDC;
wire SDD;
wire SDE;
wire SDF;
wire SDG;
wire SDH;
wire SDI;
wire SDJ;
wire SDK;
wire SDL;
wire SDM;
wire SDN;
wire SDO;
wire SDP;
wire SEA;
wire SEB;
wire SEC;
wire SED;
wire SEE;
wire SEF;
wire SEG;
wire SEH;
wire SEI;
wire SEJ;
wire SEK;
wire SEL;
wire SEM;
wire SEN;
wire SEO;
wire SEP;
wire SFA;
wire SFB;
wire SFC;
wire SFD;
wire SFE;
wire SFF;
wire SFG;
wire SFH;
wire SFI;
wire SFJ;
wire SFK;
wire SFL;
wire SFM;
wire SFN;
wire SFO;
wire SFP;
wire SGA;
wire SGB;
wire SGC;
wire SGD;
wire SGE;
wire SGF;
wire SGG;
wire SGH;
wire SGI;
wire SGJ;
wire SGK;
wire SGL;
wire SGM;
wire SGN;
wire SGO;
wire SGP;
wire SHA;
wire SHB;
wire SHC;
wire SHD;
wire SHE;
wire SHF;
wire SHG;
wire SHH;
wire SHI;
wire SHJ;
wire SHK;
wire SHL;
wire SHM;
wire SHN;
wire SHO;
wire SHP;
wire SIA;
wire SIB;
wire SIC;
wire SID;
wire SIE;
wire SIF;
wire SIG;
wire SIH;
wire SII;
wire SIJ;
wire SIK;
wire SIL;
wire SIM;
wire SIN;
wire SIO;
wire SIP;
wire SJA;
wire SJB;
wire SJC;
wire SJD;
wire SJE;
wire SJF;
wire SJG;
wire SJH;
wire SJI;
wire SJJ;
wire SJK;
wire SJL;
wire SJM;
wire SJN;
wire SJO;
wire SJP;
wire SKA;
wire SKB;
wire SKC;
wire SKD;
wire SKE;
wire SKF;
wire SKG;
wire SKH;
wire SKI;
wire SKJ;
wire SKK;
wire SKL;
wire SKM;
wire SKN;
wire SKO;
wire SKP;
wire SLA;
wire SLB;
wire SLC;
wire SLD;
wire SLE;
wire SLF;
wire SLG;
wire SLH;
wire SLI;
wire SLJ;
wire SLK;
wire SLL;
wire SLM;
wire SLN;
wire SLO;
wire SLP;
wire SMA;
wire SMB;
wire SMC;
wire SMD;
wire SME;
wire SMF;
wire SMG;
wire SMH;
wire SMI;
wire SMJ;
wire SMK;
wire SML;
wire SMM;
wire SMN;
wire SMO;
wire SMP;
wire SNA;
wire SNB;
wire SNC;
wire SND;
wire SNE;
wire SNF;
wire SNG;
wire SNH;
wire SNI;
wire SNJ;
wire SNK;
wire SNL;
wire SNM;
wire SNN;
wire SNO;
wire SNP;
wire SOA;
wire SOB;
wire SOC;
wire SOD;
wire SOE;
wire SOF;
wire SOG;
wire SOH;
wire SOI;
wire SOJ;
wire SOK;
wire SOL;
wire SOM;
wire SON;
wire SOO;
wire SOP;
wire SPA;
wire SPB;
wire SPC;
wire SPD;
wire SPE;
wire SPF;
wire SPG;
wire SPH;
wire SPI;
wire SPJ;
wire SPK;
wire SPL;
wire SPM;
wire SPN;
wire SPO;
wire SPP;

assign ZZI = 1'b1;
assign ZZO = 1'b0;
assign bea = ~BEA;  //complement 
assign beb = ~BEB;  //complement 
assign bab = ~BAB;  //complement 
assign baa = ~BAA;  //complement 
assign bec = ~BEC;  //complement 
assign bed = ~BED;  //complement 
assign bac = ~BAC;  //complement 
assign bad = ~BAD;  //complement 
assign bee = ~BEE;  //complement 
assign bef = ~BEF;  //complement 
assign bae = ~BAE;  //complement 
assign baf = ~BAF;  //complement 
assign beg = ~BEG;  //complement 
assign beh = ~BEH;  //complement 
assign wae = ~WAE;  //complement 
assign waf = ~WAF;  //complement 
assign wag = ~WAG;  //complement 
assign wah = ~WAH;  //complement 
assign bhj = ~BHJ;  //complement 
assign bhk = ~BHK;  //complement 
assign bhl = ~BHL;  //complement 
assign bag = ~BAG;  //complement 
assign bah = ~BAH;  //complement 
assign bhm = ~BHM;  //complement 
assign bhn = ~BHN;  //complement 
assign bho = ~BHO;  //complement 
assign bhp = ~BHP;  //complement 
assign aaa = ~AAA;  //complement 
assign aab = ~AAB;  //complement 
assign aac = ~AAC;  //complement 
assign aad = ~AAD;  //complement 
assign aae = ~AAE;  //complement 
assign aaf = ~AAF;  //complement 
assign aag = ~AAG;  //complement 
assign aah = ~AAH;  //complement 
assign aai = ~AAI;  //complement 
assign aaj = ~AAJ;  //complement 
assign aak = ~AAK;  //complement 
assign aal = ~AAL;  //complement 
assign maa = ~MAA;  //complement 
assign waa = ~WAA;  //complement 
assign wab = ~WAB;  //complement 
assign wac = ~WAC;  //complement 
assign wad = ~WAD;  //complement 
assign toa = qaa; 
assign TOA = ~toa; //complement 
assign tob = qaa; 
assign TOB = ~tob;  //complement 
assign toc = qaa; 
assign TOC = ~toc;  //complement 
assign tod = qaa; 
assign TOD = ~tod;  //complement 
assign WAI = ~wai;  //complement 
assign WAJ = ~waj;  //complement 
assign WAK = ~wak;  //complement 
assign WAL = ~wal;  //complement 
assign WAM = ~wam;  //complement 
assign WAN = ~wan;  //complement 
assign WAO = ~wao;  //complement 
assign WAP = ~wap;  //complement 
assign bep = ~BEP;  //complement 
assign tga = ~TGA;  //complement 
assign tgb = ~TGB;  //complement 
assign tgc = ~TGC;  //complement 
assign tgd = ~TGD;  //complement 
assign faa = ~FAA;  //complement 
assign fab = ~FAB;  //complement 
assign fac = ~FAC;  //complement 
assign fad = ~FAD;  //complement 
assign fae = ~FAE;  //complement 
assign faf = ~FAF;  //complement 
assign fag = ~FAG;  //complement 
assign fah = ~FAH;  //complement 
assign fai = ~FAI;  //complement 
assign faj = ~FAJ;  //complement 
assign fak = ~FAK;  //complement 
assign fal = ~FAL;  //complement 
assign nai = ~NAI;  //complement 
assign naj = ~NAJ;  //complement 
assign nak = ~NAK;  //complement 
assign nal = ~NAL;  //complement 
assign oaa = ~OAA;  //complement 
assign nam = ~NAM;  //complement 
assign nan = ~NAN;  //complement 
assign nao = ~NAO;  //complement 
assign nap = ~NAP;  //complement 
assign JCA =  QFA & iea & ieb  ; 
assign jca = ~JCA;  //complement 
assign JCB =  QFA & IEA & ieb  ; 
assign jcb = ~JCB;  //complement 
assign oab = ~OAB;  //complement 
assign qac = ~QAC;  //complement 
assign qbd = ~QBD;  //complement 
assign qbb = ~QBB;  //complement 
assign qbc = ~QBC;  //complement 
assign oac = ~OAC;  //complement 
assign JCC =  QFA & iea & IEB  ; 
assign jcc = ~JCC;  //complement 
assign JCD =  QFA & IEA & IEB  ; 
assign jcd = ~JCD;  //complement 
assign oad = ~OAD;  //complement 
assign JDA =  QAA & kaa & kab  ; 
assign jda = ~JDA;  //complement 
assign JDB =  QAA & KAA & kab  ; 
assign jdb = ~JDB;  //complement 
assign JDC =  QAA & kaa & KAB  ; 
assign jdc = ~JDC;  //complement 
assign JDD =  QAA & KAA & KAB  ; 
assign jdd = ~JDD;  //complement 
assign kac = ~KAC;  //complement 
assign kad = ~KAD;  //complement 
assign oae = ~OAE;  //complement 
assign JEB =  PAB & qdc  |  PAA & QDC  ; 
assign jeb = ~JEB;  //complement 
assign JEC =  PAC & qdc  |  PAB & QDC  ; 
assign jec = ~JEC;  //complement 
assign oaf = ~OAF;  //complement 
assign TWK = ~twk;  //complement 
assign TWL = ~twl;  //complement 
assign TWM = ~twm;  //complement 
assign TWN = ~twn;  //complement 
assign kae = ~KAE;  //complement 
assign kaf = ~KAF;  //complement 
assign kag = ~KAG;  //complement 
assign kah = ~KAH;  //complement 
assign naa = ~NAA;  //complement 
assign nab = ~NAB;  //complement 
assign nac = ~NAC;  //complement 
assign nad = ~NAD;  //complement 
assign kai = ~KAI;  //complement 
assign kaj = ~KAJ;  //complement 
assign kak = ~KAK;  //complement 
assign kal = ~KAL;  //complement 
assign oag = ~OAG;  //complement 
assign kam = ~KAM;  //complement 
assign kan = ~KAN;  //complement 
assign kao = ~KAO;  //complement 
assign kap = ~KAP;  //complement 
assign oah = ~OAH;  //complement 
assign nae = ~NAE;  //complement 
assign naf = ~NAF;  //complement 
assign nag = ~NAG;  //complement 
assign nah = ~NAH;  //complement 
assign bei = ~BEI;  //complement 
assign bej = ~BEJ;  //complement 
assign bai = ~BAI;  //complement 
assign baj = ~BAJ;  //complement 
assign bek = ~BEK;  //complement 
assign bel = ~BEL;  //complement 
assign bak = ~BAK;  //complement 
assign bal = ~BAL;  //complement 
assign bem = ~BEM;  //complement 
assign ben = ~BEN;  //complement 
assign bam = ~BAM;  //complement 
assign ban = ~BAN;  //complement 
assign beo = ~BEO;  //complement 
assign bao = ~BAO;  //complement 
assign bap = ~BAP;  //complement 
assign bha = ~BHA;  //complement 
assign bhb = ~BHB;  //complement 
assign bhc = ~BHC;  //complement 
assign bhd = ~BHD;  //complement 
assign bhe = ~BHE;  //complement 
assign bhf = ~BHF;  //complement 
assign bhg = ~BHG;  //complement 
assign bhh = ~BHH;  //complement 
assign bhi = ~BHI;  //complement 
assign aba = ~ABA;  //complement 
assign abb = ~ABB;  //complement 
assign abc = ~ABC;  //complement 
assign abd = ~ABD;  //complement 
assign abe = ~ABE;  //complement 
assign abf = ~ABF;  //complement 
assign abg = ~ABG;  //complement 
assign abh = ~ABH;  //complement 
assign abi = ~ABI;  //complement 
assign abj = ~ABJ;  //complement 
assign abk = ~ABK;  //complement 
assign abl = ~ABL;  //complement 
assign kaa = ~KAA;  //complement 
assign kab = ~KAB;  //complement 
assign tge = ~TGE;  //complement 
assign tgf = ~TGF;  //complement 
assign tgg = ~TGG;  //complement 
assign tgh = ~TGH;  //complement 
assign pca = ~PCA;  //complement 
assign pcb = ~PCB;  //complement 
assign pcc = ~PCC;  //complement 
assign pcd = ~PCD;  //complement 
assign pce = ~PCE;  //complement 
assign pcf = ~PCF;  //complement 
assign pcg = ~PCG;  //complement 
assign pch = ~PCH;  //complement 
assign pda = ~PDA;  //complement 
assign pdb = ~PDB;  //complement 
assign pdc = ~PDC;  //complement 
assign pdd = ~PDD;  //complement 
assign fbb = ~FBB;  //complement 
assign fbf = ~FBF;  //complement 
assign fbj = ~FBJ;  //complement 
assign fba = ~FBA;  //complement 
assign fbe = ~FBE;  //complement 
assign fbi = ~FBI;  //complement 
assign pba = ~PBA;  //complement 
assign pbb = ~PBB;  //complement 
assign pbc = ~PBC;  //complement 
assign pbd = ~PBD;  //complement 
assign oai = ~OAI;  //complement 
assign gak = ~GAK;  //complement 
assign gal = ~GAL;  //complement 
assign toe = qaa; 
assign TOE = ~toe; //complement 
assign tof = qaa; 
assign TOF = ~tof;  //complement 
assign tog = qaa; 
assign TOG = ~tog;  //complement 
assign toh = qaa; 
assign TOH = ~toh;  //complement 
assign oaj = ~OAJ;  //complement 
assign nba = ~NBA;  //complement 
assign nbb = ~NBB;  //complement 
assign nbc = ~NBC;  //complement 
assign nbd = ~NBD;  //complement 
assign nbe = ~NBE;  //complement 
assign nbf = ~NBF;  //complement 
assign nbg = ~NBG;  //complement 
assign nbh = ~NBH;  //complement 
assign oak = ~OAK;  //complement 
assign nbi = ~NBI;  //complement 
assign nbj = ~NBJ;  //complement 
assign nbk = ~NBK;  //complement 
assign nbl = ~NBL;  //complement 
assign nbm = ~NBM;  //complement 
assign nbn = ~NBN;  //complement 
assign nbo = ~NBO;  //complement 
assign nbp = ~NBP;  //complement 
assign oal = ~OAL;  //complement 
assign JED =  PAD & qdc  |  PAC & QDC  ; 
assign jed = ~JED;  //complement 
assign JEA =  PAA & qdc  |  PAD & QDC  ; 
assign jea = ~JEA;  //complement 
assign oam = ~OAM;  //complement 
assign WBI = ~wbi;  //complement 
assign WBJ = ~wbj;  //complement 
assign WBK = ~wbk;  //complement 
assign WBL = ~wbl;  //complement 
assign WBM = ~wbm;  //complement 
assign WBN = ~wbn;  //complement 
assign WBO = ~wbo;  //complement 
assign WBP = ~wbp;  //complement 
assign oan = ~OAN;  //complement 
assign wba = ~WBA;  //complement 
assign wbb = ~WBB;  //complement 
assign wbc = ~WBC;  //complement 
assign wbd = ~WBD;  //complement 
assign wbe = ~WBE;  //complement 
assign wbf = ~WBF;  //complement 
assign wbg = ~WBG;  //complement 
assign wbh = ~WBH;  //complement 
assign oao = ~OAO;  //complement 
assign gaa = ~GAA;  //complement 
assign gab = ~GAB;  //complement 
assign gac = ~GAC;  //complement 
assign gad = ~GAD;  //complement 
assign gae = ~GAE;  //complement 
assign gaf = ~GAF;  //complement 
assign oap = ~OAP;  //complement 
assign gag = ~GAG;  //complement 
assign gah = ~GAH;  //complement 
assign gai = ~GAI;  //complement 
assign gaj = ~GAJ;  //complement 
assign bfa = ~BFA;  //complement 
assign bfb = ~BFB;  //complement 
assign bba = ~BBA;  //complement 
assign bbb = ~BBB;  //complement 
assign bfc = ~BFC;  //complement 
assign bfd = ~BFD;  //complement 
assign bbc = ~BBC;  //complement 
assign bbd = ~BBD;  //complement 
assign bfe = ~BFE;  //complement 
assign bff = ~BFF;  //complement 
assign bbe = ~BBE;  //complement 
assign bbf = ~BBF;  //complement 
assign bfg = ~BFG;  //complement 
assign bfh = ~BFH;  //complement 
assign bbg = ~BBG;  //complement 
assign bbh = ~BBH;  //complement 
assign TGM = ~tgm;  //complement 
assign TGN = ~tgn;  //complement 
assign TGO = ~tgo;  //complement 
assign TGP = ~tgp;  //complement 
assign tda =  pbb & pbd  |  qbb  ; 
assign TDA = ~tda;  //complement 
assign tdb =  pbb & pbd  |  qbb  ; 
assign TDB = ~tdb;  //complement 
assign tha = ~THA;  //complement 
assign thb = ~THB;  //complement 
assign thc = ~THC;  //complement 
assign thd = ~THD;  //complement 
assign pea = ~PEA;  //complement 
assign peb = ~PEB;  //complement 
assign pec = ~PEC;  //complement 
assign ped = ~PED;  //complement 
assign the = ~THE;  //complement 
assign thf = ~THF;  //complement 
assign thg = ~THG;  //complement 
assign thh = ~THH;  //complement 
assign aca = ~ACA;  //complement 
assign acb = ~ACB;  //complement 
assign acc = ~ACC;  //complement 
assign acd = ~ACD;  //complement 
assign ace = ~ACE;  //complement 
assign acf = ~ACF;  //complement 
assign acg = ~ACG;  //complement 
assign ach = ~ACH;  //complement 
assign aci = ~ACI;  //complement 
assign acj = ~ACJ;  //complement 
assign ack = ~ACK;  //complement 
assign acl = ~ACL;  //complement 
assign mab = ~MAB;  //complement 
assign tgi = ~TGI;  //complement 
assign tgj = ~TGJ;  //complement 
assign TGK = ~tgk;  //complement 
assign TGL = ~tgl;  //complement 
assign tfe = ~TFE;  //complement 
assign tff = ~TFF;  //complement 
assign tfg = ~TFG;  //complement 
assign tfh = ~TFH;  //complement 
assign tfi = ~TFI;  //complement 
assign tfj = ~TFJ;  //complement 
assign TFK = ~tfk;  //complement 
assign TFL = ~tfl;  //complement 
assign TFM = ~tfm;  //complement 
assign TFN = ~tfn;  //complement 
assign TFO = ~tfo;  //complement 
assign TFP = ~tfp;  //complement 
assign THM = ~thm;  //complement 
assign THN = ~thn;  //complement 
assign THO = ~tho;  //complement 
assign THP = ~thp;  //complement 
assign jma = ~JMA;  //complement 
assign thi = ~THI;  //complement 
assign thj = ~THJ;  //complement 
assign THK = ~thk;  //complement 
assign THL = ~thl;  //complement 
assign tfa = ~TFA;  //complement 
assign tfb = ~TFB;  //complement 
assign tfc = ~TFC;  //complement 
assign tfd = ~TFD;  //complement 
assign oba = ~OBA;  //complement 
assign jmc = ~JMC;  //complement 
assign jmd = ~JMD;  //complement 
assign obb = ~OBB;  //complement 
assign NDM = ~ndm;  //complement 
assign NDN = ~ndn;  //complement 
assign NDO = ~ndo;  //complement 
assign NDP = ~ndp;  //complement 
assign qda = ~QDA;  //complement 
assign qdb = ~QDB;  //complement 
assign qdc = ~QDC;  //complement 
assign qfa = ~QFA;  //complement 
assign obc = ~OBC;  //complement 
assign THQ = ~thq;  //complement 
assign THR = ~thr;  //complement 
assign TGQ = ~tgq;  //complement 
assign TGR = ~tgr;  //complement 
assign TEQ = ~teq;  //complement 
assign TER = ~ter;  //complement 
assign TFQ = ~tfq;  //complement 
assign TFR = ~tfr;  //complement 
assign obd = ~OBD;  //complement 
assign tma = ~TMA;  //complement 
assign tmb = ~TMB;  //complement 
assign tmc = ~TMC;  //complement 
assign tmd = ~TMD;  //complement 
assign tme = ~TME;  //complement 
assign tmf = ~TMF;  //complement 
assign tmg = ~TMG;  //complement 
assign tmh = ~TMH;  //complement 
assign obe = ~OBE;  //complement 
assign tna = qfa; 
assign TNA = ~tna; //complement 
assign tnb = qfa; 
assign TNB = ~tnb;  //complement 
assign tnc = qfa; 
assign TNC = ~tnc;  //complement 
assign tnd = qfa; 
assign TND = ~tnd;  //complement 
assign tne = qfa; 
assign TNE = ~tne; //complement 
assign tnf = qfa; 
assign TNF = ~tnf;  //complement 
assign tng = qfa; 
assign TNG = ~tng;  //complement 
assign tnh = qfa; 
assign TNH = ~tnh;  //complement 
assign obf = ~OBF;  //complement 
assign obg = ~OBG;  //complement 
assign paa = ~PAA;  //complement 
assign jmb = ~JMB;  //complement 
assign obi = ~OBI;  //complement 
assign nda = ~NDA;  //complement 
assign ndb = ~NDB;  //complement 
assign ndc = ~NDC;  //complement 
assign ndd = ~NDD;  //complement 
assign nde = ~NDE;  //complement 
assign ndf = ~NDF;  //complement 
assign ndg = ~NDG;  //complement 
assign ndh = ~NDH;  //complement 
assign obh = ~OBH;  //complement 
assign NDI = ~ndi;  //complement 
assign NDJ = ~ndj;  //complement 
assign NDK = ~ndk;  //complement 
assign NDL = ~ndl;  //complement 
assign bfi = ~BFI;  //complement 
assign bfj = ~BFJ;  //complement 
assign bbi = ~BBI;  //complement 
assign bbj = ~BBJ;  //complement 
assign bfk = ~BFK;  //complement 
assign bfl = ~BFL;  //complement 
assign bbk = ~BBK;  //complement 
assign bbl = ~BBL;  //complement 
assign bfm = ~BFM;  //complement 
assign bfn = ~BFN;  //complement 
assign bbm = ~BBM;  //complement 
assign bbn = ~BBN;  //complement 
assign bfo = ~BFO;  //complement 
assign bfp = ~BFP;  //complement 
assign bbo = ~BBO;  //complement 
assign bbp = ~BBP;  //complement 
assign TUM = ~tum;  //complement 
assign TUN = ~tun;  //complement 
assign TUO = ~tuo;  //complement 
assign TUP = ~tup;  //complement 
assign tva = ~TVA;  //complement 
assign tvb = ~TVB;  //complement 
assign tvc = ~TVC;  //complement 
assign tvd = ~TVD;  //complement 
assign pac = ~PAC;  //complement 
assign pad = ~PAD;  //complement 
assign tua = ~TUA;  //complement 
assign tub = ~TUB;  //complement 
assign tuc = ~TUC;  //complement 
assign tud = ~TUD;  //complement 
assign tve = ~TVE;  //complement 
assign tvf = ~TVF;  //complement 
assign tvg = ~TVG;  //complement 
assign tvh = ~TVH;  //complement 
assign tue = ~TUE;  //complement 
assign tuf = ~TUF;  //complement 
assign tug = ~TUG;  //complement 
assign tuh = ~TUH;  //complement 
assign tui = ~TUI;  //complement 
assign tuj = ~TUJ;  //complement 
assign TUK = ~tuk;  //complement 
assign TUL = ~tul;  //complement 
assign ada = ~ADA;  //complement 
assign adb = ~ADB;  //complement 
assign adc = ~ADC;  //complement 
assign add = ~ADD;  //complement 
assign ade = ~ADE;  //complement 
assign adf = ~ADF;  //complement 
assign adg = ~ADG;  //complement 
assign adh = ~ADH;  //complement 
assign adi = ~ADI;  //complement 
assign adj = ~ADJ;  //complement 
assign adk = ~ADK;  //complement 
assign adl = ~ADL;  //complement 
assign TXK = ~txk;  //complement 
assign TXL = ~txl;  //complement 
assign TXM = ~txm;  //complement 
assign TXN = ~txn;  //complement 
assign pab = ~PAB;  //complement 
assign obj = ~OBJ;  //complement 
assign oed = ~OED;  //complement 
assign oee = ~OEE;  //complement 
assign oef = ~OEF;  //complement 
assign obk = ~OBK;  //complement 
assign oeg = ~OEG;  //complement 
assign oeh = ~OEH;  //complement 
assign qaa = ~QAA;  //complement 
assign obl = ~OBL;  //complement 
assign nca = ~NCA;  //complement 
assign ncb = ~NCB;  //complement 
assign ncc = ~NCC;  //complement 
assign ncd = ~NCD;  //complement 
assign nce = ~NCE;  //complement 
assign ncf = ~NCF;  //complement 
assign ncg = ~NCG;  //complement 
assign nch = ~NCH;  //complement 
assign NCI = ~nci;  //complement 
assign NCJ = ~ncj;  //complement 
assign NCK = ~nck;  //complement 
assign NCL = ~ncl;  //complement 
assign obm = ~OBM;  //complement 
assign NCM = ~ncm;  //complement 
assign NCN = ~ncn;  //complement 
assign NCO = ~nco;  //complement 
assign NCP = ~ncp;  //complement 
assign qab = ~QAB;  //complement 
assign tea = ~TEA;  //complement 
assign teb = ~TEB;  //complement 
assign tec = ~TEC;  //complement 
assign ted = ~TED;  //complement 
assign obn = ~OBN;  //complement 
assign wca = ~WCA;  //complement 
assign wcb = ~WCB;  //complement 
assign wcc = ~WCC;  //complement 
assign wcd = ~WCD;  //complement 
assign wce = ~WCE;  //complement 
assign wcf = ~WCF;  //complement 
assign wcg = ~WCG;  //complement 
assign wch = ~WCH;  //complement 
assign WCI = ~wci;  //complement 
assign WCJ = ~wcj;  //complement 
assign WCK = ~wck;  //complement 
assign WCL = ~wcl;  //complement 
assign WCM = ~wcm;  //complement 
assign WCN = ~wcn;  //complement 
assign WCO = ~wco;  //complement 
assign WCP = ~wcp;  //complement 
assign taa =  pba & pbc  |  qbc  ; 
assign TAA = ~taa;  //complement 
assign tab =  pba & pbc  |  qbc  ; 
assign TAB = ~tab;  //complement 
assign tba =  pba & pbc  |  qbb  ; 
assign TBA = ~tba;  //complement 
assign tbb =  pba & pbc  |  qbb  ; 
assign TBB = ~tbb;  //complement 
assign tca =  pbb & pbd  |  qbc  ; 
assign TCA = ~tca;  //complement 
assign tcb =  pbb & pbd  |  qbc  ; 
assign TCB = ~tcb;  //complement 
assign obo = ~OBO;  //complement 
assign twa = ~TWA;  //complement 
assign twb = ~TWB;  //complement 
assign twc = ~TWC;  //complement 
assign twd = ~TWD;  //complement 
assign twe = ~TWE;  //complement 
assign twf = ~TWF;  //complement 
assign twg = ~TWG;  //complement 
assign twh = ~TWH;  //complement 
assign obp = ~OBP;  //complement 
assign oea = ~OEA;  //complement 
assign oeb = ~OEB;  //complement 
assign twi = ~TWI;  //complement 
assign twj = ~TWJ;  //complement 
assign oec = ~OEC;  //complement 
assign bga = ~BGA;  //complement 
assign bgb = ~BGB;  //complement 
assign bca = ~BCA;  //complement 
assign bcb = ~BCB;  //complement 
assign bgc = ~BGC;  //complement 
assign bgd = ~BGD;  //complement 
assign bcc = ~BCC;  //complement 
assign bcd = ~BCD;  //complement 
assign bge = ~BGE;  //complement 
assign bgf = ~BGF;  //complement 
assign bce = ~BCE;  //complement 
assign bcf = ~BCF;  //complement 
assign bgg = ~BGG;  //complement 
assign bgh = ~BGH;  //complement 
assign bcg = ~BCG;  //complement 
assign bch = ~BCH;  //complement 
assign tei = ~TEI;  //complement 
assign tej = ~TEJ;  //complement 
assign TEK = ~tek;  //complement 
assign TEL = ~tel;  //complement 
assign TEM = ~tem;  //complement 
assign TEN = ~ten;  //complement 
assign TEO = ~teo;  //complement 
assign TEP = ~tep;  //complement 
assign jme = ~JME;  //complement 
assign wda = ~WDA;  //complement 
assign wdb = ~WDB;  //complement 
assign wdc = ~WDC;  //complement 
assign wdd = ~WDD;  //complement 
assign wde = ~WDE;  //complement 
assign wdf = ~WDF;  //complement 
assign wdg = ~WDG;  //complement 
assign wdh = ~WDH;  //complement 
assign WDI = ~wdi;  //complement 
assign WDJ = ~wdj;  //complement 
assign WDK = ~wdk;  //complement 
assign WDL = ~wdl;  //complement 
assign aea = ~AEA;  //complement 
assign aeb = ~AEB;  //complement 
assign aec = ~AEC;  //complement 
assign aed = ~AED;  //complement 
assign aee = ~AEE;  //complement 
assign aef = ~AEF;  //complement 
assign aeg = ~AEG;  //complement 
assign aeh = ~AEH;  //complement 
assign aei = ~AEI;  //complement 
assign aej = ~AEJ;  //complement 
assign aek = ~AEK;  //complement 
assign ael = ~AEL;  //complement 
assign TXO = ~txo;  //complement 
assign TXP = ~txp;  //complement 
assign TXQ = ~txq;  //complement 
assign TXR = ~txr;  //complement 
assign tee = ~TEE;  //complement 
assign tef = ~TEF;  //complement 
assign teg = ~TEG;  //complement 
assign teh = ~TEH;  //complement 
assign oca = ~OCA;  //complement 
assign tvi = ~TVI;  //complement 
assign tvj = ~TVJ;  //complement 
assign TVK = ~tvk;  //complement 
assign TVL = ~tvl;  //complement 
assign txi = ~TXI;  //complement 
assign txj = ~TXJ;  //complement 
assign ocb = ~OCB;  //complement 
assign tac =  pba & pbc  |  qbc  ; 
assign TAC = ~tac;  //complement 
assign tad =  pba & pbc  |  qbc  ; 
assign TAD = ~tad;  //complement 
assign tbc =  pba & pbc  |  qbb  ; 
assign TBC = ~tbc;  //complement 
assign tbd =  pba & pbc  |  qbb  ; 
assign TBD = ~tbd;  //complement 
assign occ = ~OCC;  //complement 
assign TVM = ~tvm;  //complement 
assign TVN = ~tvn;  //complement 
assign TVO = ~tvo;  //complement 
assign TVP = ~tvp;  //complement 
assign TUQ = ~tuq;  //complement 
assign TUR = ~tur;  //complement 
assign ocd = ~OCD;  //complement 
assign TVQ = ~tvq;  //complement 
assign TVR = ~tvr;  //complement 
assign TWO = ~two;  //complement 
assign TWP = ~twp;  //complement 
assign TWQ = ~twq;  //complement 
assign TWR = ~twr;  //complement 
assign oce = ~OCE;  //complement 
assign ocf = ~OCF;  //complement 
assign oei = ~OEI;  //complement 
assign oej = ~OEJ;  //complement 
assign ocg = ~OCG;  //complement 
assign WDM = ~wdm;  //complement 
assign WDN = ~wdn;  //complement 
assign WDO = ~wdo;  //complement 
assign WDP = ~wdp;  //complement 
assign txa = ~TXA;  //complement 
assign txb = ~TXB;  //complement 
assign txc = ~TXC;  //complement 
assign txd = ~TXD;  //complement 
assign och = ~OCH;  //complement 
assign txe = ~TXE;  //complement 
assign txf = ~TXF;  //complement 
assign txg = ~TXG;  //complement 
assign txh = ~TXH;  //complement 
assign bgi = ~BGI;  //complement 
assign bgj = ~BGJ;  //complement 
assign bci = ~BCI;  //complement 
assign bcj = ~BCJ;  //complement 
assign bgk = ~BGK;  //complement 
assign bgl = ~BGL;  //complement 
assign bck = ~BCK;  //complement 
assign bcl = ~BCL;  //complement 
assign bgm = ~BGM;  //complement 
assign bgn = ~BGN;  //complement 
assign bcm = ~BCM;  //complement 
assign bcn = ~BCN;  //complement 
assign bgo = ~BGO;  //complement 
assign bgp = ~BGP;  //complement 
assign bco = ~BCO;  //complement 
assign bcp = ~BCP;  //complement 
assign afe = ~AFE;  //complement 
assign aff = ~AFF;  //complement 
assign afg = ~AFG;  //complement 
assign afh = ~AFH;  //complement 
assign afi = ~AFI;  //complement 
assign afj = ~AFJ;  //complement 
assign afk = ~AFK;  //complement 
assign afl = ~AFL;  //complement 
assign tcc =  pbb & pbd  |  qbc  ; 
assign TCC = ~tcc;  //complement 
assign tcd =  pbb & pbd  |  qbc  ; 
assign TCD = ~tcd;  //complement 
assign FBO =  ABA & ABB & ABC & ABD  ; 
assign fbo = ~FBO;  //complement  
assign FBP =  ABE & ABF & ABG & ABH  ; 
assign fbp = ~FBP;  //complement  
assign tdc =  pbb & pbd  |  qbb  ; 
assign TDC = ~tdc;  //complement 
assign tdd =  pbb & pbd  |  qbb  ; 
assign TDD = ~tdd;  //complement 
assign oek = ~OEK;  //complement 
assign afa = ~AFA;  //complement 
assign afb = ~AFB;  //complement 
assign oel = ~OEL;  //complement 
assign oem = ~OEM;  //complement 
assign oen = ~OEN;  //complement 
assign oeo = ~OEO;  //complement 
assign oep = ~OEP;  //complement 
assign afc = ~AFC;  //complement 
assign afd = ~AFD;  //complement 
assign oci = ~OCI;  //complement 
assign off = ~OFF;  //complement 
assign ofg = ~OFG;  //complement 
assign ofh = ~OFH;  //complement 
assign ocj = ~OCJ;  //complement 
assign fbg = ~FBG;  //complement 
assign fbk = ~FBK;  //complement 
assign ock = ~OCK;  //complement 
assign tla =  qab & qac  ; 
assign TLA = ~tla;  //complement 
assign FAO =  ABA & ABB & ABC  ; 
assign fao = ~FAO;  //complement 
assign FAP =  ABE & ABF & ABG  ; 
assign fap = ~FAP;  //complement 
assign fbd = ~FBD;  //complement 
assign ocl = ~OCL;  //complement 
assign fbh = ~FBH;  //complement 
assign fbl = ~FBL;  //complement 
assign FAQ =  ABI & ABJ & ABK  ; 
assign faq = ~FAQ;  //complement 
assign ocm = ~OCM;  //complement 
assign mac = ~MAC;  //complement 
assign mad = ~MAD;  //complement 
assign mae = ~MAE;  //complement 
assign ocn = ~OCN;  //complement 
assign maf = ~MAF;  //complement 
assign mag = ~MAG;  //complement 
assign mah = ~MAH;  //complement 
assign oco = ~OCO;  //complement 
assign ofa = ~OFA;  //complement 
assign ofb = ~OFB;  //complement 
assign ocp = ~OCP;  //complement 
assign ofc = ~OFC;  //complement 
assign ofd = ~OFD;  //complement 
assign ofe = ~OFE;  //complement 
assign fbc = ~FBC;  //complement 
assign mai = ~MAI;  //complement 
assign bda = ~BDA;  //complement 
assign bdb = ~BDB;  //complement 
assign mam = ~MAM;  //complement 
assign bdc = ~BDC;  //complement 
assign bdd = ~BDD;  //complement 
assign maj = ~MAJ;  //complement 
assign bde = ~BDE;  //complement 
assign bdf = ~BDF;  //complement 
assign bdg = ~BDG;  //complement 
assign bdh = ~BDH;  //complement 
assign mak = ~MAK;  //complement 
assign mal = ~MAL;  //complement 
assign man = ~MAN;  //complement 
assign mao = ~MAO;  //complement 
assign map = ~MAP;  //complement 
assign aga = ~AGA;  //complement 
assign agb = ~AGB;  //complement 
assign agc = ~AGC;  //complement 
assign agd = ~AGD;  //complement 
assign age = ~AGE;  //complement 
assign agf = ~AGF;  //complement 
assign agg = ~AGG;  //complement 
assign agh = ~AGH;  //complement 
assign agi = ~AGI;  //complement 
assign agj = ~AGJ;  //complement 
assign agk = ~AGK;  //complement 
assign agl = ~AGL;  //complement 
assign oda = ~ODA;  //complement 
assign odb = ~ODB;  //complement 
assign maq = ~MAQ;  //complement 
assign odc = ~ODC;  //complement 
assign mar = ~MAR;  //complement 
assign mas = ~MAS;  //complement 
assign odd = ~ODD;  //complement 
assign ode = ~ODE;  //complement 
assign mat = ~MAT;  //complement 
assign odf = ~ODF;  //complement 
assign mau = ~MAU;  //complement 
assign mav = ~MAV;  //complement 
assign odg = ~ODG;  //complement 
assign ofi = ~OFI;  //complement 
assign odh = ~ODH;  //complement 
assign jmf = ~JMF;  //complement 
assign bdi = ~BDI;  //complement 
assign bdj = ~BDJ;  //complement 
assign jmg = ~JMG;  //complement 
assign jmh = ~JMH;  //complement 
assign bdk = ~BDK;  //complement 
assign bdl = ~BDL;  //complement 
assign bdm = ~BDM;  //complement 
assign bdn = ~BDN;  //complement 
assign bdo = ~BDO;  //complement 
assign bdp = ~BDP;  //complement 
assign oha = ~OHA;  //complement 
assign ohb = ~OHB;  //complement 
assign ohc = ~OHC;  //complement 
assign ohd = ~OHD;  //complement 
assign ohe = ~OHE;  //complement 
assign ohf = ~OHF;  //complement 
assign ohg = ~OHG;  //complement 
assign ohh = ~OHH;  //complement 
assign aha = ~AHA;  //complement 
assign ahb = ~AHB;  //complement 
assign ahc = ~AHC;  //complement 
assign ahd = ~AHD;  //complement 
assign ahe = ~AHE;  //complement 
assign ahf = ~AHF;  //complement 
assign ahg = ~AHG;  //complement 
assign ahh = ~AHH;  //complement 
assign ahi = ~AHI;  //complement 
assign ahj = ~AHJ;  //complement 
assign ahk = ~AHK;  //complement 
assign ahl = ~AHL;  //complement 
assign maw = ~MAW;  //complement 
assign max = ~MAX;  //complement 
assign odi = ~ODI;  //complement 
assign ofn = ~OFN;  //complement 
assign ofo = ~OFO;  //complement 
assign ofp = ~OFP;  //complement 
assign odj = ~ODJ;  //complement 
assign odk = ~ODK;  //complement 
assign odl = ~ODL;  //complement 
assign odm = ~ODM;  //complement 
assign odn = ~ODN;  //complement 
assign odo = ~ODO;  //complement 
assign ofj = ~OFJ;  //complement 
assign ofk = ~OFK;  //complement 
assign odp = ~ODP;  //complement 
assign ofl = ~OFL;  //complement 
assign ofm = ~OFM;  //complement 
assign iaa = ~IAA; //complement 
assign iab = ~IAB; //complement 
assign iac = ~IAC; //complement 
assign iad = ~IAD; //complement 
assign iae = ~IAE; //complement 
assign iaf = ~IAF; //complement 
assign iag = ~IAG; //complement 
assign iah = ~IAH; //complement 
assign iai = ~IAI; //complement 
assign iaj = ~IAJ; //complement 
assign iak = ~IAK; //complement 
assign ial = ~IAL; //complement 
assign iam = ~IAM; //complement 
assign ian = ~IAN; //complement 
assign iao = ~IAO; //complement 
assign iap = ~IAP; //complement 
assign iba = ~IBA; //complement 
assign ibb = ~IBB; //complement 
assign ibc = ~IBC; //complement 
assign ibd = ~IBD; //complement 
assign ibe = ~IBE; //complement 
assign ibf = ~IBF; //complement 
assign ibg = ~IBG; //complement 
assign ibh = ~IBH; //complement 
assign ibi = ~IBI; //complement 
assign ibj = ~IBJ; //complement 
assign ibk = ~IBK; //complement 
assign ibl = ~IBL; //complement 
assign ibm = ~IBM; //complement 
assign ibn = ~IBN; //complement 
assign ibo = ~IBO; //complement 
assign ibp = ~IBP; //complement 
assign ica = ~ICA; //complement 
assign icb = ~ICB; //complement 
assign icc = ~ICC; //complement 
assign icd = ~ICD; //complement 
assign ice = ~ICE; //complement 
assign icf = ~ICF; //complement 
assign icg = ~ICG; //complement 
assign ich = ~ICH; //complement 
assign ici = ~ICI; //complement 
assign icj = ~ICJ; //complement 
assign ick = ~ICK; //complement 
assign icl = ~ICL; //complement 
assign icm = ~ICM; //complement 
assign icn = ~ICN; //complement 
assign ico = ~ICO; //complement 
assign icp = ~ICP; //complement 
assign ida = ~IDA; //complement 
assign idb = ~IDB; //complement 
assign idc = ~IDC; //complement 
assign idd = ~IDD; //complement 
assign ide = ~IDE; //complement 
assign idf = ~IDF; //complement 
assign idg = ~IDG; //complement 
assign idh = ~IDH; //complement 
assign idi = ~IDI; //complement 
assign idj = ~IDJ; //complement 
assign idk = ~IDK; //complement 
assign idl = ~IDL; //complement 
assign idm = ~IDM; //complement 
assign idn = ~IDN; //complement 
assign ido = ~IDO; //complement 
assign idp = ~IDP; //complement 
assign iea = ~IEA; //complement 
assign ieb = ~IEB; //complement 
assign iec = ~IEC; //complement 
assign ied = ~IED; //complement 
assign iee = ~IEE; //complement 
assign ief = ~IEF; //complement 
assign ieg = ~IEG; //complement 
assign ieh = ~IEH; //complement 
assign iei = ~IEI; //complement 
assign iej = ~IEJ; //complement 
assign iek = ~IEK; //complement 
assign iel = ~IEL; //complement 
assign iem = ~IEM; //complement 
assign ien = ~IEN; //complement 
assign ieo = ~IEO; //complement 
assign iep = ~IEP; //complement 
assign ifa = ~IFA; //complement 
assign ifb = ~IFB; //complement 
assign ifc = ~IFC; //complement 
assign ifd = ~IFD; //complement 
assign ife = ~IFE; //complement 
assign ifff  = ~IFFF ; //complement 
assign ifg = ~IFG; //complement 
assign ifh = ~IFH; //complement 
assign ifi = ~IFI; //complement 
assign ifj = ~IFJ; //complement 
assign ifk = ~IFK; //complement 
assign ifl = ~IFL; //complement 
assign ifm = ~IFM; //complement 
assign ifn = ~IFN; //complement 
assign ifo = ~IFO; //complement 
assign ifp = ~IFP; //complement 
assign iga = ~IGA; //complement 
assign igb = ~IGB; //complement 
assign igc = ~IGC; //complement 
assign igd = ~IGD; //complement 
assign ige = ~IGE; //complement 
assign igf = ~IGF; //complement 
assign igg = ~IGG; //complement 
assign igh = ~IGH; //complement 
assign igi = ~IGI; //complement 
assign igj = ~IGJ; //complement 
assign igk = ~IGK; //complement 
assign igl = ~IGL; //complement 
assign igm = ~IGM; //complement 
assign ign = ~IGN; //complement 
assign igo = ~IGO; //complement 
assign igp = ~IGP; //complement 
assign iha = ~IHA; //complement 
assign ihb = ~IHB; //complement 
assign iia = ~IIA; //complement 
assign iib = ~IIB; //complement 
assign ija = ~IJA; //complement 
assign ijb = ~IJB; //complement 
assign ijc = ~IJC; //complement 
assign ijd = ~IJD; //complement 
always@(posedge IZZ )
   begin 
 BEA <=  BEA & tca & tda  |  NAA & TCA  |  IAA & TDA  ; 
 BEB <=  BEB & tca & tda  |  NAB & TCA  |  IAB & TDA  ; 
 BAB <=  BAB & taa & tba  |  NAB & TAA  |  IAB & TBA  ; 
 BAA <=  BAA & taa & tba  |  NAA & TAA  |  IAA & TBA  ; 
 BEC <=  BEC & tca & tda  |  NAC & TCA  |  IAC & TDA  ; 
 BED <=  BED & tca & tda  |  NAD & TCA  |  IAD & TDA  ; 
 BAC <=  BAC & taa & tba  |  NAC & TAA  |  IAC & TBA  ; 
 BAD <=  BAD & taa & tba  |  NAD & TAA  |  IAD & TBA  ; 
 BEE <=  BEE & tca & tda  |  NAE & TCA  |  IAE & TDA  ; 
 BEF <=  BEF & tca & tda  |  NAF & TCA  |  IAF & TDA  ; 
 BAE <=  BAE & taa & tba  |  NAE & TAA  |  IAE & TBA  ; 
 BAF <=  BAF & taa & tba  |  NAF & TAA  |  IAF & TBA  ; 
 BEG <=  BEG & tca & tda  |  NAG & TCA  |  IAG & TDA  ; 
 BEH <=  BEH & tca & tda  |  NAH & TCA  |  IAH & TDA  ; 
 WAE <= PEA ; 
 WAF <= PEA ; 
 WAG <= PEA ; 
 WAH <= PEA ; 
 BHJ <=  BHJ & tcd & tdd  |  NDJ & TCD  |  IDJ & TDD  ; 
 BHK <=  BHK & tcd & tdd  |  NDK & TCD  |  IDK & TDD  ; 
 BHL <=  BHL & tcd & tdd  |  NDL & TCD  |  IDL & TDD  ; 
 BAG <=  BAG & taa & tba  |  NAG & TAA  |  IAG & TBA  ; 
 BAH <=  BAH & taa & tba  |  NAH & TAA  |  IAH & TBA  ; 
 BHM <=  BHM & tcd & tdd  |  NDM & TCD  |  IDM & TDD  ; 
 BHN <=  BHN & tcd & tdd  |  NDN & TCD  |  IDN & TDD  ; 
 BHO <=  BHO & tcd & tdd  |  NDO & TCD  |  IDO & TDD  ; 
 BHP <=  BHP & tcd & tdd  |  NDP & TCD  |  IDP & TDD  ; 
 AAA <=  GAA & TMA  |  IEC & TNA  |  KAC & TOA  ; 
 AAB <=  GAB & TMA  |  IED & TNA  |  KAD & TOA  ; 
 AAC <=  GAC & TMA  |  IEE & TNA  |  KAE & TOA  ; 
 AAD <=  GAD & TMA  |  IEF & TNA  |  KAF & TOA  ; 
 AAE <=  GAE & TMA  |  IEG & TNA  |  KAG & TOA  ; 
 AAF <=  GAF & TMA  |  IEH & TNA  |  KAH & TOA  ; 
 AAG <=  GAG & TMA  |  IEI & TNA  |  KAI & TOA  ; 
 AAH <=  GAH & TMA  |  IEJ & TNA  |  KAJ & TOA  ; 
 AAI <=  GAI & TMB  |  IEK & TNB  |  KAK & TOB  ; 
 AAJ <=  GAJ & TMB  |  IEL & TNB  |  KAL & TOB  ; 
 AAK <=  GAK & TMB  |  IEM & TNB  |  KAM & TOB  ; 
 AAL <=  GAL & TMB  |  IEN & TNB  |  KAN & TOB  ; 
 MAA <=  BAA & bab & bac  |  baa & BAB & bac  |  baa & bab & BAC  |  BAA & BAB & BAC  ;
 WAA <= PEA ; 
 WAB <= PEA ; 
 WAC <= PEA ; 
 WAD <= PEA ; 
 wai <= pea ; 
 waj <= pea ; 
 wak <= pea ; 
 wal <= pea ; 
 wam <= pea ; 
 wan <= pea ; 
 wao <= pea ; 
 wap <= pea ; 
 BEP <=  BEP & tcb & tdb  |  NAP & TCB  |  IAP & TDB  ; 
 TGA <= PCC ; 
 TGB <= PCC ; 
 TGC <= PCC ; 
 TGD <= PCC ; 
 FAA <= ABA ; 
 FAB <= ABB ; 
 FAC <= ABC ; 
 FAD <= ABD ; 
 FAE <= ABE ; 
 FAF <= ABF ; 
 FAG <= ABG ; 
 FAH <= ABH ; 
 FAI <= ABI ; 
 FAJ <= ABJ ; 
 FAK <= ABK ; 
 FAL <= ABL ; 
 NAI <= IEI ; 
 NAJ <= IEJ ; 
 NAK <= IEK ; 
 NAL <= IEL ; 
 OAA <=  SAA & TEA  |  SEA & TFA  |  SIA & TGA  |  SMA & THA  ; 
 NAM <= IEM ; 
 NAN <= IEN ; 
 NAO <= IEO ; 
 NAP <= IEP ; 
 OAB <=  SAB & TEB  |  SEB & TFB  |  SIB & TGB  |  SMB & THB  ; 
 QAC <= QAB ; 
 QBD <= IJB ; 
 QBB <= IJB ; 
 QBC <= IJC ; 
 OAC <=  SAC & TEA  |  SEC & TFA  |  SIC & TGA  |  SMC & THA  ; 
 OAD <=  SAD & TEB  |  SED & TFB  |  SID & TGB  |  SMD & THB  ; 
 KAC <= IGC ; 
 KAD <= IGD ; 
 OAE <=  SAE & TEC  |  SEE & TFC  |  SIE & TGC  |  SME & THC  ; 
 OAF <=  SAF & TED  |  SEF & TFD  |  SIF & TGD  |  SMF & THD  ; 
 twk <= pcc ; 
 twl <= pcc ; 
 twm <= pcc ; 
 twn <= pcc ; 
 KAE <= IGE ; 
 KAF <= IGF ; 
 KAG <= IGG ; 
 KAH <= IGH ; 
 NAA <= IEA ; 
 NAB <= IEB ; 
 NAC <= IEC ; 
 NAD <= IED ; 
 KAI <= IGI ; 
 KAJ <= IGJ ; 
 KAK <= IGK ; 
 KAL <= IGL ; 
 OAG <=  SAG & TEC  |  SEG & TFC  |  SIG & TGC  |  SMG & THC  ; 
 KAM <= IGM ; 
 KAN <= IGN ; 
 KAO <= IGO ; 
 KAP <= IGP ; 
 OAH <=  SAH & TED  |  SEH & TFD  |  SIH & TGD  |  SMH & THD  ; 
 NAE <= IEE ; 
 NAF <= IEF ; 
 NAG <= IEG ; 
 NAH <= IEH ; 
 BEI <=  BEI & tcb & tdb  |  NAI & TCB  |  IAI & TDB  ; 
 BEJ <=  BEJ & tcb & tdb  |  NAJ & TCB  |  IAJ & TDB  ; 
 BAI <=  BAI & tab & tbb  |  NAI & TAB  |  IAI & TBB  ; 
 BAJ <=  BAJ & tab & tbb  |  NAJ & TAB  |  IAJ & TBB  ; 
 BEK <=  BEK & tcb & tdb  |  NAK & TCB  |  IAK & TDB  ; 
 BEL <=  BEL & tcb & tdb  |  NAL & TCB  |  IAL & TDB  ; 
 BAK <=  BAK & tab & tbb  |  NAK & TAB  |  IAK & TBB  ; 
 BAL <=  BAL & tab & tbb  |  NAL & TAB  |  IAL & TBB  ; 
 BEM <=  BEM & tcb & tdb  |  NAM & TCB  |  IAM & TDB  ; 
 BEN <=  BEN & tcb & tdb  |  NAN & TCB  |  IAN & TDB  ; 
 BAM <=  BAM & tab & tbb  |  NAM & TAB  |  IAM & TBB  ; 
 BAN <=  BAN & tab & tbb  |  NAN & TAB  |  IAN & TBB  ; 
 BEO <=  BEO & tcb & tdb  |  NAO & TCB  |  IAO & TDB  ; 
 BAO <=  BAO & tab & tbb  |  NAO & TAB  |  IAO & TBB  ; 
 BAP <=  BAP & tab & tbb  |  NAP & TAB  |  IAP & TBB  ; 
 BHA <=  BHA & tcc & tdc  |  NDC & TCC  |  IDC & TDC  ; 
 BHB <=  BHB & tcc & tdc  |  NDB & TCC  |  IDB & TDC  ; 
 BHC <=  BHC & tcc & tdc  |  NDC & TCC  |  IDC & TDC  ; 
 BHD <=  BHD & tcc & tdc  |  NDD & TCC  |  IDD & TDC  ; 
 BHE <=  BHE & tcc & tdc  |  NDE & TCC  |  IDE & TDC  ; 
 BHF <=  BHF & tcc & tdc  |  NDF & TCC  |  IDF & TDC  ; 
 BHG <=  BHG & tcc & tdc  |  NDG & TCC  |  IDG & TDC  ; 
 BHH <=  BHH & tcc & tdc  |  NDH & TCC  |  IDH & TDC  ; 
 BHI <=  BHI & tcd & tdd  |  NDI & TCD  |  IDI & TDD  ; 
 ABA <=  AEA & TMC  |  IEC & TNC  |  KAC & TOC  ; 
 ABB <=  AEB & TMC  |  IED & TNC  |  KAD & TOC  ; 
 ABC <=  AEC & TMC  |  IEE & TNC  |  KAE & TOC  ; 
 ABD <=  AED & TMC  |  IEF & TNC  |  KAF & TOC  ; 
 ABE <=  AEE & TMC  |  IEG & TNC  |  KAG & TOC  ; 
 ABF <=  AEF & TMC  |  IEH & TNC  |  KAH & TOC  ; 
 ABG <=  AEG & TMC  |  IEI & TNC  |  KAI & TOC  ; 
 ABH <=  AEH & TMC  |  IEJ & TNC  |  KAJ & TOC  ; 
 ABI <=  AEI & TMD  |  IEK & TND  |  KAK & TOD  ; 
 ABJ <=  AEJ & TMD  |  IEL & TND  |  KAL & TOD  ; 
 ABK <=  AEK & TMD  |  IEM & TND  |  KAM & TOD  ; 
 ABL <=  AEL & TMD  |  IEN & TND  |  KAN & TOD  ; 
 KAA <= IGA & tla |  KAA & TLA ; 
 KAB <= IGB & tla |  KAB & TLA ; 
 TGE <= PCC ; 
 TGF <= PCC ; 
 TGG <= PCC ; 
 TGH <= PCC ; 
 PCA <= PBA ; 
 PCB <= PBB ; 
 PCC <= PBC ; 
 PCD <= PBD ; 
 PCE <= PBA ; 
 PCF <= PBB ; 
 PCG <= PBC ; 
 PCH <= PBD ; 
 PDA <= QBD & PAA ; 
 PDB <= QBD & PAB ; 
 PDC <= QBD & PAC ; 
 PDD <= QBD & PAD ; 
 FBB <= aba & ABB |  ABA & abb ; 
 FBF <= abe & ABF |  ABE & abf ; 
 FBJ <= abi & ABJ |  ABI & abj ; 
 FBA <= aba ; 
 FBE <= abe ; 
 FBI <= abi ; 
 PBA <= PAA ; 
 PBB <= PAB ; 
 PBC <= PAC ; 
 PBD <= PAD ; 
 OAI <=  SAI & TEE  |  SEI & TFE  |  SII & TGE  |  SMI & THE  ; 
 GAK <= FAK & fbp |  FBK & FBP ; 
 GAL <= FAL & fbp |  FBL & FBP ; 
 OAJ <=  SAJ & TEF  |  SEJ & TFF  |  SIJ & TGF  |  SMJ & THF  ; 
 NBA <= IFA ; 
 NBB <= IFB ; 
 NBC <= IFC ; 
 NBD <= IFD ; 
 NBE <= IFE ; 
 NBF <= IFFF  ; 
 NBG <= IFG ; 
 NBH <= IFH ; 
 OAK <=  SAK & TEE  |  SEK & TFE  |  SIK & TGE  |  SMK & THE  ; 
 NBI <= IFI ; 
 NBJ <= IFJ ; 
 NBK <= IFK ; 
 NBL <= IFL ; 
 NBM <= IFM ; 
 NBN <= IFN ; 
 NBO <= IFO ; 
 NBP <= IFP ; 
 OAL <=  SAL & TEF  |  SEL & TFF  |  SIL & TGF  |  SML & THF  ; 
 OAM <=  SAM & TEG  |  SEM & TFG  |  SIM & TGG  |  SMM & THG  ; 
 wbi <= peb ; 
 wbj <= peb ; 
 wbk <= peb ; 
 wbl <= peb ; 
 wbm <= peb ; 
 wbn <= peb ; 
 wbo <= peb ; 
 wbp <= peb ; 
 OAN <=  SAN & TEH  |  SEN & TFH  |  SIN & TGH  |  SMN & THH  ; 
 WBA <= PEB ; 
 WBB <= PEB ; 
 WBC <= PEB ; 
 WBD <= PEB ; 
 WBE <= PEB ; 
 WBF <= PEB ; 
 WBG <= PEB ; 
 WBH <= PEB ; 
 OAO <=  SAO & TEG  |  SEO & TFG  |  SIO & TGG  |  SMO & THG  ; 
 GAA <= FBA ; 
 GAB <= FBB ; 
 GAC <= FBC ; 
 GAD <= FBD ; 
 GAE <= FAE & fbo |  FBE & FBO ; 
 GAF <= FAF & fbo |  FBF & FBO ; 
 OAP <=  SAP & TEH  |  SEP & TFH  |  SIP & TGH  |  SMP & THH  ; 
 GAG <= FAG & fbo |  FBG & FBO ; 
 GAH <= FAH & fbo |  FBH & FBO ; 
 GAI <= FAI & fbp |  FBI & FBP ; 
 GAJ <= FAJ & fbp |  FBJ & FBP ; 
 BFA <=  BFA & tca & tda  |  NBA & TCA  |  IBA & TDA  ; 
 BFB <=  BFB & tca & tda  |  NBB & TCA  |  IBB & TDA  ; 
 BBA <=  BBA & taa & tba  |  NBA & TAA  |  IBA & TBA  ; 
 BBB <=  BBB & taa & tba  |  NBB & TAA  |  IBB & TBA  ; 
 BFC <=  BFC & tca & tda  |  NBC & TCA  |  IBC & TDA  ; 
 BFD <=  BFD & tca & tda  |  NBD & TCA  |  IBD & TDA  ; 
 BBC <=  BBC & taa & tba  |  NBC & TAA  |  IBC & TBA  ; 
 BBD <=  BBD & taa & tba  |  NBD & TAA  |  IBD & TBA  ; 
 BFE <=  BFE & tca & tda  |  NBE & TCA  |  IBE & TDA  ; 
 BFF <=  BFF & tca & tda  |  NBF & TCA  |  IBF & TDA  ; 
 BBE <=  BBE & taa & tba  |  NBE & TAA  |  IBE & TBA  ; 
 BBF <=  BBF & taa & tba  |  NBF & TAA  |  IBF & TBA  ; 
 BFG <=  BFG & tca & tda  |  NBG & TCA  |  IBG & TDA  ; 
 BFH <=  BFH & tca & tda  |  NBH & TCA  |  IBH & TDA  ; 
 BBG <=  BBG & taa & tba  |  NBG & TAA  |  IBG & TBA  ; 
 BBH <=  BBH & taa & tba  |  NBH & TAA  |  IBH & TBA  ; 
 tgm <= pcc ; 
 tgn <= pcc ; 
 tgo <= pcc ; 
 tgp <= pcc ; 
 THA <= PCD ; 
 THB <= PCD ; 
 THC <= PCD ; 
 THD <= PCD ; 
 PEA <=  PDA  |  PAA & QBD  ; 
 PEB <=  PDB  |  PAB & QBD  ; 
 PEC <=  PDC  |  PAC & QBD  ; 
 PED <=  PDD  |  PAD & QBD  ; 
 THE <= PCD ; 
 THF <= PCD ; 
 THG <= PCD ; 
 THH <= PCD ; 
 ACA <=  AFA & TME  |  IEC & TNE  |  KAC & TOE  ; 
 ACB <=  AFB & TME  |  IED & TNE  |  KAD & TOE  ; 
 ACC <=  AFC & TME  |  IEE & TNE  |  KAE & TOE  ; 
 ACD <=  AFD & TME  |  IEF & TNE  |  KAF & TOE  ; 
 ACE <=  AFE & TME  |  IEG & TNE  |  KAG & TOE  ; 
 ACF <=  AFF & TME  |  IEH & TNE  |  KAH & TOE  ; 
 ACG <=  AFG & TME  |  IEI & TNE  |  KAI & TOE  ; 
 ACH <=  AFH & TME  |  IEJ & TNE  |  KAJ & TOE  ; 
 ACI <=  AFI & TMF  |  IEK & TNF  |  KAK & TOF  ; 
 ACJ <=  AFJ & TMF  |  IEL & TNF  |  KAL & TOF  ; 
 ACK <=  AFK & TMF  |  IEM & TNF  |  KAM & TOF  ; 
 ACL <=  AFL & TMF  |  IEN & TNF  |  KAN & TOF  ; 
 MAB <=  BAD & bae & baf  |  bad & BAE & baf  |  bad & bae & BAF  |  BAD & BAE & BAF  ;
 TGI <= PCC ; 
 TGJ <= PCC ; 
 tgk <= pcc ; 
 tgl <= pcc ; 
 TFE <= PCB ; 
 TFF <= PCB ; 
 TFG <= PCB ; 
 TFH <= PCB ; 
 TFI <= PCB ; 
 TFJ <= PCB ; 
 tfk <= pcb ; 
 tfl <= pcb ; 
 tfm <= pcb ; 
 tfn <= pcb ; 
 tfo <= pcb ; 
 tfp <= pcb ; 
 thm <= pcd ; 
 thn <= pcd ; 
 tho <= pcd ; 
 thp <= pcd ; 
 JMA <=  MAA & mab & mac  |  maa & MAB & mac  |  maa & mab & MAC  |  MAA & MAB & MAC  ;
 THI <= PCD ; 
 THJ <= PCD ; 
 thk <= pcd ; 
 thl <= pcd ; 
 TFA <= PCB ; 
 TFB <= PCB ; 
 TFC <= PCB ; 
 TFD <= PCB ; 
 OBA <=  SBA & TEK  |  SFA & TFK  |  SJA & TGK  |  SNA & THK  ; 
 JMC <=  MAG & mah & mai  |  mag & MAH & mai  |  mag & mah & MAI  |  MAG & MAH & MAI  ;
 JMD <=  MAJ & mak & mal  |  maj & MAK & mal  |  maj & mak & MAL  |  MAJ & MAK & MAL  ;
 OBB <=  SBB & TEL  |  SFB & TFL  |  SJB & TGL  |  SNB & THL  ; 
 ndm <= ifp ; 
 ndn <= ifp ; 
 ndo <= ifp ; 
 ndp <= ifp ; 
 QDA <= IJD ; 
 QDB <= IJD ; 
 QDC <= QDB ; 
 QFA <= IJA ; 
 OBC <=  SBC & TEK  |  SFC & TFK  |  SJC & TGK  |  SNC & THK  ; 
 thq <= pcd ; 
 thr <= pcd ; 
 tgq <= pcc ; 
 tgr <= pcc ; 
 teq <= pca ; 
 ter <= pca ; 
 tfq <= pcb ; 
 tfr <= pcb ; 
 OBD <=  SBD & TEL  |  SFD & TFL  |  SJD & TGL  |  SND & THL  ; 
 TMA <= qaa & PCE ; 
 TMB <= qaa & PCE ; 
 TMC <= qaa & qfa ; 
 TMD <= qaa & qfa ; 
 TME <= qaa & qfa ; 
 TMF <= qaa & qfa ; 
 TMG <= qaa & qfa ; 
 TMH <= qaa & qfa ; 
 OBE <=  SBE & TEM  |  SFE & TFM  |  SJE & TGM  |  SNE & THM  ; 
 OBF <=  SBF & TEN  |  SFF & TFN  |  SJF & TGN  |  SNF & THM  ; 
 OBG <=  SBG & TEM  |  SFG & TFM  |  SJG & TGM  |  SNG & THM  ; 
 PAA <=  JCA  |  JDA  |  JEA  ; 
 JMB <=  MAD & mae & maf  |  mad & MAE & maf  |  mad & mae & MAF  |  MAD & MAE & MAF  ;
 OBI <=  SBI & TEO  |  SFI & TFO  |  SJI & TGO  |  SNI & THO  ; 
 NDA <= IFP ; 
 NDB <= IFP ; 
 NDC <= IFP ; 
 NDD <= IFP ; 
 NDE <= IFP ; 
 NDF <= IFP ; 
 NDG <= IFP ; 
 NDH <= IFP ; 
 OBH <=  SBH & TEN  |  SFH & TFN  |  SJH & TGN  |  SNH & THN  ; 
 ndi <= ifp ; 
 ndj <= ifp ; 
 ndk <= ifp ; 
 ndl <= ifp ; 
 BFI <=  BFI & tcb & tdb  |  NBI & TCB  |  IBI & TDB  ; 
 BFJ <=  BFJ & tcb & tdb  |  NBJ & TCB  |  IBJ & TDB  ; 
 BBI <=  BBI & tab & tbb  |  NBI & TAB  |  IBI & TBB  ; 
 BBJ <=  BBJ & tab & tbb  |  NBJ & TAB  |  IBJ & TBB  ; 
 BFK <=  BFK & tcb & tdb  |  NBK & TCB  |  IBK & TDB  ; 
 BFL <=  BFL & tcb & tdb  |  NBL & TCB  |  IBL & TDB  ; 
 BBK <=  BBK & tab & tbb  |  NBK & TAB  |  IBK & TBB  ; 
 BBL <=  BBL & tab & tbb  |  NBL & TAB  |  IBL & TBB  ; 
 BFM <=  BFM & tcb & tdb  |  NBM & TCB  |  IBM & TDB  ; 
 BFN <=  BFN & tcb & tdb  |  NBN & TCB  |  IBN & TDB  ; 
 BBM <=  BBM & tab & tbb  |  NBM & TAB  |  IBM & TBB  ; 
 BBN <=  BBN & tab & tbb  |  NBN & TAB  |  IBN & TBB  ; 
 BFO <=  BFO & tcb & tdb  |  NBO & TCB  |  IBO & TDB  ; 
 BFP <=  BFP & tcb & tdb  |  NBP & TCB  |  IBP & TDB  ; 
 BBO <=  BBO & tab & tbb  |  NBO & TAB  |  IBO & TBB  ; 
 BBP <=  BBP & tab & tbb  |  NBP & TAB  |  IBP & TBB  ; 
 tum <= pca ; 
 tun <= pca ; 
 tuo <= pca ; 
 tup <= pca ; 
 TVA <= PCB ; 
 TVB <= PCB ; 
 TVC <= PCB ; 
 TVD <= PCB ; 
 PAC <=  JCC  |  JDC  |  JEC  ; 
 PAD <=  JCD  |  JDD  |  JED  ; 
 TUA <= PCA ; 
 TUB <= PCA ; 
 TUC <= PCA ; 
 TUD <= PCA ; 
 TVE <= PCB ; 
 TVF <= PCB ; 
 TVG <= PCB ; 
 TVH <= PCB ; 
 TUE <= PCA ; 
 TUF <= PCA ; 
 TUG <= PCA ; 
 TUH <= PCA ; 
 TUI <= PCA ; 
 TUJ <= PCA ; 
 tuk <= pca ; 
 tul <= pca ; 
 ADA <=  AGA & TMG  |  IEC & TNG  |  KAC & TOG  ; 
 ADB <=  AGB & TMG  |  IED & TNG  |  KAD & TOG  ; 
 ADC <=  AGC & TMG  |  IEE & TNG  |  KAE & TOG  ; 
 ADD <=  AGD & TMG  |  IEF & TNG  |  KAF & TOG  ; 
 ADE <=  AGE & TMG  |  IEG & TNG  |  KAG & TOG  ; 
 ADF <=  AGF & TMG  |  IEH & TNG  |  KAH & TOG  ; 
 ADG <=  AGG & TMG  |  IEI & TNG  |  KAI & TOG  ; 
 ADH <=  AGH & TMG  |  IEJ & TNG  |  KAJ & TOG  ; 
 ADI <=  AGI & TMH  |  IEK & TNH  |  KAK & TOH  ; 
 ADJ <=  AGJ & TMH  |  IEL & TNH  |  KAL & TOH  ; 
 ADK <=  AGK & TMH  |  IEM & TNH  |  KAM & TOH  ; 
 ADL <=  AGL & TMH  |  IEN & TNH  |  KAN & TOH  ; 
 txk <= pcd ; 
 txl <= pcd ; 
 txm <= pcd ; 
 txn <= pcd ; 
 PAB <=  JCB  |  JDB  |  JEB  ; 
 OBJ <=  SBJ & TEP  |  SFJ & TFP  |  SJJ & TGP  |  SNJ & THP  ; 
 OED <=  SCD & TUB  |  SGD & TVB  |  SKD & TWB  |  SOD & TXB  ; 
 OEE <=  SCE & TUC  |  SGE & TVC  |  SKE & TWC  |  SOE & TXC  ; 
 OEF <=  SCF & TUD  |  SGF & TVD  |  SKF & TWD  |  SOF & TXD  ; 
 OBK <=  SBK & TEO  |  SFK & TFO  |  SJK & TGO  |  SNK & THO  ; 
 OEG <=  SCG & TUC  |  SGG & TVC  |  SKG & TWC  |  SOG & TXC  ; 
 OEH <=  SCH & TUD  |  SGH & TVD  |  SKH & TWD  |  SOH & TXD  ; 
 QAA <=  IIA & IHA & IHB  |  QAC  ; 
 OBL <=  SBL & TEP  |  SFL & TFP  |  SJL & TGP  |  SNL & THP  ; 
 NCA <= IFP ; 
 NCB <= IFP ; 
 NCC <= IFP ; 
 NCD <= IFP ; 
 NCE <= IFP ; 
 NCF <= IFP ; 
 NCG <= IFP ; 
 NCH <= IFP ; 
 nci <= ifp ; 
 ncj <= ifp ; 
 nck <= ifp ; 
 ncl <= ifp ; 
 OBM <=  SBM & TEQ  |  SFM & TFQ  |  SJM & TGQ  |  SNM & THQ  ; 
 ncm <= ifp ; 
 ncn <= ifp ; 
 nco <= ifp ; 
 ncp <= ifp ; 
 QAB <=  IIB & IHA & IHB  ; 
 TEA <= PCA ; 
 TEB <= PCA ; 
 TEC <= PCA ; 
 TED <= PCA ; 
 OBN <=  SBN & TER  |  SFN & TFR  |  SJN & TGR  |  SNN & THR  ; 
 WCA <= PEC ; 
 WCB <= PEC ; 
 WCC <= PEC ; 
 WCD <= PEC ; 
 WCE <= PEC ; 
 WCF <= PEC ; 
 WCG <= PEC ; 
 WCH <= PEC ; 
 wci <= pec ; 
 wcj <= pec ; 
 wck <= pec ; 
 wcl <= pec ; 
 wcm <= pec ; 
 wcn <= pec ; 
 wco <= pec ; 
 wcp <= pec ; 
 OBO <=  SBO & TEQ  |  SFO & TFQ  |  SJO & TGQ  |  SNO & THQ  ; 
 TWA <= PCC ; 
 TWB <= PCC ; 
 TWC <= PCC ; 
 TWD <= PCC ; 
 TWE <= PCC ; 
 TWF <= PCC ; 
 TWG <= PCC ; 
 TWH <= PCC ; 
 OBP <=  SBP & TER  |  SFP & TFR  |  SJP & TGR  |  SNP & THR  ; 
 OEA <=  SCA & TUA  |  SGA & TVA  |  SKA & TWA  |  SOA & TXA  ; 
 OEB <=  SCB & TUB  |  SGB & TVB  |  SKB & TWB  |  SOB & TXB  ; 
 TWI <= PCC ; 
 TWJ <= PCC ; 
 OEC <=  SCC & TUA  |  SGC & TVA  |  SKC & TWA  |  SOC & TXA  ; 
 BGA <=  BGA & tcc & tdc  |  NCC & TCC  |  ICC & TDC  ; 
 BGB <=  BGB & tcc & tdc  |  NCB & TCC  |  ICB & TDC  ; 
 BCA <=  BCA & tac & tbc  |  NCC & TAC  |  ICC & TBC  ; 
 BCB <=  BCB & tac & tbc  |  NCB & TAC  |  ICB & TBC  ; 
 BGC <=  BGC & tcc & tdc  |  NCC & TCC  |  ICC & TDC  ; 
 BGD <=  BGD & tcc & tdc  |  NCD & TCC  |  ICD & TDC  ; 
 BCC <=  BCC & tac & tbc  |  NCC & TAC  |  ICC & TBC  ; 
 BCD <=  BCD & tac & tbc  |  NCD & TAC  |  ICD & TBC  ; 
 BGE <=  BGE & tcc & tdc  |  NCE & TCC  |  ICE & TDC  ; 
 BGF <=  BGF & tcc & tdc  |  NCF & TCC  |  ICF & TDC  ; 
 BCE <=  BCE & tac & tbc  |  NCE & TAC  |  ICE & TBC  ; 
 BCF <=  BCF & tac & tbc  |  NCF & TAC  |  ICF & TBC  ; 
 BGG <=  BGG & tcc & tdc  |  NCG & TCC  |  ICG & TDC  ; 
 BGH <=  BGH & tcc & tdc  |  NCH & TCC  |  ICH & TDC  ; 
 BCG <=  BCG & tac & tbc  |  NCG & TAC  |  ICG & TBC  ; 
 BCH <=  BCH & tac & tbc  |  NCH & TAC  |  ICH & TBC  ; 
 TEI <= PCA ; 
 TEJ <= PCA ; 
 tek <= pca ; 
 tel <= pca ; 
 tem <= pca ; 
 ten <= pca ; 
 teo <= pca ; 
 tep <= pca ; 
 JME <=  MAM & man & mao  |  mam & MAN & mao  |  mam & man & MAO  |  MAM & MAN & MAO  ;
 WDA <= PED ; 
 WDB <= PED ; 
 WDC <= PED ; 
 WDD <= PED ; 
 WDE <= PED ; 
 WDF <= PED ; 
 WDG <= PED ; 
 WDH <= PED ; 
 wdi <= ped ; 
 wdj <= ped ; 
 wdk <= ped ; 
 wdl <= ped ; 
 AEA <=  GAA & TMA  |  IEC & TNA  |  KAC & TOA  ; 
 AEB <=  GAB & TMA  |  IED & TNA  |  KAD & TOA  ; 
 AEC <=  GAC & TMA  |  IEE & TNA  |  KAE & TOA  ; 
 AED <=  GAD & TMA  |  IEF & TNA  |  KAF & TOA  ; 
 AEE <=  GAE & TMA  |  IEG & TNA  |  KAG & TOA  ; 
 AEF <=  GAF & TMA  |  IEH & TNA  |  KAH & TOA  ; 
 AEG <=  GAG & TMA  |  IEI & TNA  |  KAI & TOA  ; 
 AEH <=  GAH & TMA  |  IEJ & TNA  |  KAJ & TOA  ; 
 AEI <=  GAI & TMB  |  IEK & TNB  |  KAK & TOB  ; 
 AEJ <=  GAJ & TMB  |  IEL & TNB  |  KAL & TOB  ; 
 AEK <=  GAK & TMB  |  IEM & TNB  |  KAM & TOB  ; 
 AEL <=  GAL & TMB  |  IEN & TNB  |  KAN & TOB  ; 
 txo <= pcd ; 
 txp <= pcd ; 
 txq <= pcd ; 
 txr <= pcd ; 
 TEE <= PCA ; 
 TEF <= PCA ; 
 TEG <= PCA ; 
 TEH <= PCA ; 
 OCA <=  SCA & TEA  |  SGA & TFA  |  SKA & TGA  |  SOA & THA  ; 
 TVI <= PCB ; 
 TVJ <= PCB ; 
 tvk <= pcb ; 
 tvl <= pcb ; 
 TXI <= PCD ; 
 TXJ <= PCD ; 
 OCB <=  SCB & TEB  |  SGB & TFB  |  SKB & TGB  |  SOB & THB  ; 
 OCC <=  SCC & TEA  |  SGC & TFA  |  SKC & TGA  |  SOC & THA  ; 
 tvm <= pcb ; 
 tvn <= pcb ; 
 tvo <= pcb ; 
 tvp <= pcb ; 
 tuq <= pca ; 
 tur <= pca ; 
 OCD <=  SCD & TEB  |  SGD & TFB  |  SKD & TGB  |  SOD & THB  ; 
 tvq <= pcb ; 
 tvr <= pcb ; 
 two <= pcc ; 
 twp <= pcc ; 
 twq <= pcc ; 
 twr <= pcc ; 
 OCE <=  SCE & TEC  |  SGE & TFC  |  SKE & TGC  |  SOE & THC  ; 
 OCF <=  SCF & TED  |  SGF & TFD  |  SKF & TGD  |  SOF & THD  ; 
 OEI <=  SCI & TUE  |  SGI & TVE  |  SKI & TWE  |  SOI & TXE  ; 
 OEJ <=  SCJ & TUF  |  SGJ & TVF  |  SKJ & TWF  |  SOJ & TXF  ; 
 OCG <=  SCG & TEC  |  SGG & TFC  |  SKG & TGC  |  SOG & THC  ; 
 wdm <= ped ; 
 wdn <= ped ; 
 wdo <= ped ; 
 wdp <= ped ; 
 TXA <= PCD ; 
 TXB <= PCD ; 
 TXC <= PCD ; 
 TXD <= PCD ; 
 OCH <=  SCH & TED  |  SGH & TFD  |  SKH & TGD  |  SOH & THD  ; 
 TXE <= PCD ; 
 TXF <= PCD ; 
 TXG <= PCD ; 
 TXH <= PCD ; 
 BGI <=  BGI & tcd & tdd  |  NCI & TCD  |  ICI & TDD  ; 
 BGJ <=  BGJ & tcd & tdd  |  NCJ & TCD  |  ICJ & TDD  ; 
 BCI <=  BCI & tad & tbd  |  NCI & TAD  |  ICI & TBD  ; 
 BCJ <=  BCJ & tad & tbd  |  NCJ & TAD  |  ICJ & TBD  ; 
 BGK <=  BGK & tcd & tdd  |  NCK & TCD  |  ICK & TDD  ; 
 BGL <=  BGL & tcd & tdd  |  NCL & TCD  |  ICL & TDD  ; 
 BCK <=  BCK & tad & tbd  |  NCK & TAD  |  ICK & TBD  ; 
 BCL <=  BCL & tad & tbd  |  NCL & TAD  |  ICL & TBD  ; 
 BGM <=  BGM & tcd & tdd  |  NCM & TCD  |  ICM & TDD  ; 
 BGN <=  BGN & tcd & tdd  |  NCN & TCD  |  ICN & TDD  ; 
 BCM <=  BCM & tad & tbd  |  NCM & TAD  |  ICM & TBD  ; 
 BCN <=  BCN & tad & tbd  |  NCN & TAD  |  ICN & TBD  ; 
 BGO <=  BGO & tcd & tdd  |  NCO & TCD  |  ICO & TDD  ; 
 BGP <=  BGP & tcd & tdd  |  NCP & TCD  |  ICP & TDD  ; 
 BCO <=  BCO & tad & tbd  |  NCO & TAD  |  ICO & TBD  ; 
 BCP <=  BCP & tad & tbd  |  NCP & TAD  |  ICP & TBD  ; 
 AFE <=  AEE & TMC  |  IEG & TNC  |  KAG & TOC  ; 
 AFF <=  AEF & TMC  |  IEH & TNC  |  KAH & TOC  ; 
 AFG <=  AEG & TMC  |  IEI & TNC  |  KAI & TOC  ; 
 AFH <=  AEH & TMC  |  IEJ & TNC  |  KAJ & TOC  ; 
 AFI <=  AEI & TMD  |  IEK & TND  |  KAK & TOD  ; 
 AFJ <=  AEJ & TMD  |  IEL & TND  |  KAL & TOD  ; 
 AFK <=  AEK & TMD  |  IEM & TND  |  KAM & TOD  ; 
 AFL <=  AEL & TMD  |  IEN & TND  |  KAN & TOD  ; 
 OEK <=  SCK & TUE  |  SGK & TVE  |  SKK & TWE  |  SOK & TXE  ; 
 AFA <=  AEA & TMC  |  IEC & TNC  |  KAC & TOC  ; 
 AFB <=  AEB & TMC  |  IED & TNC  |  KAD & TOC  ; 
 OEL <=  SCL & TUF  |  SGL & TVF  |  SKL & TWF  |  SOL & TXF  ; 
 OEM <=  SCM & TUG  |  SGM & TVG  |  SKM & TWG  |  SOM & TXG  ; 
 OEN <=  SCN & TUH  |  SGN & TVH  |  SKN & TWH  |  SON & TXH  ; 
 OEO <=  SCO & TUG  |  SGO & TVG  |  SKO & TWG  |  SOO & TXG  ; 
 OEP <=  SCP & TUH  |  SGP & TVH  |  SKP & TWH  |  SOP & TXH  ; 
 AFC <=  AEC & TMC  |  IEE & TNC  |  KAE & TOC  ; 
 AFD <=  AED & TMC  |  IEF & TNC  |  KAF & TOC  ; 
 OCI <=  SCI & TEE  |  SGI & TFE  |  SKI & TGE  |  SOI & THE  ; 
 OFF <=  SDF & TUN  |  SHF & TVN  |  SLF & TWN  |  SPF & TXM  ; 
 OFG <=  SDG & TUM  |  SHG & TVM  |  SLG & TWM  |  SPG & TXM  ; 
 OFH <=  SDH & TUN  |  SHH & TVN  |  SLH & TWN  |  SPH & TXN  ; 
 OCJ <=  SCJ & TEF  |  SGJ & TFF  |  SKJ & TGF  |  SOJ & THF  ; 
 FBG <=  ABE & ABF & abg  |  ABG & abe  |  ABG & abf  ; 
 FBK <=  ABI & ABJ & abk  |  ABK & abi  |  ABK & abj  ; 
 OCK <=  SCK & TEE  |  SGK & TFE  |  SKK & TGE  |  SOK & THE  ; 
 FBD <=  FAO & abd  |  ABD & aba  |  ABD & abb  |  ABD & abc  ; 
 OCL <=  SCL & TEF  |  SGL & TFF  |  SKL & TGF  |  SOL & THF  ; 
 FBH <=  FAP & abh  |  ABH & abe  |  ABH & abf  |  ABH & abg  ; 
 FBL <=  FAQ & abl  |  ABL & abi  |  ABL & abj  |  ABL & abk  ; 
 OCM <=  SCM & TEG  |  SGM & TFG  |  SKM & TGG  |  SOM & THG  ; 
 MAC <=  BAG & bah & bai  |  bag & BAH & bai  |  bag & bah & BAI  |  BAG & BAH & BAI  ;
 MAD <=  BAJ & bak & bal  |  baj & BAK & bal  |  baj & bak & BAL  |  BAJ & BAK & BAL  ;
 MAE <=  BAM & ban & bao  |  bam & BAN & bao  |  bam & ban & BAO  |  BAM & BAN & BAO  ;
 OCN <=  SCN & TEH  |  SGN & TFH  |  SKN & TGH  |  SON & THH  ; 
 MAF <=  BAP  |  BAP  ;
 MAG <=  BBA & bbb & bbc  |  bba & BBB & bbc  |  bba & bbb & BBC  |  BBA & BBB & BBC  ;
 MAH <=  BBD & bbe & bbf  |  bbd & BBE & bbf  |  bbd & bbe & BBF  |  BBD & BBE & BBF  ;
 OCO <=  SCO & TEG  |  SGO & TFG  |  SKO & TGG  |  SOO & THG  ; 
 OFA <=  SDA & TUK  |  SHA & TVK  |  SLA & TWK  |  SPA & TXK  ; 
 OFB <=  SDB & TUL  |  SHB & TVL  |  SLB & TWL  |  SPB & TXL  ; 
 OCP <=  SCP & TEH  |  SGP & TFH  |  SKP & TGH  |  SOP & THH  ; 
 OFC <=  SDC & TUK  |  SHC & TVK  |  SLC & TWK  |  SPC & TXK  ; 
 OFD <=  SDD & TUL  |  SHD & TVL  |  SLD & TWL  |  SPD & TXL  ; 
 OFE <=  SDE & TUM  |  SHE & TVM  |  SLE & TWM  |  SPE & TXM  ; 
 FBC <=  ABA & ABB & abc  |  ABC & aba  |  ABC & abb  ; 
 MAI <=  BBG & bbh & bbi  |  bbg & BBH & bbi  |  bbg & bbh & BBI  |  BBG & BBH & BBI  ;
 BDA <=  BDA & tac & tbc  |  NDC & TAC  |  IDC & TBC  ; 
 BDB <=  BDB & tac & tbc  |  NDB & TAC  |  IDB & TBC  ; 
 MAM <=  BCA & bcb & bcc  |  bca & BCB & bcc  |  bca & bcb & BCC  |  BCA & BCB & BCC  ;
 BDC <=  BDC & tac & tbc  |  NDC & TAC  |  IDC & TBC  ; 
 BDD <=  BDD & tac & tbc  |  NDD & TAC  |  IDD & TBC  ; 
 MAJ <=  BBJ & bbk & bbl  |  bbj & BBK & bbl  |  bbj & bbk & BBL  |  BBJ & BBK & BBL  ;
 BDE <=  BDE & tac & tbc  |  NDE & TAC  |  IDE & TBC  ; 
 BDF <=  BDF & tac & tbc  |  NDF & TAC  |  IDF & TBC  ; 
 BDG <=  BDG & tac & tbc  |  NDG & TAC  |  IDG & TBC  ; 
 BDH <=  BDH & tac & tbc  |  NDH & TAC  |  IDH & TBC  ; 
 MAK <=  BBM & bbn & bbo  |  bbm & BBN & bbo  |  bbm & bbn & BBO  |  BBM & BBN & BBO  ;
 MAL <=  BBP  |  BBP  ;
 MAN <=  BCD & bce & bcf  |  bcd & BCE & bcf  |  bcd & bce & BCF  |  BCD & BCE & BCF  ;
 MAO <=  BCG & bch & bci  |  bcg & BCH & bci  |  bcg & bch & BCI  |  BCG & BCH & BCI  ;
 MAP <=  BCJ & bck & bcl  |  bcj & BCK & bcl  |  bcj & bck & BCL  |  BCJ & BCK & BCL  ;
 AGA <=  AFA & TME  |  IEC & TNE  |  KAC & TOE  ; 
 AGB <=  AFB & TME  |  IED & TNE  |  KAD & TOE  ; 
 AGC <=  AFC & TME  |  IEE & TNE  |  KAE & TOE  ; 
 AGD <=  AFD & TME  |  IEF & TNE  |  KAF & TOE  ; 
 AGE <=  AFE & TME  |  IEG & TNE  |  KAG & TOE  ; 
 AGF <=  AFF & TME  |  IEH & TNE  |  KAH & TOE  ; 
 AGG <=  AFG & TME  |  IEI & TNE  |  KAI & TOE  ; 
 AGH <=  AFH & TME  |  IEJ & TNE  |  KAJ & TOE  ; 
 AGI <=  AFI & TMF  |  IEK & TNF  |  KAK & TOF  ; 
 AGJ <=  AFJ & TMF  |  IEL & TNF  |  KAL & TOF  ; 
 AGK <=  AFK & TMF  |  IEM & TNF  |  KAM & TOF  ; 
 AGL <=  AFL & TMF  |  IEN & TNF  |  KAN & TOF  ; 
 ODA <=  SDA & TEK  |  SHA & TFK  |  SLA & TGK  |  SPA & THK  ; 
 ODB <=  SDB & TEL  |  SHB & TFL  |  SLB & TGL  |  SPB & THL  ; 
 MAQ <=  BCM & bcn & bco  |  bcm & BCN & bco  |  bcm & bcn & BCO  |  BCM & BCN & BCO  ;
 ODC <=  SDC & TEK  |  SHC & TFK  |  SLC & TGK  |  SPC & THK  ; 
 MAR <=  BCP  |  BCP  ;
 MAS <=  BDA & bdb & bdc  |  bda & BDB & bdc  |  bda & bdb & BDC  |  BDA & BDB & BDC  ;
 ODD <=  SDD & TEL  |  SHD & TFL  |  SLD & TGL  |  SPD & THL  ; 
 ODE <=  SDE & TEM  |  SHE & TFM  |  SLE & TGM  |  SPE & THM  ; 
 MAT <=  BDD & bde & bdf  |  bdd & BDE & bdf  |  bdd & bde & BDF  |  BDD & BDE & BDF  ;
 ODF <=  SDF & TEN  |  SHF & TFN  |  SLF & TGN  |  SPF & THM  ; 
 MAU <=  BDG & bdh & bdi  |  bdg & BDH & bdi  |  bdg & bdh & BDI  |  BDG & BDH & BDI  ;
 MAV <=  BDJ & bdk & bdl  |  bdj & BDK & bdl  |  bdj & bdk & BDL  |  BDJ & BDK & BDL  ;
 ODG <=  SDG & TEM  |  SHG & TFM  |  SLG & TGM  |  SPG & THM  ; 
 OFI <=  SDI & TUO  |  SHI & TVO  |  SLI & TWO  |  SPI & TXO  ; 
 ODH <=  SDH & TEN  |  SHH & TFN  |  SLH & TGN  |  SPH & THN  ; 
 JMF <=  MAP & maq & mar  |  map & MAQ & mar  |  map & maq & MAR  |  MAP & MAQ & MAR  ;
 BDI <=  BDI & tad & tbd  |  NDI & TAD  |  IDI & TBD  ; 
 BDJ <=  BDJ & tad & tbd  |  NDJ & TAD  |  IDJ & TBD  ; 
 JMG <=  MAS & mat & mau  |  mas & MAT & mau  |  mas & mat & MAU  |  MAS & MAT & MAU  ;
 JMH <=  MAV & maw & max  |  mav & MAW & max  |  mav & maw & MAX  |  MAV & MAW & MAX  ;
 BDK <=  BDK & tad & tbd  |  NDK & TAD  |  IDK & TBD  ; 
 BDL <=  BDL & tad & tbd  |  NDL & TAD  |  IDL & TBD  ; 
 BDM <=  BDM & tad & tbd  |  NDM & TAD  |  IDM & TBD  ; 
 BDN <=  BDN & tad & tbd  |  NDN & TAD  |  IDN & TBD  ; 
 BDO <=  BDO & tad & tbd  |  NDO & TAD  |  IDO & TBD  ; 
 BDP <=  BDP & tad & tbd  |  NDP & TAD  |  IDP & TBD  ; 
 OHA <= JMA ; 
 OHB <= JMB ; 
 OHC <= JMC ; 
 OHD <= JMD ; 
 OHE <= JME ; 
 OHF <= JMF ; 
 OHG <= JMG ; 
 OHH <= JMH ; 
 AHA <=  AGA & TMG  |  IEC & TNG  |  KAC & TOG  ; 
 AHB <=  AGB & TMG  |  IED & TNG  |  KAD & TOG  ; 
 AHC <=  AGC & TMG  |  IEE & TNG  |  KAE & TOG  ; 
 AHD <=  AGD & TMG  |  IEF & TNG  |  KAF & TOG  ; 
 AHE <=  AGE & TMG  |  IEG & TNG  |  KAG & TOG  ; 
 AHF <=  AGF & TMG  |  IEH & TNG  |  KAH & TOG  ; 
 AHG <=  AGG & TMG  |  IEI & TNG  |  KAI & TOG  ; 
 AHH <=  AGH & TMG  |  IEJ & TNG  |  KAJ & TOG  ; 
 AHI <=  AGI & TMH  |  IEK & TNH  |  KAK & TOH  ; 
 AHJ <=  AGJ & TMH  |  IEL & TNH  |  KAL & TOH  ; 
 AHK <=  AGK & TMH  |  IEM & TNH  |  KAM & TOH  ; 
 AHL <=  AGL & TMH  |  IEN & TNH  |  KAN & TOH  ; 
 MAW <=  BDM & bdn & bdo  |  bdm & BDN & bdo  |  bdm & bdn & BDO  |  BDM & BDN & BDO  ;
 MAX <=  BDP  |  BDP  ;
 ODI <=  SDI & TEO  |  SHI & TFO  |  SLI & TGO  |  SPI & THO  ; 
 OFN <=  SDN & TUR  |  SHN & TVR  |  SLN & TWR  |  SPN & TXR  ; 
 OFO <=  SDO & TUQ  |  SHO & TVQ  |  SLO & TWQ  |  SPO & TXQ  ; 
 OFP <=  SDP & TUR  |  SHP & TVR  |  SLP & TWR  |  SPP & TXR  ; 
 ODJ <=  SDJ & TEP  |  SHJ & TFP  |  SLJ & TGP  |  SPJ & THP  ; 
 ODK <=  SDK & TEO  |  SHK & TFO  |  SLK & TGO  |  SPK & THO  ; 
 ODL <=  SDL & TEP  |  SHL & TFP  |  SLL & TGP  |  SPL & THP  ; 
 ODM <=  SDM & TEQ  |  SHM & TFQ  |  SLM & TGQ  |  SPM & THQ  ; 
 ODN <=  SDN & TER  |  SHN & TFR  |  SLN & TGR  |  SPN & THR  ; 
 ODO <=  SDO & TEQ  |  SHO & TFQ  |  SLO & TGQ  |  SPO & THQ  ; 
 OFJ <=  SDJ & TUP  |  SHJ & TVP  |  SLJ & TWP  |  SPJ & TXP  ; 
 OFK <=  SDK & TUO  |  SHK & TVO  |  SLK & TWO  |  SPK & TXO  ; 
 ODP <=  SDP & TER  |  SHP & TFR  |  SLP & TGR  |  SPP & THR  ; 
 OFL <=  SDL & TUP  |  SHL & TVP  |  SLL & TWP  |  SPL & TXP  ; 
 OFM <=  SDM & TUQ  |  SHM & TVQ  |  SLM & TWQ  |  SPM & TXQ  ; 
end
ram_4096x1 sinst_000(SAA,BAA,{AAA,AAB,AAC,AAD,AAE,AAF,AAG,AAH,AAI,AAJ,AAK,AAL}, ZZI, WAA, IZZ); 
ram_4096x1 sinst_001(SEA,BEA,{ABA,ABB,ABC,ABD,ABE,ABF,ABG,ABH,ABI,ABJ,ABK,ABL}, ZZI, WBA, IZZ); 
ram_4096x1 sinst_002(SIA,BAA,{ACA,ACB,ACC,ACD,ACE,ACF,ACG,ACH,ACI,ACJ,ACK,ACL}, ZZI, WCA, IZZ); 
ram_4096x1 sinst_003(SAB,BAB,{aaa,aab,aac,aad,aae,aaf,aag,aah,aai,aaj,aak,aal}, ZZI, WAB, IZZ); 
ram_4096x1 sinst_004(SEB,BEB,{aba,abb,abc,abd,abe,abf,abg,abh,abi,abj,abk,abl}, ZZI, WBB, IZZ); 
ram_4096x1 sinst_005(SIB,BAB,{aca,acb,acc,acd,ace,acf,acg,ach,aci,acj,ack,acl}, ZZI, WCB, IZZ); 
ram_4096x1 sinst_006(SAC,BAC,{AEA,AEB,AEC,AED,AEE,AEF,AEG,AEH,AEI,AEJ,AEK,AEL}, ZZI, WAC, IZZ); 
ram_4096x1 sinst_007(SEC,BEC,{AFA,AFB,AFC,AFD,AFE,AFF,AFG,AFH,AFI,AFJ,AFK,AFL}, ZZI, WBC, IZZ); 
ram_4096x1 sinst_008(SIC,BAC,{AGA,AGB,AGC,AGD,AGE,AGF,AGG,AGH,AGI,AGJ,AGK,AGL}, ZZI, WCC, IZZ); 
ram_4096x1 sinst_009(SAD,BAD,{aea,aeb,aec,aed,aee,aef,aeg,aeh,aei,aej,aek,ael}, ZZI, WAD, IZZ); 
ram_4096x1 sinst_010(SED,BED,{afa,afb,afc,afd,afe,aff,afg,afh,afi,afj,afk,afl}, ZZI, WBD, IZZ); 
ram_4096x1 sinst_011(SID,BAD,{aga,agb,agc,agd,age,agf,agg,agh,agi,agj,agk,agl}, ZZI, WCD, IZZ); 
ram_4096x1 sinst_012(SAE,BAE,{AAA,AAB,AAC,AAD,AAE,AAF,AAG,AAH,AAI,AAJ,AAK,AAL}, ZZI, WAE, IZZ); 
ram_4096x1 sinst_013(SEE,BEE,{ABA,ABB,ABC,ABD,ABE,ABF,ABG,ABH,ABI,ABJ,ABK,ABL}, ZZI, WBE, IZZ); 
ram_4096x1 sinst_014(SIE,BAE,{ACA,ACB,ACC,ACD,ACE,ACF,ACG,ACH,ACI,ACJ,ACK,ACL}, ZZI, WCE, IZZ); 
ram_4096x1 sinst_015(SAF,BAF,{aaa,aab,aac,aad,aae,aaf,aag,aah,aai,aaj,aak,aal}, ZZI, WAF, IZZ); 
ram_4096x1 sinst_016(SEF,BEF,{aba,abb,abc,abd,abe,abf,abg,abh,abi,abj,abk,abl}, ZZI, WBF, IZZ); 
ram_4096x1 sinst_017(SIH,BAH,{aga,agb,agc,agd,age,agf,agg,agh,agi,agj,agk,agl}, ZZI, WCH, IZZ); 
ram_4096x1 sinst_018(SIF,BAF,{aca,acb,acc,acd,ace,acf,acg,ach,aci,acj,ack,acl}, ZZI, WCF, IZZ); 
ram_4096x1 sinst_019(SAG,BAG,{AEA,AEB,AEC,AED,AEE,AEF,AEG,AEH,AEI,AEJ,AEK,AEL}, ZZI, WAG, IZZ); 
ram_4096x1 sinst_020(SEG,BEG,{AFA,AFB,AFC,AFD,AFE,AFF,AFG,AFH,AFI,AFJ,AFK,AFL}, ZZI, WBG, IZZ); 
ram_4096x1 sinst_021(SIG,BAG,{AGA,AGB,AGC,AGD,AGE,AGF,AGG,AGH,AGI,AGJ,AGK,AGL}, ZZI, WCG, IZZ); 
ram_4096x1 sinst_022(SAH,BAH,{aea,aeb,aec,aed,aee,aef,aeg,aeh,aei,aej,aek,ael}, ZZI, WAH, IZZ); 
ram_4096x1 sinst_023(SEH,BEH,{afa,afb,afc,afd,afe,aff,afg,afh,afi,afj,afk,afl}, ZZI, WBH, IZZ); 
ram_4096x1 sinst_024(SMA,BEA,{ADA,ADB,ADC,ADD,ADE,ADF,ADG,ADH,ADI,ADJ,ADK,ADL}, ZZI, WDA, IZZ); 
ram_4096x1 sinst_025(SMB,BEB,{ada,adb,adc,add,ade,adf,adg,adh,adi,adj,adk,adl}, ZZI, WDB, IZZ); 
ram_4096x1 sinst_026(SMC,BEC,{AHA,AHB,AHC,AHD,AHE,AHF,AHG,AHH,AHI,AHJ,AHK,AHL}, ZZI, WDC, IZZ); 
ram_4096x1 sinst_027(SMD,BED,{aha,ahb,ahc,ahd,ahe,ahf,ahg,ahh,ahi,ahj,ahk,ahl}, ZZI, WDD, IZZ); 
ram_4096x1 sinst_028(SME,BEE,{ADA,ADB,ADC,ADD,ADE,ADF,ADG,ADH,ADI,ADJ,ADK,ADL}, ZZI, WDE, IZZ); 
ram_4096x1 sinst_029(SMF,BEF,{ada,adb,adc,add,ade,adf,adg,adh,adi,adj,adk,adl}, ZZI, WDF, IZZ); 
ram_4096x1 sinst_030(SMG,BEG,{AHA,AHB,AHC,AHD,AHE,AHF,AHG,AHH,AHI,AHJ,AHK,AHL}, ZZI, WDG, IZZ); 
ram_4096x1 sinst_031(SMH,BEH,{aha,ahb,ahc,ahd,ahe,ahf,ahg,ahh,ahi,ahj,ahk,ahl}, ZZI, WDH, IZZ); 
ram_4096x1 sinst_032(SAI,BAI,{AAA,AAB,AAC,AAD,AAE,AAF,AAG,AAH,AAI,AAJ,AAK,AAL}, ZZI, WAI, IZZ); 
ram_4096x1 sinst_033(SEI,BEI,{ABA,ABB,ABC,ABD,ABE,ABF,ABG,ABH,ABI,ABJ,ABK,ABL}, ZZI, WBI, IZZ); 
ram_4096x1 sinst_034(SII,BAI,{ACA,ACB,ACC,ACD,ACE,ACF,ACG,ACH,ACI,ACJ,ACK,ACL}, ZZI, WCI, IZZ); 
ram_4096x1 sinst_035(SAJ,BAJ,{aaa,aab,aac,aad,aae,aaf,aag,aah,aai,aaj,aak,aal}, ZZI, WAJ, IZZ); 
ram_4096x1 sinst_036(SEJ,BEJ,{aba,abb,abc,abd,abe,abf,abg,abh,abi,abj,abk,abl}, ZZI, WBJ, IZZ); 
ram_4096x1 sinst_037(SIJ,BAJ,{aca,acb,acc,acd,ace,acf,acg,ach,aci,acj,ack,acl}, ZZI, WCJ, IZZ); 
ram_4096x1 sinst_038(SAK,BAK,{AEA,AEB,AEC,AED,AEE,AEF,AEG,AEH,AEI,AEJ,AEK,AEL}, ZZI, WAK, IZZ); 
ram_4096x1 sinst_039(SEK,BEK,{AFA,AFB,AFC,AFD,AFE,AFF,AFG,AFH,AFI,AFJ,AFK,AFL}, ZZI, WBK, IZZ); 
ram_4096x1 sinst_040(SIK,BAK,{AGA,AGB,AGC,AGD,AGE,AGF,AGG,AGH,AGI,AGJ,AGK,AGL}, ZZI, WCK, IZZ); 
ram_4096x1 sinst_041(SAL,BAL,{aea,aeb,aec,aed,aee,aef,aeg,aeh,aei,aej,aek,ael}, ZZI, WAL, IZZ); 
ram_4096x1 sinst_042(SEL,BEL,{afa,afb,afc,afd,afe,aff,afg,afh,afi,afj,afk,afl}, ZZI, WBL, IZZ); 
ram_4096x1 sinst_043(SIL,BAL,{aga,agb,agc,agd,age,agf,agg,agh,agi,agj,agk,agl}, ZZI, WCL, IZZ); 
ram_4096x1 sinst_044(SAM,BAM,{AAA,AAB,AAC,AAD,AAE,AAF,AAG,AAH,AAI,AAJ,AAK,AAL}, ZZI, WAM, IZZ); 
ram_4096x1 sinst_045(SEM,BEM,{ABA,ABB,ABC,ABD,ABE,ABF,ABG,ABH,ABI,ABJ,ABK,ABL}, ZZI, WBM, IZZ); 
ram_4096x1 sinst_046(SIM,BAM,{ACA,ACB,ACC,ACD,ACE,ACF,ACG,ACH,ACI,ACJ,ACK,ACL}, ZZI, WCM, IZZ); 
ram_4096x1 sinst_047(SAN,BAN,{aaa,aab,aac,aad,aae,aaf,aag,aah,aai,aaj,aak,aal}, ZZI, WAN, IZZ); 
ram_4096x1 sinst_048(SEN,BEN,{aba,abb,abc,abd,abe,abf,abg,abh,abi,abj,abk,abl}, ZZI, WBN, IZZ); 
ram_4096x1 sinst_049(SIN,BAN,{aca,acb,acc,acd,ace,acf,acg,ach,aci,acj,ack,acl}, ZZI, WCN, IZZ); 
ram_4096x1 sinst_050(SAO,BAO,{AEA,AEB,AEC,AED,AEE,AEF,AEG,AEH,AEI,AEJ,AEK,AEL}, ZZI, WAO, IZZ); 
ram_4096x1 sinst_051(SEO,BEO,{AFA,AFB,AFC,AFD,AFE,AFF,AFG,AFH,AFI,AFJ,AFK,AFL}, ZZI, WBO, IZZ); 
ram_4096x1 sinst_052(SIO,BAO,{AGA,AGB,AGC,AGD,AGE,AGF,AGG,AGH,AGI,AGJ,AGK,AGL}, ZZI, WCO, IZZ); 
ram_4096x1 sinst_053(SAP,BAP,{aea,aeb,aec,aed,aee,aef,aeg,aeh,aei,aej,aek,ael}, ZZI, WAP, IZZ); 
ram_4096x1 sinst_054(SEP,BEP,{afa,afb,afc,afd,afe,aff,afg,afh,afi,afj,afk,afl}, ZZI, WBP, IZZ); 
ram_4096x1 sinst_055(SIP,BAP,{aga,agb,agc,agd,age,agf,agg,agh,agi,agj,agk,agl}, ZZI, WCP, IZZ); 
ram_4096x1 sinst_056(SMI,BEI,{ADA,ADB,ADC,ADD,ADE,ADF,ADG,ADH,ADI,ADJ,ADK,ADL}, ZZI, WDI, IZZ); 
ram_4096x1 sinst_057(SMJ,BEJ,{ada,adb,adc,add,ade,adf,adg,adh,adi,adj,adk,adl}, ZZI, WDJ, IZZ); 
ram_4096x1 sinst_058(SMK,BEK,{AHA,AHB,AHC,AHD,AHE,AHF,AHG,AHH,AHI,AHJ,AHK,AHL}, ZZI, WDK, IZZ); 
ram_4096x1 sinst_059(SML,BEL,{aha,ahb,ahc,ahd,ahe,ahf,ahg,ahh,ahi,ahj,ahk,ahl}, ZZI, WDL, IZZ); 
ram_4096x1 sinst_060(SMM,BEM,{ADA,ADB,ADC,ADD,ADE,ADF,ADG,ADH,ADI,ADJ,ADK,ADL}, ZZI, WDM, IZZ); 
ram_4096x1 sinst_061(SMN,BEN,{ada,adb,adc,add,ade,adf,adg,adh,adi,adj,adk,adl}, ZZI, WDN, IZZ); 
ram_4096x1 sinst_062(SMO,BEO,{AHA,AHB,AHC,AHD,AHE,AHF,AHG,AHH,AHI,AHJ,AHK,AHL}, ZZI, WDO, IZZ); 
ram_4096x1 sinst_063(SMP,BEP,{aha,ahb,ahc,ahd,ahe,ahf,ahg,ahh,ahi,ahj,ahk,ahl}, ZZI, WDP, IZZ); 
ram_4096x1 sinst_064(SBA,BBA,{AAA,AAB,AAC,AAD,AAE,AAF,AAG,AAH,AAI,AAJ,AAK,AAL}, ZZI, WAA, IZZ); 
ram_4096x1 sinst_065(SFA,BFA,{ABA,ABB,ABC,ABD,ABE,ABF,ABG,ABH,ABI,ABJ,ABK,ABL}, ZZI, WBA, IZZ); 
ram_4096x1 sinst_066(SJA,BBA,{ACA,ACB,ACC,ACD,ACE,ACF,ACG,ACH,ACI,ACJ,ACK,ACL}, ZZI, WCA, IZZ); 
ram_4096x1 sinst_067(SBB,BBB,{aaa,aab,aac,aad,aae,aaf,aag,aah,aai,aaj,aak,aal}, ZZI, WAB, IZZ); 
ram_4096x1 sinst_068(SFB,BFB,{aba,abb,abc,abd,abe,abf,abg,abh,abi,abj,abk,abl}, ZZI, WBB, IZZ); 
ram_4096x1 sinst_069(SJB,BBB,{aca,acb,acc,acd,ace,acf,acg,ach,aci,acj,ack,acl}, ZZI, WCB, IZZ); 
ram_4096x1 sinst_070(SBC,BBC,{AEA,AEB,AEC,AED,AEE,AEF,AEG,AEH,AEI,AEJ,AEK,AEL}, ZZI, WAC, IZZ); 
ram_4096x1 sinst_071(SFC,BFC,{AFA,AFB,AFC,AFD,AFE,AFF,AFG,AFH,AFI,AFJ,AFK,AFL}, ZZI, WBC, IZZ); 
ram_4096x1 sinst_072(SJC,BBC,{AGA,AGB,AGC,AGD,AGE,AGF,AGG,AGH,AGI,AGJ,AGK,AGL}, ZZI, WCC, IZZ); 
ram_4096x1 sinst_073(SBD,BBD,{aea,aeb,aec,aed,aee,aef,aeg,aeh,aei,aej,aek,ael}, ZZI, WAD, IZZ); 
ram_4096x1 sinst_074(SFD,BFD,{afa,afb,afc,afd,afe,aff,afg,afh,afi,afj,afk,afl}, ZZI, WBD, IZZ); 
ram_4096x1 sinst_075(SJD,BBD,{aga,agb,agc,agd,age,agf,agg,agh,agi,agj,agk,agl}, ZZI, WCD, IZZ); 
ram_4096x1 sinst_076(SBE,BBE,{AAA,AAB,AAC,AAD,AAE,AAF,AAG,AAH,AAI,AAJ,AAK,AAL}, ZZI, WAE, IZZ); 
ram_4096x1 sinst_077(SFE,BFE,{ABA,ABB,ABC,ABD,ABE,ABF,ABG,ABH,ABI,ABJ,ABK,ABL}, ZZI, WBE, IZZ); 
ram_4096x1 sinst_078(SJE,BBE,{ACA,ACB,ACC,ACD,ACE,ACF,ACG,ACH,ACI,ACJ,ACK,ACL}, ZZI, WCE, IZZ); 
ram_4096x1 sinst_079(SBF,BBF,{aaa,aab,aac,aad,aae,aaf,aag,aah,aai,aaj,aak,aal}, ZZI, WAF, IZZ); 
ram_4096x1 sinst_080(SFF,BFF,{aba,abb,abc,abd,abe,abf,abg,abh,abi,abj,abk,abl}, ZZI, WBF, IZZ); 
ram_4096x1 sinst_081(SJF,BBF,{aca,acb,acc,acd,ace,acf,acg,ach,aci,acj,ack,acl}, ZZI, WCF, IZZ); 
ram_4096x1 sinst_082(SBG,BBG,{AEA,AEB,AEC,AED,AEE,AEF,AEG,AEH,AEI,AEJ,AEK,AEL}, ZZI, WAG, IZZ); 
ram_4096x1 sinst_083(SFG,BFG,{AFA,AFB,AFC,AFD,AFE,AFF,AFG,AFH,AFI,AFJ,AFK,AFL}, ZZI, WBG, IZZ); 
ram_4096x1 sinst_084(SJG,BBG,{AGA,AGB,AGC,AGD,AGE,AGF,AGG,AGH,AGI,AGJ,AGK,AGL}, ZZI, WCG, IZZ); 
ram_4096x1 sinst_085(SBH,BBH,{aea,aeb,aec,aed,aee,aef,aeg,aeh,aei,aej,aek,ael}, ZZI, WAH, IZZ); 
ram_4096x1 sinst_086(SFH,BFH,{afa,afb,afc,afd,afe,aff,afg,afh,afi,afj,afk,afl}, ZZI, WBH, IZZ); 
ram_4096x1 sinst_087(SJH,BBH,{aga,agb,agc,agd,age,agf,agg,agh,agi,agj,agk,agl}, ZZI, WCH, IZZ); 
ram_4096x1 sinst_088(SNA,BFA,{ADA,ADB,ADC,ADD,ADE,ADF,ADG,ADH,ADI,ADJ,ADK,ADL}, ZZI, WDA, IZZ); 
ram_4096x1 sinst_089(SNB,BFB,{ada,adb,adc,add,ade,adf,adg,adh,adi,adj,adk,adl}, ZZI, WDB, IZZ); 
ram_4096x1 sinst_090(SNC,BFC,{AHA,AHB,AHC,AHD,AHE,AHF,AHG,AHH,AHI,AHJ,AHK,AHL}, ZZI, WDC, IZZ); 
ram_4096x1 sinst_091(SND,BFD,{aha,ahb,ahc,ahd,ahe,ahf,ahg,ahh,ahi,ahj,ahk,ahl}, ZZI, WDD, IZZ); 
ram_4096x1 sinst_092(SNE,BFE,{ADA,ADB,ADC,ADD,ADE,ADF,ADG,ADH,ADI,ADJ,ADK,ADL}, ZZI, WDE, IZZ); 
ram_4096x1 sinst_093(SNF,BFF,{ada,adb,adc,add,ade,adf,adg,adh,adi,adj,adk,adl}, ZZI, WDF, IZZ); 
ram_4096x1 sinst_094(SNG,BFG,{AHA,AHB,AHC,AHD,AHE,AHF,AHG,AHH,AHI,AHJ,AHK,AHL}, ZZI, WDG, IZZ); 
ram_4096x1 sinst_095(SNH,BFH,{aha,ahb,ahc,ahd,ahe,ahf,ahg,ahh,ahi,ahj,ahk,ahl}, ZZI, WDH, IZZ); 
ram_4096x1 sinst_096(SBI,BBI,{AAA,AAB,AAC,AAD,AAE,AAF,AAG,AAH,AAI,AAJ,AAK,AAL}, ZZI, WAI, IZZ); 
ram_4096x1 sinst_097(SNI,BFI,{ADA,ADB,ADC,ADD,ADE,ADF,ADG,ADH,ADI,ADJ,ADK,ADL}, ZZI, WDI, IZZ); 
ram_4096x1 sinst_098(SFI,BFI,{ABA,ABB,ABC,ABD,ABE,ABF,ABG,ABH,ABI,ABJ,ABK,ABL}, ZZI, WBI, IZZ); 
ram_4096x1 sinst_099(SJI,BBI,{ACA,ACB,ACC,ACD,ACE,ACF,ACG,ACH,ACI,ACJ,ACK,ACL}, ZZI, WCI, IZZ); 
ram_4096x1 sinst_100(SBJ,BBJ,{aaa,aab,aac,aad,aae,aaf,aag,aah,aai,aaj,aak,aal}, ZZI, WAJ, IZZ); 
ram_4096x1 sinst_101(SNJ,BFJ,{ada,adb,adc,add,ade,adf,adg,adh,adi,adj,adk,adl}, ZZI, WDJ, IZZ); 
ram_4096x1 sinst_102(SFJ,BFJ,{aba,abb,abc,abd,abe,abf,abg,abh,abi,abj,abk,abl}, ZZI, WBJ, IZZ); 
ram_4096x1 sinst_103(SJJ,BBJ,{aca,acb,acc,acd,ace,acf,acg,ach,aci,acj,ack,acl}, ZZI, WCJ, IZZ); 
ram_4096x1 sinst_104(SBK,BBK,{AEA,AEB,AEC,AED,AEE,AEF,AEG,AEH,AEI,AEJ,AEK,AEL}, ZZI, WAK, IZZ); 
ram_4096x1 sinst_105(SNK,BFK,{AHA,AHB,AHC,AHD,AHE,AHF,AHG,AHH,AHI,AHJ,AHK,AHL}, ZZI, WDK, IZZ); 
ram_4096x1 sinst_106(SFK,BFK,{AFA,AFB,AFC,AFD,AFE,AFF,AFG,AFH,AFI,AFJ,AFK,AFL}, ZZI, WBK, IZZ); 
ram_4096x1 sinst_107(SJK,BBK,{AGA,AGB,AGC,AGD,AGE,AGF,AGG,AGH,AGI,AGJ,AGK,AGL}, ZZI, WCK, IZZ); 
ram_4096x1 sinst_108(SBL,BBL,{aea,aeb,aec,aed,aee,aef,aeg,aeh,aei,aej,aek,ael}, ZZI, WAL, IZZ); 
ram_4096x1 sinst_109(SNL,BFL,{aha,ahb,ahc,ahd,ahe,ahf,ahg,ahh,ahi,ahj,ahk,ahl}, ZZI, WDL, IZZ); 
ram_4096x1 sinst_110(SFL,BFL,{afa,afb,afc,afd,afe,aff,afg,afh,afi,afj,afk,afl}, ZZI, WBL, IZZ); 
ram_4096x1 sinst_111(SJL,BBL,{aga,agb,agc,agd,age,agf,agg,agh,agi,agj,agk,agl}, ZZI, WCL, IZZ); 
ram_4096x1 sinst_112(SBM,BBM,{AAA,AAB,AAC,AAD,AAE,AAF,AAG,AAH,AAI,AAJ,AAK,AAL}, ZZI, WAM, IZZ); 
ram_4096x1 sinst_113(SNM,BFM,{ADA,ADB,ADC,ADD,ADE,ADF,ADG,ADH,ADI,ADJ,ADK,ADL}, ZZI, WDM, IZZ); 
ram_4096x1 sinst_114(SFM,BFM,{ABA,ABB,ABC,ABD,ABE,ABF,ABG,ABH,ABI,ABJ,ABK,ABL}, ZZI, WBM, IZZ); 
ram_4096x1 sinst_115(SJM,BBM,{ACA,ACB,ACC,ACD,ACE,ACF,ACG,ACH,ACI,ACJ,ACK,ACL}, ZZI, WCM, IZZ); 
ram_4096x1 sinst_116(SBN,BBN,{aaa,aab,aac,aad,aae,aaf,aag,aah,aai,aaj,aak,aal}, ZZI, WAN, IZZ); 
ram_4096x1 sinst_117(SNN,BFN,{ada,adb,adc,add,ade,adf,adg,adh,adi,adj,adk,adl}, ZZI, WDN, IZZ); 
ram_4096x1 sinst_118(SFN,BFN,{aba,abb,abc,abd,abe,abf,abg,abh,abi,abj,abk,abl}, ZZI, WBN, IZZ); 
ram_4096x1 sinst_119(SJN,BBN,{aca,acb,acc,acd,ace,acf,acg,ach,aci,acj,ack,acl}, ZZI, WCN, IZZ); 
ram_4096x1 sinst_120(SBO,BBO,{AEA,AEB,AEC,AED,AEE,AEF,AEG,AEH,AEI,AEJ,AEK,AEL}, ZZI, WAO, IZZ); 
ram_4096x1 sinst_121(SNO,BFO,{AHA,AHB,AHC,AHD,AHE,AHF,AHG,AHH,AHI,AHJ,AHK,AHL}, ZZI, WDO, IZZ); 
ram_4096x1 sinst_122(SFO,BFO,{AFA,AFB,AFC,AFD,AFE,AFF,AFG,AFH,AFI,AFJ,AFK,AFL}, ZZI, WBO, IZZ); 
ram_4096x1 sinst_123(SJO,BBO,{AGA,AGB,AGC,AGD,AGE,AGF,AGG,AGH,AGI,AGJ,AGK,AGL}, ZZI, WCO, IZZ); 
ram_4096x1 sinst_124(SBP,BBP,{aea,aeb,aec,aed,aee,aef,aeg,aeh,aei,aej,aek,ael}, ZZI, WAP, IZZ); 
ram_4096x1 sinst_125(SFP,BFP,{afa,afb,afc,afd,afe,aff,afg,afh,afi,afj,afk,afl}, ZZI, WBP, IZZ); 
ram_4096x1 sinst_126(SNP,BFP,{aha,ahb,ahc,ahd,ahe,ahf,ahg,ahh,ahi,ahj,ahk,ahl}, ZZI, WDP, IZZ); 
ram_4096x1 sinst_127(SJP,BBP,{aga,agb,agc,agd,age,agf,agg,agh,agi,agj,agk,agl}, ZZI, WCP, IZZ); 
ram_4096x1 sinst_128(SCA,BCA,{AAA,AAB,AAC,AAD,AAE,AAF,AAG,AAH,AAI,AAJ,AAK,AAL}, ZZI, WAA, IZZ); 
ram_4096x1 sinst_129(SGA,BGA,{ABA,ABB,ABC,ABD,ABE,ABF,ABG,ABH,ABI,ABJ,ABK,ABL}, ZZI, WBA, IZZ); 
ram_4096x1 sinst_130(SKA,BCA,{ACA,ACB,ACC,ACD,ACE,ACF,ACG,ACH,ACI,ACJ,ACK,ACL}, ZZI, WCA, IZZ); 
ram_4096x1 sinst_131(SCB,BCB,{aaa,aab,aac,aad,aae,aaf,aag,aah,aai,aaj,aak,aal}, ZZI, WAB, IZZ); 
ram_4096x1 sinst_132(SGB,BGB,{aba,abb,abc,abd,abe,abf,abg,abh,abi,abj,abk,abl}, ZZI, WBB, IZZ); 
ram_4096x1 sinst_133(SKB,BCB,{aca,acb,acc,acd,ace,acf,acg,ach,aci,acj,ack,acl}, ZZI, WCB, IZZ); 
ram_4096x1 sinst_134(SCC,BCC,{AEA,AEB,AEC,AED,AEE,AEF,AEG,AEH,AEI,AEJ,AEK,AEL}, ZZI, WAC, IZZ); 
ram_4096x1 sinst_135(SGC,BGC,{AFA,AFB,AFC,AFD,AFE,AFF,AFG,AFH,AFI,AFJ,AFK,AFL}, ZZI, WBC, IZZ); 
ram_4096x1 sinst_136(SKC,BCC,{AGA,AGB,AGC,AGD,AGE,AGF,AGG,AGH,AGI,AGJ,AGK,AGL}, ZZI, WCC, IZZ); 
ram_4096x1 sinst_137(SCD,BCD,{aea,aeb,aec,aed,aee,aef,aeg,aeh,aei,aej,aek,ael}, ZZI, WAD, IZZ); 
ram_4096x1 sinst_138(SGD,BGD,{afa,afb,afc,afd,afe,aff,afg,afh,afi,afj,afk,afl}, ZZI, WBD, IZZ); 
ram_4096x1 sinst_139(SKD,BCD,{aga,agb,agc,agd,age,agf,agg,agh,agi,agj,agk,agl}, ZZI, WCD, IZZ); 
ram_4096x1 sinst_140(SCE,BCE,{AAA,AAB,AAC,AAD,AAE,AAF,AAG,AAH,AAI,AAJ,AAK,AAL}, ZZI, WAE, IZZ); 
ram_4096x1 sinst_141(SGE,BGE,{ABA,ABB,ABC,ABD,ABE,ABF,ABG,ABH,ABI,ABJ,ABK,ABL}, ZZI, WBE, IZZ); 
ram_4096x1 sinst_142(SKE,BCE,{ACA,ACB,ACC,ACD,ACE,ACF,ACG,ACH,ACI,ACJ,ACK,ACL}, ZZI, WCE, IZZ); 
ram_4096x1 sinst_143(SCF,BCF,{aaa,aab,aac,aad,aae,aaf,aag,aah,aai,aaj,aak,aal}, ZZI, WAF, IZZ); 
ram_4096x1 sinst_144(SGF,BGF,{aba,abb,abc,abd,abe,abf,abg,abh,abi,abj,abk,abl}, ZZI, WBF, IZZ); 
ram_4096x1 sinst_145(SKF,BCF,{aca,acb,acc,acd,ace,acf,acg,ach,aci,acj,ack,acl}, ZZI, WCF, IZZ); 
ram_4096x1 sinst_146(SCG,BCG,{AEA,AEB,AEC,AED,AEE,AEF,AEG,AEH,AEI,AEJ,AEK,AEL}, ZZI, WAG, IZZ); 
ram_4096x1 sinst_147(SGG,BGG,{AFA,AFB,AFC,AFD,AFE,AFF,AFG,AFH,AFI,AFJ,AFK,AFL}, ZZI, WBG, IZZ); 
ram_4096x1 sinst_148(SKG,BCG,{AGA,AGB,AGC,AGD,AGE,AGF,AGG,AGH,AGI,AGJ,AGK,AGL}, ZZI, WCG, IZZ); 
ram_4096x1 sinst_149(SCH,BCH,{aea,aeb,aec,aed,aee,aef,aeg,aeh,aei,aej,aek,ael}, ZZI, WAH, IZZ); 
ram_4096x1 sinst_150(SGH,BGH,{afa,afb,afc,afd,afe,aff,afg,afh,afi,afj,afk,afl}, ZZI, WBH, IZZ); 
ram_4096x1 sinst_151(SKH,BCH,{aga,agb,agc,agd,age,agf,agg,agh,agi,agj,agk,agl}, ZZI, WCH, IZZ); 
ram_4096x1 sinst_152(SOA,BGA,{ADA,ADB,ADC,ADD,ADE,ADF,ADG,ADH,ADI,ADJ,ADK,ADL}, ZZI, WDA, IZZ); 
ram_4096x1 sinst_153(SOB,BGB,{ada,adb,adc,add,ade,adf,adg,adh,adi,adj,adk,adl}, ZZI, WDB, IZZ); 
ram_4096x1 sinst_154(SOC,BGC,{AHA,AHB,AHC,AHD,AHE,AHF,AHG,AHH,AHI,AHJ,AHK,AHL}, ZZI, WDC, IZZ); 
ram_4096x1 sinst_155(SOD,BGD,{aha,ahb,ahc,ahd,ahe,ahf,ahg,ahh,ahi,ahj,ahk,ahl}, ZZI, WDD, IZZ); 
ram_4096x1 sinst_156(SOE,BGE,{ADA,ADB,ADC,ADD,ADE,ADF,ADG,ADH,ADI,ADJ,ADK,ADL}, ZZI, WDE, IZZ); 
ram_4096x1 sinst_157(SOF,BGF,{ada,adb,adc,add,ade,adf,adg,adh,adi,adj,adk,adl}, ZZI, WDF, IZZ); 
ram_4096x1 sinst_158(SOG,BGG,{AHA,AHB,AHC,AHD,AHE,AHF,AHG,AHH,AHI,AHJ,AHK,AHL}, ZZI, WDG, IZZ); 
ram_4096x1 sinst_159(SOH,BGH,{aha,ahb,ahc,ahd,ahe,ahf,ahg,ahh,ahi,ahj,ahk,ahl}, ZZI, WDH, IZZ); 
ram_4096x1 sinst_160(SCI,BCI,{AAA,AAB,AAC,AAD,AAE,AAF,AAG,AAH,AAI,AAJ,AAK,AAL}, ZZI, WAI, IZZ); 
ram_4096x1 sinst_161(SGI,BGI,{ABA,ABB,ABC,ABD,ABE,ABF,ABG,ABH,ABI,ABJ,ABK,ABL}, ZZI, WBI, IZZ); 
ram_4096x1 sinst_162(SKI,BCI,{ACA,ACB,ACC,ACD,ACE,ACF,ACG,ACH,ACI,ACJ,ACK,ACL}, ZZI, WCI, IZZ); 
ram_4096x1 sinst_163(SCJ,BCJ,{aaa,aab,aac,aad,aae,aaf,aag,aah,aai,aaj,aak,aal}, ZZI, WAJ, IZZ); 
ram_4096x1 sinst_164(SGJ,BGJ,{aba,abb,abc,abd,abe,abf,abg,abh,abi,abj,abk,abl}, ZZI, WBJ, IZZ); 
ram_4096x1 sinst_165(SKJ,BCJ,{aca,acb,acc,acd,ace,acf,acg,ach,aci,acj,ack,acl}, ZZI, WCJ, IZZ); 
ram_4096x1 sinst_166(SCK,BCK,{AEA,AEB,AEC,AED,AEE,AEF,AEG,AEH,AEI,AEJ,AEK,AEL}, ZZI, WAK, IZZ); 
ram_4096x1 sinst_167(SGK,BGK,{AFA,AFB,AFC,AFD,AFE,AFF,AFG,AFH,AFI,AFJ,AFK,AFL}, ZZI, WBK, IZZ); 
ram_4096x1 sinst_168(SKK,BCK,{AGA,AGB,AGC,AGD,AGE,AGF,AGG,AGH,AGI,AGJ,AGK,AGL}, ZZI, WCK, IZZ); 
ram_4096x1 sinst_169(SCL,BCL,{aea,aeb,aec,aed,aee,aef,aeg,aeh,aei,aej,aek,ael}, ZZI, WAL, IZZ); 
ram_4096x1 sinst_170(SGL,BGL,{afa,afb,afc,afd,afe,aff,afg,afh,afi,afj,afk,afl}, ZZI, WBL, IZZ); 
ram_4096x1 sinst_171(SKL,BCL,{aga,agb,agc,agd,age,agf,agg,agh,agi,agj,agk,agl}, ZZI, WCL, IZZ); 
ram_4096x1 sinst_172(SCM,BCM,{AAA,AAB,AAC,AAD,AAE,AAF,AAG,AAH,AAI,AAJ,AAK,AAL}, ZZI, WAM, IZZ); 
ram_4096x1 sinst_173(SGM,BGM,{ABA,ABB,ABC,ABD,ABE,ABF,ABG,ABH,ABI,ABJ,ABK,ABL}, ZZI, WBM, IZZ); 
ram_4096x1 sinst_174(SKM,BCM,{ACA,ACB,ACC,ACD,ACE,ACF,ACG,ACH,ACI,ACJ,ACK,ACL}, ZZI, WCM, IZZ); 
ram_4096x1 sinst_175(SCN,BCN,{aaa,aab,aac,aad,aae,aaf,aag,aah,aai,aaj,aak,aal}, ZZI, WAN, IZZ); 
ram_4096x1 sinst_176(SGN,BGN,{aba,abb,abc,abd,abe,abf,abg,abh,abi,abj,abk,abl}, ZZI, WBN, IZZ); 
ram_4096x1 sinst_177(SKN,BCN,{aca,acb,acc,acd,ace,acf,acg,ach,aci,acj,ack,acl}, ZZI, WCN, IZZ); 
ram_4096x1 sinst_178(SCO,BCO,{AEA,AEB,AEC,AED,AEE,AEF,AEG,AEH,AEI,AEJ,AEK,AEL}, ZZI, WAO, IZZ); 
ram_4096x1 sinst_179(SGO,BGO,{AFA,AFB,AFC,AFD,AFE,AFF,AFG,AFH,AFI,AFJ,AFK,AFL}, ZZI, WBO, IZZ); 
ram_4096x1 sinst_180(SKO,BCO,{AGA,AGB,AGC,AGD,AGE,AGF,AGG,AGH,AGI,AGJ,AGK,AGL}, ZZI, WCO, IZZ); 
ram_4096x1 sinst_181(SCP,BCP,{aea,aeb,aec,aed,aee,aef,aeg,aeh,aei,aej,aek,ael}, ZZI, WAP, IZZ); 
ram_4096x1 sinst_182(SGP,BGP,{afa,afb,afc,afd,afe,aff,afg,afh,afi,afj,afk,afl}, ZZI, WBP, IZZ); 
ram_4096x1 sinst_183(SKP,BCP,{aga,agb,agc,agd,age,agf,agg,agh,agi,agj,agk,agl}, ZZI, WCP, IZZ); 
ram_4096x1 sinst_184(SOI,BGI,{ADA,ADB,ADC,ADD,ADE,ADF,ADG,ADH,ADI,ADJ,ADK,ADL}, ZZI, WDI, IZZ); 
ram_4096x1 sinst_185(SOJ,BGJ,{ada,adb,adc,add,ade,adf,adg,adh,adi,adj,adk,adl}, ZZI, WDJ, IZZ); 
ram_4096x1 sinst_186(SOK,BGK,{AHA,AHB,AHC,AHD,AHE,AHF,AHG,AHH,AHI,AHJ,AHK,AHL}, ZZI, WDK, IZZ); 
ram_4096x1 sinst_187(SOL,BGL,{ada,adb,adc,add,ade,adf,adg,adh,adi,adj,adk,adl}, ZZI, WDL, IZZ); 
ram_4096x1 sinst_188(SOM,BGM,{ADA,ADB,ADC,ADD,ADE,ADF,ADG,ADH,ADI,ADJ,ADK,ADL}, ZZI, WDM, IZZ); 
ram_4096x1 sinst_189(SON,BGN,{ada,adb,adc,add,ade,adf,adg,adh,adi,adj,adk,adl}, ZZI, WDN, IZZ); 
ram_4096x1 sinst_190(SOO,BGO,{AHA,AHB,AHC,AHD,AHE,AHF,AHG,AHH,AHI,AHJ,AHK,AHL}, ZZI, WDO, IZZ); 
ram_4096x1 sinst_191(SOP,BGP,{aha,ahb,ahc,ahd,ahe,ahf,ahg,ahh,ahi,ahj,ahk,ahl}, ZZI, WDP, IZZ); 
ram_4096x1 sinst_192(SDA,BDA,{AAA,AAB,AAC,AAD,AAE,AAF,AAG,AAH,AAI,AAJ,AAK,AAL}, ZZI, WAA, IZZ); 
ram_4096x1 sinst_193(SHA,BHA,{ABA,ABB,ABC,ABD,ABE,ABF,ABG,ABH,ABI,ABJ,ABK,ABL}, ZZI, WBA, IZZ); 
ram_4096x1 sinst_194(SLA,BDA,{ACA,ACB,ACC,ACD,ACE,ACF,ACG,ACH,ACI,ACJ,ACK,ACL}, ZZI, WCA, IZZ); 
ram_4096x1 sinst_195(SDB,BDB,{aaa,aab,aac,aad,aae,aaf,aag,aah,aai,aaj,aak,aal}, ZZI, WAB, IZZ); 
ram_4096x1 sinst_196(SHB,BHB,{aba,abb,abc,abd,abe,abf,abg,abh,abi,abj,abk,abl}, ZZI, WBB, IZZ); 
ram_4096x1 sinst_197(SLB,BDB,{aca,acb,acc,acd,ace,acf,acg,ach,aci,acj,ack,acl}, ZZI, WCB, IZZ); 
ram_4096x1 sinst_198(SDC,BDC,{AAA,AAB,AAC,AAD,AAE,AAF,AAG,AAH,AAI,AAJ,AAK,AAL}, ZZI, WAC, IZZ); 
ram_4096x1 sinst_199(SHC,BHC,{AFA,AFB,AFC,AFD,AFE,AFF,AFG,AFH,AFI,AFJ,AFK,AFL}, ZZI, WBC, IZZ); 
ram_4096x1 sinst_200(SLC,BDC,{AGA,AGB,AGC,AGD,AGE,AGF,AGG,AGH,AGI,AGJ,AGK,AGL}, ZZI, WCC, IZZ); 
ram_4096x1 sinst_201(SDD,BDD,{aea,aeb,aec,aed,aee,aef,aeg,aeh,aei,aej,aek,ael}, ZZI, WAD, IZZ); 
ram_4096x1 sinst_202(SHD,BHD,{afa,afb,afc,afd,afe,aff,afg,afh,afi,afj,afk,afl}, ZZI, WBD, IZZ); 
ram_4096x1 sinst_203(SLD,BDD,{aga,agb,agc,agd,age,agf,agg,agh,agi,agj,agk,agl}, ZZI, WCD, IZZ); 
ram_4096x1 sinst_204(SDE,BDE,{AAA,AAB,AAC,AAD,AAE,AAF,AAG,AAH,AAI,AAJ,AAK,AAL}, ZZI, WAE, IZZ); 
ram_4096x1 sinst_205(SHE,BHE,{ABA,ABB,ABC,ABD,ABE,ABF,ABG,ABH,ABI,ABJ,ABK,ABL}, ZZI, WBE, IZZ); 
ram_4096x1 sinst_206(SLE,BDE,{ACA,ACB,ACC,ACD,ACE,ACF,ACG,ACH,ACI,ACJ,ACK,ACL}, ZZI, WCE, IZZ); 
ram_4096x1 sinst_207(SDF,BDF,{aaa,aab,aac,aad,aae,aaf,aag,aah,aai,aaj,aak,aal}, ZZI, WAF, IZZ); 
ram_4096x1 sinst_208(SHF,BHF,{aba,abb,abc,abd,abe,abf,abg,abh,abi,abj,abk,abl}, ZZI, WBF, IZZ); 
ram_4096x1 sinst_209(SLF,BDF,{aca,acb,acc,acd,ace,acf,acg,ach,aci,acj,ack,acl}, ZZI, WCF, IZZ); 
ram_4096x1 sinst_210(SDG,BDG,{AEA,AEB,AEC,AED,AEE,AEF,AEG,AEH,AEI,AEJ,AEK,AEL}, ZZI, WAG, IZZ); 
ram_4096x1 sinst_211(SHG,BHG,{AFA,AFB,AFC,AFD,AFE,AFF,AFG,AFH,AFI,AFJ,AFK,AFL}, ZZI, WBG, IZZ); 
ram_4096x1 sinst_212(SLG,BDG,{AGA,AGB,AGC,AGD,AGE,AGF,AGG,AGH,AGI,AGJ,AGK,AGL}, ZZI, WCG, IZZ); 
ram_4096x1 sinst_213(SDH,BDH,{aea,aeb,aec,aed,aee,aef,aeg,aeh,aei,aej,aek,ael}, ZZI, WAH, IZZ); 
ram_4096x1 sinst_214(SHH,BHH,{afa,afb,afc,afd,afe,aff,afg,afh,afi,afj,afk,afl}, ZZI, WBH, IZZ); 
ram_4096x1 sinst_215(SLH,BDH,{aga,agb,agc,agd,age,agf,agg,agh,agi,agj,agk,agl}, ZZI, WCH, IZZ); 
ram_4096x1 sinst_216(SPI,BHI,{ADA,ADB,ADC,ADD,ADE,ADF,ADG,ADH,ADI,ADJ,ADK,ADL}, ZZI, WDI, IZZ); 
ram_4096x1 sinst_217(SPB,BHB,{ada,adb,adc,add,ade,adf,adg,adh,adi,adj,adk,adl}, ZZI, WDB, IZZ); 
ram_4096x1 sinst_218(SPJ,BHJ,{ada,adb,adc,add,ade,adf,adg,adh,adi,adj,adk,adl}, ZZI, WDJ, IZZ); 
ram_4096x1 sinst_219(SPC,BHC,{AHA,AHB,AHC,AHD,AHE,AHF,AHG,AHH,AHI,AHJ,AHK,AHL}, ZZI, WDC, IZZ); 
ram_4096x1 sinst_220(SPK,BHK,{AHA,AHB,AHC,AHD,AHE,AHF,AHG,AHH,AHI,AHJ,AHK,AHL}, ZZI, WDK, IZZ); 
ram_4096x1 sinst_221(SPL,BHL,{aha,ahb,ahc,ahd,ahe,ahf,ahg,ahh,ahi,ahj,ahk,ahl}, ZZI, WDL, IZZ); 
ram_4096x1 sinst_222(SPD,BHD,{aha,ahb,ahc,ahd,ahe,ahf,ahg,ahh,ahi,ahj,ahk,ahl}, ZZI, WDD, IZZ); 
ram_4096x1 sinst_223(SPE,BHE,{ADA,ADB,ADC,ADD,ADE,ADF,ADG,ADH,ADI,ADJ,ADK,ADL}, ZZI, WDE, IZZ); 
ram_4096x1 sinst_224(SPM,BHM,{ADA,ADB,ADC,ADD,ADE,ADF,ADG,ADH,ADI,ADJ,ADK,ADL}, ZZI, WDM, IZZ); 
ram_4096x1 sinst_225(SPF,BHF,{ada,adb,adc,add,ade,adf,adg,adh,adi,adj,adk,adl}, ZZI, WDF, IZZ); 
ram_4096x1 sinst_226(SPN,BHN,{ada,adb,adc,add,ade,adf,adg,adh,adi,adj,adk,adl}, ZZI, WDN, IZZ); 
ram_4096x1 sinst_227(SPG,BHG,{AHA,AHB,AHC,AHD,AHE,AHF,AHG,AHH,AHI,AHJ,AHK,AHL}, ZZI, WDG, IZZ); 
ram_4096x1 sinst_228(SPO,BHO,{AHA,AHB,AHC,AHD,AHE,AHF,AHG,AHH,AHI,AHJ,AHK,AHL}, ZZI, WDO, IZZ); 
ram_4096x1 sinst_229(SPH,BHH,{aha,ahb,ahc,ahd,ahe,ahf,ahg,ahh,ahi,ahj,ahk,ahl}, ZZI, WDH, IZZ); 
ram_4096x1 sinst_230(SPP,BHP,{aha,ahb,ahc,ahd,ahe,ahf,ahg,ahh,ahi,ahj,ahk,ahl}, ZZI, WDP, IZZ); 
ram_4096x1 sinst_231(SPA,BHA,{ADA,ADB,ADC,ADD,ADE,ADF,ADG,ADH,ADI,ADJ,ADK,ADL}, ZZI, WDA, IZZ); 
ram_4096x1 sinst_232(SDI,BDI,{AAA,AAB,AAC,AAD,AAE,AAF,AAG,AAH,AAI,AAJ,AAK,AAL}, ZZI, WAI, IZZ); 
ram_4096x1 sinst_233(SHI,BHI,{ABA,ABB,ABC,ABD,ABE,ABF,ABG,ABH,ABI,ABJ,ABK,ABL}, ZZI, WBI, IZZ); 
ram_4096x1 sinst_234(SLI,BDI,{ACA,ACB,ACC,ACD,ACE,ACF,ACG,ACH,ACI,ACJ,ACK,ACL}, ZZI, WCI, IZZ); 
ram_4096x1 sinst_235(SDJ,BDJ,{aaa,aab,aac,aad,aae,aaf,aag,aah,aai,aaj,aak,aal}, ZZI, WAJ, IZZ); 
ram_4096x1 sinst_236(SHJ,BHJ,{aba,abb,abc,abd,abe,abf,abg,abh,abi,abj,abk,abl}, ZZI, WBJ, IZZ); 
ram_4096x1 sinst_237(SLJ,BDJ,{aca,acb,acc,acd,ace,acf,acg,ach,aci,acj,ack,acl}, ZZI, WCJ, IZZ); 
ram_4096x1 sinst_238(SDK,BDK,{AEA,AEB,AEC,AED,AEE,AEF,AEG,AEH,AEI,AEJ,AEK,AEL}, ZZI, WAK, IZZ); 
ram_4096x1 sinst_239(SHK,BHK,{AFA,AFB,AFC,AFD,AFE,AFF,AFG,AFH,AFI,AFJ,AFK,AFL}, ZZI, WBK, IZZ); 
ram_4096x1 sinst_240(SLK,BDK,{AGA,AGB,AGC,AGD,AGE,AGF,AGG,AGH,AGI,AGJ,AGK,AGL}, ZZI, WCK, IZZ); 
ram_4096x1 sinst_241(SDL,BDL,{aea,aeb,aec,aed,aee,aef,aeg,aeh,aei,aej,aek,ael}, ZZI, WAL, IZZ); 
ram_4096x1 sinst_242(SHL,BHL,{afa,afb,afc,afd,afe,aff,afg,afh,afi,afj,afk,afl}, ZZI, WBL, IZZ); 
ram_4096x1 sinst_243(SLL,BDL,{aga,agb,agc,agd,age,agf,agg,agh,agi,agj,agk,agl}, ZZI, WCL, IZZ); 
ram_4096x1 sinst_244(SDM,BDM,{AAA,AAB,AAC,AAD,AAE,AAF,AAG,AAH,AAI,AAJ,AAK,AAL}, ZZI, WAM, IZZ); 
ram_4096x1 sinst_245(SHM,BHM,{ABA,ABB,ABC,ABD,ABE,ABF,ABG,ABH,ABI,ABJ,ABK,ABL}, ZZI, WBM, IZZ); 
ram_4096x1 sinst_246(SLM,BDM,{ACA,ACB,ACC,ACD,ACE,ACF,ACG,ACH,ACI,ACJ,ACK,ACL}, ZZI, WCM, IZZ); 
ram_4096x1 sinst_247(SDN,BDN,{aaa,aab,aac,aad,aae,aaf,aag,aah,aai,aaj,aak,aal}, ZZI, WAN, IZZ); 
ram_4096x1 sinst_248(SHN,BHN,{aba,abb,abc,abd,abe,abf,abg,abh,abi,abj,abk,abl}, ZZI, WBN, IZZ); 
ram_4096x1 sinst_249(SLN,BDN,{aca,acb,acc,acd,ace,acf,acg,ach,aci,acj,ack,acl}, ZZI, WCN, IZZ); 
ram_4096x1 sinst_250(SDO,BDO,{AEA,AEB,AEC,AED,AEE,AEF,AEG,AEH,AEI,AEJ,AEK,AEL}, ZZI, WAO, IZZ); 
ram_4096x1 sinst_251(SHO,BHO,{AFA,AFB,AFC,AFD,AFE,AFF,AFG,AFH,AFI,AFJ,AFK,AFL}, ZZI, WBO, IZZ); 
ram_4096x1 sinst_252(SLO,BDO,{AGA,AGB,AGC,AGD,AGE,AGF,AGG,AGH,AGI,AGJ,AGK,AGL}, ZZI, WCO, IZZ); 
ram_4096x1 sinst_253(SDP,BDP,{aea,aeb,aec,aed,aee,aef,aeg,aeh,aei,aej,aek,ael}, ZZI, WAP, IZZ); 
ram_4096x1 sinst_254(SHP,BHP,{afa,afb,afc,afd,afe,aff,afg,afh,afi,afj,afk,afl}, ZZI, WBP, IZZ); 
ram_4096x1 sinst_255(SLP,BDP,{aga,agb,agc,agd,age,agf,agg,agh,agi,agj,agk,agl}, ZZI, WCP, IZZ); 
endmodule;
