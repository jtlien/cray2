

module cpu_top(input sysclock,
               input         ihold, // just to prevent issue at 0
               input         iedataval,
               input         iedatahold,
               input [23:0]  quad0memparcel,
               input [23:0]  quad1memparcel,
               input [23:0]  quad2memparcel,
               input [23:0]  quad3memparcel,
               input [5:0]   quad0memdest,
               input [5:0]   quad1memdest,
               input [5:0]   quad2memdest,
               input [5:0]   quad3memdest,
	       input [1:0]   qd0release,
	       input [1:0]   qd1release,
	       input [1:0]   qd2release,
	       input [1:0]   qd3release,
	       input [7:0]   kaconsoletora,
	       input [31:0]  erroraddr,
               input [31:0]  tfbaseaddr,
               input  setbaseaddr,
	       input [19:0]  flooptoea,
	       output [4:0]  bankptrtoqb,
               output [23:0] quad0packet,
               output [23:0] quad1packet,
               output [23:0] quad2packet,
               output [23:0] quad3packet,
	       output [19:0] floopfrmeb,
               output [19:0] consoletonextra,
	       output        raloadbytenext,
               output [63:0] s2regval,
               output [31:0] a3regval
          );


   
wire enablecmrangetotf;
wire gaf0;
wire gaf1;
wire barreltesttoie;
wire branchpreambletoie;
wire branchintoie;
wire branchouttoie;
wire branchfallthrutoie;
wire fetchcmletetoif;
wire indlightlgoissue; 
wire ragatesqrthardround; 

 wire araddrtotf[0:31];
 wire ensignbit[0:8];
 wire enterbasetf;
 wire nxtcpup1blockref;
 wire nxtcpup2blockref;
 wire gatewdfromib;
 wire iolentoie[0:8];
 wire blockreftonext;
 wire goga;
 wire gaj0;
 wire gaj1;
 wire gak0;
   
 wire jafgacnt[0:1];
 wire jakgacnt;
 wire akshtogb[0:15];
 wire akshtovr[0:15];
 wire instpartoif[0:15];
 wire bankarivfromtf[0:2];
 wire stkbnd[0:1];
 wire enablebypass;
 wire stackboundary;
 wire clearreadadr;
 wire clearreadadr1;
 wire boundflagtotf;
 wire fetchcmpltoif;
 wire boundaryflagtoif;
 wire exchangedatafromjb[0:15];
 wire exchangedatafromja[0:15];
 wire sregbrdata[0:8];
 wire aregbrdata[0:8];
 wire barrelresp;
 wire boundaryseq;
 wire fetchinprog;
 wire goissueif[0:1];
 wire advanceqif;
 wire conflicktchain;
 wire semaphorefromea[0:2];
 wire deadstarttoif;
 wire enterpfromea;
 wire enterbafromea;
 wire enterlafromea;
 wire startfromea;
 wire enablecmrangetest;
 wire phasetoif;
 wire quad0bufferbusy;
 wire quad1bufferbusy;
 wire quad2bufferbusy;
 wire quad3bufferbusy;
 wire vlengthtoif[0:7];
 wire iolengthtoif[0:7];
 wire externalseq[0:2];
 wire refreshfromea;
 wire addresstota[0:31];
 wire ifcontroltota[0:24];
 wire gosdatatotb;
 wire goebdatatotb;
 wire retrytotb;
 wire brout[0:7];
 wire parcelptr[0:1];
 wire memportbusyfromif;
 wire holdissuefromif;
 wire gobranchfromif;
 wire semaphorefl_0[0:1];
 wire semaphorefl_1[0:1];
 wire semaphorefl_2[0:1];
 wire semaphorefl_3[0:1];
 wire setsematoea;
 wire clrsematoea;
 wire holdadvtojb1;
 wire holdadvtojb2;
 wire ifindlights[0:14];
 wire vectorshiftenable;
 wire enterardtowa;
 wire deadstartjc0;
 wire bcritetojc1[0:3];
 //wire phasefromjb;
 wire deadstartfromea;
 wire backupfromtf;
 wire phasetotd;
 wire enablesecded;
 wire validaddtotf;
 wire reproshtdata;
 wire refreshtotf;
 wire tfflagtolights[0:9];
 wire vectorenablefromjb;     

wire ltwaystation[0:15];
wire readparity;
wire fetcharrival[0:2];
wire fetcharrivaltoeb[0:2];
wire bankarrivfromtf[0:3];
wire ieindlights[0:23];
wire backupcnd[0:4];
wire validaddrtotf;
wire reproshfdata;
wire cmrangeerrortoea;
wire gatewdfromia;
wire blockreftonextp1;
wire blockreftonextp2;
wire blockreftonextp3;
wire refreshenblout;
wire functiondcdlights[0:7];
wire refreshenable;
wire nxtcpublockref;
wire nextcpup1blockref;
wire nextcpup2blockref;
wire phasetojb;
wire tailgatejb; 
wire shregdatajb[0:7];
wire adderselga;
wire addrtotc[0:31];
wire advanceqjb;
wire advlmadrtowa;
wire amtoar[0:31];
wire aradrtotf[0:31];
wire ardatatoincr;
wire aregsrctoar[0:5];
wire arfanouttojb[0:31];
wire arreadout[0:2];
wire arsigntest;
wire artoam[0:31];
wire artoas[0:7];
wire artofirstadder;
wire artoifviajb[0:31];
wire arzerotesta;
wire arzerotestb;
wire basetothirdaddr;
wire begvecttojc1[0:7];
wire begvecttojc0[0:7];
wire bp0mergetb1[0:4];
wire bp1mergetb1[0:4];
wire bp2mergetb1[0:4];
wire bp3mergetb1[0:4];
wire branchout;
wire branchpreamble;
wire bufferdataqd0;
wire bufferdataqd1;
wire bufferdataqd2;
wire bufferdataqd3;
wire bwritetojc0[0:3];
wire bwritetojc1[0:3];
wire carrietosecondaddr;
wire clearvectorlenvl;
wire clrsemaphore;
wire clrtoja[0:4];
wire cmdatatoeb[0:63];
wire cmdatatoie[0:63];
wire cmdesttoeb[0:63];
wire cmdesttoie[0:63];
wire coeftofb[0:47];
wire commemtovr[0:63];
wire commemtoeb[0:63];
wire commemtoie[0:63];
   
wire constoverflfc;
wire constreadwa;
wire constwritewa;
wire cunderflowtofc;
wire datareadyja;
wire deadstarteb;
wire deadstartia;
wire deadstartib;
wire deadstartie;
wire deadstartie1;
wire deadstartif;
wire deadstartjb;
wire deadstartjc1;
wire deadstartjc2;
wire deadstartqb;
wire deadstartra;
wire deadstarttc;
wire deadstartvl;
wire deadstrtja;
wire doublebiterror;
wire eaclock;
wire ebaddrtotf[0:31];
wire ebdatatb[0:63];
wire enablecmrangetest;
wire enablecmrangeea;
wire enablecmtoif;
wire enableexectoib;
wire enableexectoif;
wire enablefarangeerr;
wire enablefmrangeerr;
wire enableiota[0:1];
wire enablerangeerr;
wire enablerangerrfc;
wire endsequencetoeb;
wire enteradtowa;
wire enterbaseib;
wire enterbaseif;
wire enterbasetff;
wire enterlimitib;
wire enterlimitif;
wire enterlimittf;
wire enterltoar;
wire enterpib;
wire enterpif;
wire entervrtowa;
wire exittoea;
wire exptofc[0:16];
wire exterreftoib;
wire exterreftoif;
wire fbgoadd;
wire fbsubtractmode;
wire fctovr[0:63];
wire fetchcompletetoif;
wire flooptoeb[0:31];
wire fprangeerrfc;
wire fprangeerrme;
wire gathertest;
wire gatovr[0:63];
wire gbtovr[0:63];
wire goaddrmul;
wire goaddtofc;
wire gocons122174;
wire gocons123175;
wire goissuetoif[0:1];
wire goissuetojb[0:1];
wire goissuetojc0[0:1];
wire goissuetojc1[0:1];
wire goissuetowa[0:1];
wire goquadrant[0:3];
wire gosharedreg;
wire gostreamgb;
wire gowritetoeb;
wire hiwaterenable;
wire holdadvjc[0:1];
wire holdinincrement;
wire holdissueja;
wire holdissueic;
   
wire holdreadaddr;
wire holdtofirstaddr;
wire holdtosecondaddr;
wire ifaddrtotf[0:31];
wire ibinincrement;
wire ibufftoja[0:63];
wire idletoea;
wire ifinincrement;
wire indlightadvanceque;
wire indlightgateparcel[0:3];
wire indlightgoissue;
wire indlightrankcfull;
wire indlightrankefull;
wire incrtofirst;
wire incrtothirdaddr;
wire indlightip[0:31];
wire instbufadr[0:4];
wire instbufptr[0:9];
wire instpartoib[0:15];
wire instpartojb[0:15];
wire interrupttoib;
wire interrupttoif;
wire ioaddrtothirdaddr;
wire iolentoif[0:6];
wire jabranch;
wire jafacnt[0:4];
wire jagacnt[0:3];
wire jagbcnt[0:5];
wire jamecnt[0:5];
wire japarcel[0:1];
wire javacntr[0:3];
wire javbcntr[0:4];
wire javlcnt[0:6];
//wire jaarcntr[0:3];
wire jbatoar[0:31];
wire jbtovr[0:63];
wire jclocal[0:1];
wire jblengthlight[0:7];
wire jbindlight[0:5];
wire jkdatatoea[0:5];
wire jopfotoma[0:47];
wire jopfotomb[0:47];
wire jopfotomc[0:47];
wire jopfotomd[0:47];
wire kadeadstart;
wire kopfotoma[0:47];
wire kopfotomb[0:47];
wire kopfotomc[0:47];
wire kopfotomd[0:47];
wire lmaddrtoea[0:31];
wire lmadvancevec;
wire lmbanktoea[0:3];
wire lmbeginref;
wire lmparityea[0:7];
wire lmparityeafrvr[0:7];
   
wire lmwritemode;
wire looptofirstaddr;
wire ludatain[0:7];
wire lufotoma[0:9];
wire lufotomb[0:9];
wire lufotomc[0:31];
wire lufotomd[0:9];
wire luoddevenadd;
wire magatejdata;
wire magatekdata;
wire magatekdatadel;
wire magatekdatatoj;
wire maholdjdata;
wire mambflcar[0:15];
wire mambftlcar[0:15];
wire mambslcar[0:15];
wire mambtlcar[0:15];
wire marestomea[0:47];
wire marestomeb[0:47];
wire masellookup;
wire mbgatejdata;
wire mbgatekdata;
wire mbgatekdatadel;
wire mbgatekdatatoj;
wire mbholdjdata;
wire mbitercntl;
wire mbmcfitlcar[0:1];
wire mbmcflcar[0:13];
wire mbmcftlcar[0:1];
wire mbmcslcar[0:9];
wire mbmctlcar[0:5];
wire mbrestomea[0:9];
wire mbrestomeb[0:9];
wire mbrestomec[0:3];
wire mbsellookup;
wire mchardrnd[0:5];
wire rarndbit[0:1];
wire mcitercntl;
wire mcmdflcar[0:8];
wire mcmdftlcar[0:1];
wire mcmdslcar[0:7];
wire mcmdtlcar[0:3];
wire mcrestomea[0:12];
wire mcrestomeb[0:12];
wire mcrestomec[0:12];
wire mcsellookup;
wire mditercntl;
wire mdludata[0:14];
wire mdrestomea[0:27];
wire mdrestomeb[0:27];
wire mdrndbit[0:2];
wire mdsellookup;
wire mdselsqrtsh;
wire mefloatrnd;
wire mefuenable;
wire memarivtojc0[0:4];
wire memarivtojc1[0:4];
wire membackup0;
wire membackup2;
wire membackup3;
wire membsyja[0:1];
wire memdestcode[5:0];
wire memdestja[0:3];
wire mereciprnd;
wire mesqrtrnd;
wire metovr[0:63];
wire modechcnt[0:2];
wire newpregtoif[0:31];
wire normalizecnt12;
wire normalizecnt[0:5];
wire p0pktdata[0:23];
wire p1pktdata[0:23];
wire p2pktdata[0:23];
wire p3pktdata[0:23];
wire packreqq0[0:23];
wire packreqq1[0:23];
wire packreqq2[0:23];
wire packreqq3[0:23];
wire parceltowa[0:15];
wire phasejbtoas;
wire phasejbtocm[0:4];
wire phasejbtotm[0:5];
wire phasejbtonxtjb;
wire pkgphasetb;
wire pregtoam[0:31];
wire pregtoea[0:31];
wire qb0quadrela[0:1];
wire qb1quadrela[0:1];
wire qb2quadrela[0:1];
wire qb3quadrela[0:1];
wire rafourtyeight;
wire ragatejdata;
wire ragatekdata;
wire ragatekdatadel;
wire ragatekdatatoj;
wire ragaterecip;
wire ragatesqrt;
wire raholdjdata;
wire raloadbyte;
wire radeadstartnext;
wire raparityerror;
wire raselrecip;
wire readmodetoib;
wire readmodetoif;
wire recyclebd;
wire refreshinprog;
wire reliota[0:1];
wire relvitojb;
wire resumetoie;
wire rpacketquad0[0:23];
wire rpacketquad1[0:23];
wire rpacketquad2[0:23];
wire rpacketquad3[0:23];
wire scaldesttovr0[0:5];
wire scaldesttovr1[0:5];
wire scaldesttovr2[0:5];
wire scaldesttovr3[0:5];
wire scaldesttovr4[0:5];
wire scaldesttovr5[0:5];
wire scaldesttovr6[0:5];
wire scaldesttovr7[0:5];
wire scaljtovl[0:63];
wire scdatatoga[0:63];
wire sect0tofc[0:1];
wire sect1tofc[0:1];
wire sect2tofc[0:1];
wire selextdata;
wire selsidata;
wire semaphoreptr[0:2];
wire shdatatogb[0:63];
wire shftcnt[0:7];
wire shftcoef[0:47];
wire shftcoeflo;
wire shftcontogb[0:2];
wire shftovfl[0:2];
wire shifteqminus1;
wire shregoddeven;
wire shregtype1;
wire shregtype2;
wire shtambtovb[0:6];
wire shtovflvb;
wire signtofc[0:63];
wire singlebiterror;
wire sregsrctoam[0:5];
wire stackbndtotf;
wire stackmodetoib;
wire stackmodetoif;
wire subtracttoar;
wire addtoar;   
wire syndrome[0:7];
wire togglesign;
wire unlikesigns;
wire validsqrt;
wire v0addr1[0:5];
wire v0addr2[0:5];
wire v0addr3[0:5];
wire v0addr4[0:5];
wire v0addr5[0:5];
wire v0addr6[0:5];
wire v0addr7[0:5];
wire v0addr8[0:5];
wire v0vectmode[0:7];
wire v0vectstep[0:7];
wire v1addr1[0:5];
wire v1addr2[0:5];
wire v1addr3[0:5];
wire v1addr4[0:5];
wire v1addr5[0:5];
wire v1addr6[0:5];
wire v1addr7[0:5];
wire v1addr8[0:5];
wire v1vectmode[0:7];
wire v1vectstep[0:7];
wire v2addr1[0:5];
wire v2addr2[0:5];
wire v2addr3[0:5];
wire v2addr4[0:5];
wire v2addr5[0:5];
wire v2addr6[0:5];
wire v2addr7[0:5];
wire v2addr8[0:5];
wire v2vectmode[0:7];
wire v2vectstep[0:7];
wire v3addr1[0:5];
wire v3addr2[0:5];
wire v3addr3[0:5];
wire v3addr4[0:5];
wire v3addr5[0:5];
wire v3addr6[0:5];
wire v3addr7[0:5];
wire v3addr8[0:5];
wire v3vectmode[0:7];
wire v3vectstep[0:7];
wire v4addr1[0:5];
wire v4addr2[0:5];
wire v4addr3[0:5];
wire v4addr4[0:5];
wire v4addr5[0:5];
wire v4addr6[0:5];
wire v4addr7[0:5];
wire v4addr8[0:5];
wire v4vectmode[0:7];
wire v4vectstep[0:7];
wire v5addr1[0:5];
wire v5addr2[0:5];
wire v5addr3[0:5];
wire v5addr4[0:5];
wire v5addr5[0:5];
wire v5addr6[0:5];
wire v5addr7[0:5];
wire v5addr8[0:5];
wire v5vectmode[0:7];
wire v5vectstep[0:7];
wire v6addr1[0:5];
wire v6addr2[0:5];
wire v6addr3[0:5];
wire v6addr4[0:5];
wire v6addr5[0:5];
wire v6addr6[0:5];
wire v6addr7[0:5];
wire v6addr8[0:5];
wire v6vectmode[0:7];
wire v6vectstep[0:7];
wire v7addr1[0:5];
wire v7addr2[0:5];
wire v7addr3[0:5];
wire v7addr4[0:5];
wire v7addr5[0:5];
wire v7addr6[0:5];
wire v7addr7[0:5];
wire v7addr8[0:5];
wire v7vectmode[0:7];
wire v7vectstep[0:7];
wire vasregsign;
   
wire vasregzero[0:7];
wire vatovb[0:63];
wire vbtovr[0:63];
wire vec0rel;
wire vec1rel;
wire vec2rel;
wire vec3rel;
wire vec4rel;
wire vec5rel;
wire vec6rel;
wire vec7rel;
wire vectlentoam[0:5];
wire vectlentoib[0:5];
wire vectlentoif[0:5];
wire vectlentojb[0:5];
wire vectlentojc0[0:5];
wire vectlentojc1[0:5];
wire vector1srccode[0:6];
wire vector2srccode[0:6];
wire vector3srccode[0:6];
wire vector4srccode[0:6];
wire vector5srccode[0:6];
wire vector6srccode[0:6];
wire vector7srccode[0:6];
wire vector8srccode[0:6];
wire vectorcodeam[0:6];
wire vectorlencntl;
wire vectormode[0:1];
wire vltovr[0:63];
wire vraddrtotf[0:31];
wire vrdatatb[0:63];
wire vrdatatbrel[0:63];
wire vrtoar[0:63];
wire vrtofaj[0:63];
wire vrtofak[0:63];
wire vrtolm[0:63];
wire vrtocm[0:63];
wire vrtomulj[0:63];
wire vrtomulk[0:63];
wire vrtosecondadder;
wire vrtovaj[0:63];
wire vrtovak[0:63];
wire vrtovb[0:63];
wire vrtovlk[0:63];
wire wadatalm[0:63];
wire watoar[0:63];
wire watovr[0:63];      
wire raintoranxt[0:7];
wire wajamecnt[0:5];
wire mccotwoseven;
   

                         
assign memdestcode[0] = ifcontroltota[0];
assign memdestcode[1] = ifcontroltota[1];
assign memdestcode[2] = ifcontroltota[2];
assign memdestcode[3] = ifcontroltota[3];
assign memdestcode[4] = ifcontroltota[4];
assign memdestcode[5] = ifcontroltota[5];
   
assign validaddtotf = ifcontroltota[6];
assign reproshtdata = ifcontroltota[7];
assign enablecmrangetotf = ifcontroltota[8];
assign gathertest = ifcontroltota[10];
//assign phasejbtotm[0] = ifcontroltota[11];
assign incrtofirst = ifcontroltota[11];
assign artofirstadder = ifcontroltota[12];
//assign looptofirstaddr = ifcontroltota[13];
assign holdtofirstaddr = ifcontroltota[13];
assign vrtosecondadder = ifcontroltota[14];
assign carrietosecondaddr = ifcontroltota[15];
assign holdtosecondaddr = ifcontroltota[16];
assign ioaddrtothirdaddr = ifcontroltota[17];
assign incrtothirdaddr = ifcontroltota[18];
assign basetothirdaddr = ifcontroltota[19];
assign ardatatoincr = ifcontroltota[20];
assign ifinincrement = ifcontroltota[21];
assign holdinincrement = ifcontroltota[22];
assign enterbasetf = ifcontroltota[23];
assign enterlimittf = ifcontroltota[24];

am am0 (
.IAA(artoam[0]),
.IAB(artoam[1]),
.IAC(artoam[2]),
.IAD(artoam[3]),
.IAE(artoam[4]),
.IAF(artoam[5]),
.IAG(artoam[6]),
.IAH(artoam[7]),
.IAI(artoam[8]),
.IAJ(artoam[9]),
.IAK(artoam[10]),
.IAL(artoam[11]),
.IAM(artoam[12]),
.IAN(artoam[13]),
.IAO(artoam[14]),
.IAP(artoam[15]),
.IBA(artoam[16]),
.IBB(artoam[17]),
.IBC(artoam[18]),
.IBD(artoam[19]),
.IBE(artoam[20]),
.IBF(artoam[21]),
.IBG(artoam[22]),
.IBH(artoam[23]),
.IBI(artoam[24]),
.IBJ(artoam[25]),
.IBK(artoam[26]),
.IBL(artoam[27]),
.IBM(artoam[28]),
.IBN(artoam[29]),
.IBO(artoam[30]),
.IBP(artoam[31]),
.ICA(pregtoam[0]),
.ICB(pregtoam[1]),
.ICC(pregtoam[2]),
.ICD(pregtoam[3]),
.ICE(pregtoam[4]),
.ICF(pregtoam[5]),
.ICG(pregtoam[6]),
.ICH(pregtoam[7]),
.ICI(pregtoam[8]),
.ICJ(pregtoam[9]),
.ICK(pregtoam[10]),
.ICL(pregtoam[11]),
.ICM(pregtoam[12]),
.ICN(pregtoam[13]),
.ICO(pregtoam[14]),
.ICP(pregtoam[15]),
.IDA(pregtoam[16]),
.IDB(pregtoam[17]),
.IDC(pregtoam[18]),
.IDD(pregtoam[19]),
.IDE(pregtoam[20]),
.IDF(pregtoam[21]),
.IDG(pregtoam[22]),
.IDH(pregtoam[23]),
.IDI(pregtoam[24]),
.IDJ(pregtoam[25]),
.IDK(pregtoam[26]),
.IDL(pregtoam[27]),
.IDM(pregtoam[28]),
.IDN(pregtoam[29]),
.IDO(pregtoam[30]),
.IDP(pregtoam[31]),
.IEA(vectlentoam[0]),
.IEB(vectlentoam[1]),
.IEC(vectlentoam[2]),
.IED(vectlentoam[3]),
.IEE(vectlentoam[4]),
.IEF(vectlentoam[5]),
.IFA(vectorcodeam[0]),
.IFB(vectorcodeam[1]),
.IFC(vectorcodeam[2]),
.IFD(vectorcodeam[3]),
.IFE(vectorcodeam[4]),
.IFFF(vectorcodeam[5]),
.IFG(vectorcodeam[6]),
.IGA(sregsrctoam[0]),
.IGB(sregsrctoam[1]),
.IGC(sregsrctoam[2]),
.IGD(sregsrctoam[3]),
.IGE(sregsrctoam[4]),
.IGF(sregsrctoam[5]),
.IHA(goaddrmul),
.IZZ(sysclock),
.IZH(ihold),
.OAA(amtoar[0]),
.OAB(amtoar[1]),
.OAC(amtoar[2]),
.OAD(amtoar[3]),
.OAE(amtoar[4]),
.OAF(amtoar[5]),
.OAG(amtoar[6]),
.OAH(amtoar[7]),
.OAI(amtoar[8]),
.OAJ(amtoar[9]),
.OAK(amtoar[10]),
.OAL(amtoar[11]),
.OAM(amtoar[12]),
.OAN(amtoar[13]),
.OAO(amtoar[14]),
.OAP(amtoar[15]),
.OBA(amtoar[16]),
.OBB(amtoar[17]),
.OBC(amtoar[18]),
.OBD(amtoar[19]),
.OBE(amtoar[20]),
.OBF(amtoar[21]),
.OBG(amtoar[22]),
.OBH(amtoar[23]),
.OBI(amtoar[24]),
.OBJ(amtoar[25]),
.OBK(amtoar[26]),
.OBL(amtoar[27]),
.OBM(amtoar[28]),
.OBN(amtoar[29]),
.OBO(amtoar[30]),
.OBP(amtoar[31]),
.OCA(pregtoea[0]),
.OCB(pregtoea[1]),
.OCC(pregtoea[2]),
.OCD(pregtoea[3]),
.OCE(pregtoea[4]),
.OCF(pregtoea[5]),
.OCG(pregtoea[6]),
.OCH(pregtoea[7]),
.OCI(pregtoea[8]),
.OCJ(pregtoea[9]),
.OCK(pregtoea[10]),
.OCL(pregtoea[11]),
.OCM(pregtoea[12]),
.OCN(pregtoea[13]),
.OCO(pregtoea[14]),
.OCP(pregtoea[15]),
.ODA(pregtoea[16]),
.ODB(pregtoea[17]),
.ODC(pregtoea[18]),
.ODD(pregtoea[19]),
.ODE(pregtoea[20]),
.ODF(pregtoea[21]),
.ODG(pregtoea[22]),
.ODH(pregtoea[23]),
.ODI(pregtoea[24]),
.ODJ(pregtoea[25]),
.ODK(pregtoea[26]),
.ODL(pregtoea[27]),
.ODM(pregtoea[28]),
.ODN(pregtoea[29]),
.ODO(pregtoea[30]),
.ODP(pregtoea[31]),
.OEA(vectlentoif[0]),
.OEB(vectlentoif[1]),
.OEC(vectlentoif[2]),
.OED(vectlentoif[3]),
.OEE(vectlentoif[4]),
.OEF(vectlentoif[5]),
.OFA(vectlentojb[0]),
.OFB(vectlentojb[1]),
.OFC(vectlentojb[2]),
.OFD(vectlentojb[3]),
.OFE(vectlentojb[4]),
.OFF(vectlentojb[5]),
.OGA(vectlentojc0[0]),
.OGB(vectlentojc0[1]),
.OGC(vectlentojc0[2]),
.OGD(vectlentojc0[3]),
.OGE(vectlentojc0[4]),
.OGF(vectlentojc0[5]),
.OHA(vectlentojc1[0]),
.OHB(vectlentojc1[1]),
.OHC(vectlentojc1[2]),
.OHD(vectlentojc1[3]),
.OHE(vectlentojc1[4]),
.OHF(vectlentojc1[5]),
.OIA(vector1srccode[0]),
.OIB(vector1srccode[1]),
.OIC(vector1srccode[2]),
.OID(vector1srccode[3]),
.OIE(vector1srccode[4]),
.OIF(vector1srccode[5]),
.OIG(vector1srccode[6]),
.OIH(scaldesttovr0[0]),
.OII(scaldesttovr0[1]),
.OIJ(scaldesttovr0[2]),
.OIK(scaldesttovr0[3]),
.OIL(scaldesttovr0[4]),
.OIM(scaldesttovr0[5]),
.OJA(vector2srccode[0]),
.OJB(vector2srccode[1]),
.OJC(vector2srccode[2]),
.OJD(vector2srccode[3]),
.OJE(vector2srccode[4]),
.OJF(vector2srccode[5]),
.OJG(vector2srccode[6]),
.OJH(scaldesttovr1[0]),
.OJI(scaldesttovr1[1]),
.OJJ(scaldesttovr1[2]),
.OJK(scaldesttovr1[3]),
.OJL(scaldesttovr1[4]),
.OJM(scaldesttovr1[5]),
.OKA(vector3srccode[0]),
.OKB(vector3srccode[1]),
.OKC(vector3srccode[2]),
.OKD(vector3srccode[3]),
.OKE(vector3srccode[4]),
.OKF(vector3srccode[5]),
.OKG(vector3srccode[6]),
.OKH(scaldesttovr2[0]),
.OKI(scaldesttovr2[1]),
.OKJ(scaldesttovr2[2]),
.OKK(scaldesttovr2[3]),
.OKL(scaldesttovr2[4]),
.OKM(scaldesttovr2[5]),
.OLA(vector4srccode[0]),
.OLB(vector4srccode[1]),
.OLC(vector4srccode[2]),
.OLD(vector4srccode[3]),
.OLE(vector4srccode[4]),
.OLF(vector4srccode[5]),
.OLG(vector4srccode[6]),
.OLH(scaldesttovr3[0]),
.OLI(scaldesttovr3[1]),
.OLJ(scaldesttovr3[2]),
.OLK(scaldesttovr3[3]),
.OLL(scaldesttovr3[4]),
.OLM(scaldesttovr3[5]),
.OMA(vector5srccode[0]),
.OMB(vector5srccode[1]),
.OMC(vector5srccode[2]),
.OMD(vector5srccode[3]),
.OME(vector5srccode[4]),
.OMF(vector5srccode[5]),
.OMG(vector5srccode[6]),
.OMH(scaldesttovr4[0]),
.OMI(scaldesttovr4[1]),
.OMJ(scaldesttovr4[2]),
.OMK(scaldesttovr4[3]),
.OML(scaldesttovr4[4]),
.OMM(scaldesttovr4[5]),
.ONA(vector6srccode[0]),
.ONB(vector6srccode[1]),
.ONC(vector6srccode[2]),
.OND(vector6srccode[3]),
.ONE(vector6srccode[4]),
.ONF(vector6srccode[5]),
.ONG(vector6srccode[6]),
.ONH(scaldesttovr5[0]),
.ONI(scaldesttovr5[1]),
.ONJ(scaldesttovr5[2]),
.ONK(scaldesttovr5[3]),
.ONL(scaldesttovr5[4]),
.ONM(scaldesttovr5[5]),
.OOA(vector7srccode[0]),
.OOB(vector7srccode[1]),
.OOC(vector7srccode[2]),
.OOD(vector7srccode[3]),
.OOE(vector7srccode[4]),
.OOF(vector7srccode[5]),
.OOG(vector7srccode[6]),
.OOH(scaldesttovr6[0]),
.OOI(scaldesttovr6[1]),
.OOJ(scaldesttovr6[2]),
.OOK(scaldesttovr6[3]),
.OOL(scaldesttovr6[4]),
.OOM(scaldesttovr6[5]),
.OPA(vector8srccode[0]),
.OPB(vector8srccode[1]),
.OPC(vector8srccode[2]),
.OPD(vector8srccode[3]),
.OPE(vector8srccode[4]),
.OPF(vector8srccode[5]),
.OPG(vector8srccode[6]),
.OPH(scaldesttovr7[0]),
.OPI(scaldesttovr7[1]),
.OPJ(scaldesttovr7[2]),
.OPK(scaldesttovr7[3]),
.OPL(scaldesttovr7[4]),
.OPM(scaldesttovr7[5])
);
  
ar ar0 (
.IAA(watoar[0]),
.IAB(watoar[1]),
.IAC(watoar[2]),
.IAD(watoar[3]),
.IAE(watoar[4]),
.IAF(watoar[5]),
.IAG(watoar[6]),
.IAH(watoar[7]),
.IAI(watoar[8]),
.IAJ(watoar[9]),
.IAK(watoar[10]),
.IAL(watoar[11]),
.IAM(watoar[12]),
.IAN(watoar[13]),
.IAO(watoar[14]),
.IAP(watoar[15]),
.IBA(watoar[16]),
.IBB(watoar[17]),
.IBC(watoar[18]),
.IBD(watoar[19]),
.IBE(watoar[20]),
.IBF(watoar[21]),
.IBG(watoar[22]),
.IBH(watoar[23]),
.IBI(watoar[24]),
.IBJ(watoar[25]),
.IBK(watoar[26]),
.IBL(watoar[27]),
.IBM(watoar[28]),
.IBN(watoar[29]),
.IBO(watoar[30]),
.IBP(watoar[31]),
.ICA(vrtoar[0]),
.ICB(vrtoar[1]),
.ICC(vrtoar[2]),
.ICD(vrtoar[3]),
.ICE(vrtoar[4]),
.ICF(vrtoar[5]),
.ICG(vrtoar[6]),
.ICH(vrtoar[7]),
.ICI(vrtoar[8]),
.ICJ(vrtoar[9]),
.ICK(vrtoar[10]),
.ICL(vrtoar[11]),
.ICM(vrtoar[12]),
.ICN(vrtoar[13]),
.ICO(vrtoar[14]),
.ICP(vrtoar[15]),
.IDA(vrtoar[16]),
.IDB(vrtoar[17]),
.IDC(vrtoar[18]),
.IDD(vrtoar[19]),
.IDE(vrtoar[20]),
.IDF(vrtoar[21]),
.IDG(vrtoar[22]),
.IDH(vrtoar[23]),
.IDI(vrtoar[24]),
.IDJ(vrtoar[25]),
.IDK(vrtoar[26]),
.IDL(vrtoar[27]),
.IDM(vrtoar[28]),
.IDN(vrtoar[29]),
.IDO(vrtoar[30]),
.IDP(vrtoar[31]),
.IEA(jbatoar[0]),
.IEB(jbatoar[1]),
.IEC(jbatoar[2]),
.IED(jbatoar[3]),
.IEE(jbatoar[4]),
.IEF(jbatoar[5]),
.IEG(jbatoar[6]),
.IEH(jbatoar[7]),
.IEI(jbatoar[8]),
.IEJ(jbatoar[9]),
.IEK(jbatoar[10]),
.IEL(jbatoar[11]),
.IEM(jbatoar[12]),
.IEN(jbatoar[13]),
.IEO(jbatoar[14]),
.IEP(jbatoar[15]),
.IFA(jbatoar[16]),
.IFB(jbatoar[17]),
.IFC(jbatoar[18]),
.IFD(jbatoar[19]),
.IFE(jbatoar[20]),
.IFFF(jbatoar[21]),
.IFG(jbatoar[22]),
.IFH(jbatoar[23]),
.IFI(jbatoar[24]),
.IFJ(jbatoar[25]),
.IFK(jbatoar[26]),
.IFL(jbatoar[27]),
.IFM(jbatoar[28]),
.IFN(jbatoar[29]),
.IFO(jbatoar[30]),
.IFP(jbatoar[31]),
.IGA(amtoar[0]),
.IGB(amtoar[1]),
.IGC(amtoar[2]),
.IGD(amtoar[3]),
.IGE(amtoar[4]),
.IGF(amtoar[5]),
.IGG(amtoar[6]),
.IGH(amtoar[7]),
.IGI(amtoar[8]),
.IGJ(amtoar[9]),
.IGK(amtoar[10]),
.IGL(amtoar[11]),
.IGM(amtoar[12]),
.IGN(amtoar[13]),
.IGO(amtoar[14]),
.IGP(amtoar[15]),
.IHA(amtoar[16]),
.IHB(amtoar[17]),
.IHC(amtoar[18]),
.IHD(amtoar[19]),
.IHE(amtoar[20]),
.IHF(amtoar[21]),
.IHG(amtoar[22]),
.IHH(amtoar[23]),
.IHI(amtoar[24]),
.IHJ(amtoar[25]),
.IHK(amtoar[26]),
.IHL(amtoar[27]),
.IHM(amtoar[28]),
.IHN(amtoar[29]),
.IHO(amtoar[30]),
.IHP(amtoar[31]),
.IIA(arreadout[0]),
.IIB(arreadout[1]),
.IIC(arreadout[2]),
.IJA(aregsrctoar[0]),
.IJB(aregsrctoar[1]),
.IJC(aregsrctoar[2]),
.IJD(aregsrctoar[3]),
.IJE(aregsrctoar[4]),
.IJF(aregsrctoar[5]),
.IKA(subtracttoar),
.IKB(addtoar),
.ILA(enterltoar),
.IMA(),
.IZZ (sysclock),
.OAA(wadatalm[0]),
.OAB(wadatalm[1]),
.OAC(wadatalm[2]),
.OAD(wadatalm[3]),
.OAE(wadatalm[4]),
.OAF(wadatalm[5]),
.OAG(wadatalm[6]),
.OAH(wadatalm[7]),
.OAI(wadatalm[8]),
.OAJ(wadatalm[9]),
.OAK(wadatalm[10]),
.OAL(wadatalm[11]),
.OAM(wadatalm[12]),
.OAN(wadatalm[13]),
.OAO(wadatalm[14]),
.OAP(wadatalm[15]),
.OBA(wadatalm[16]),
.OBB(wadatalm[17]),
.OBC(wadatalm[18]),
.OBD(wadatalm[19]),
.OBE(wadatalm[20]),
.OBF(wadatalm[21]),
.OBG(wadatalm[22]),
.OBH(wadatalm[23]),
.OBI(wadatalm[24]),
.OBJ(wadatalm[25]),
.OBK(wadatalm[26]),
.OBL(wadatalm[27]),
.OBM(wadatalm[28]),
.OBN(wadatalm[29]),
.OBO(wadatalm[30]),
.OBP(wadatalm[31]),
.OCA(araddrtotf[0]),
.OCB(araddrtotf[1]),
.OCC(araddrtotf[2]),
.OCD(araddrtotf[3]),
.OCE(araddrtotf[4]),
.OCF(araddrtotf[5]),
.OCG(araddrtotf[6]),
.OCH(araddrtotf[7]),
.OCI(araddrtotf[8]),
.OCJ(araddrtotf[9]),
.OCK(araddrtotf[10]),
.OCL(araddrtotf[11]),
.OCM(araddrtotf[12]),
.OCN(araddrtotf[13]),
.OCO(araddrtotf[14]),
.OCP(araddrtotf[15]),
.ODA(araddrtotf[16]),
.ODB(araddrtotf[17]),
.ODC(araddrtotf[18]),
.ODD(araddrtotf[19]),
.ODE(araddrtotf[20]),
.ODF(araddrtotf[21]),
.ODG(araddrtotf[22]),
.ODH(araddrtotf[23]),
.ODI(araddrtotf[24]),
.ODJ(araddrtotf[25]),
.ODK(araddrtotf[26]),
.ODL(araddrtotf[27]),
.ODM(araddrtotf[28]),
.ODN(araddrtotf[29]),
.ODO(araddrtotf[30]),
.ODP(araddrtotf[31]),
.OEA(arfanouttojb[0]),
.OEB(arfanouttojb[1]),
.OEC(arfanouttojb[2]),
.OED(arfanouttojb[3]),
.OEE(arfanouttojb[4]),
.OEF(arfanouttojb[5]),
.OEG(arfanouttojb[6]),
.OEH(arfanouttojb[7]),
.OEI(arfanouttojb[8]),
.OEJ(arfanouttojb[9]),
.OEK(arfanouttojb[10]),
.OEL(arfanouttojb[11]),
.OEM(arfanouttojb[12]),
.OEN(arfanouttojb[13]),
.OEO(arfanouttojb[14]),
.OEP(arfanouttojb[15]),
.OFA(arfanouttojb[16]),
.OFB(arfanouttojb[17]),
.OFC(arfanouttojb[18]),
.OFD(arfanouttojb[19]),
.OFE(arfanouttojb[20]),
.OFF(arfanouttojb[21]),
.OFG(arfanouttojb[22]),
.OFH(arfanouttojb[23]),
.OFI(arfanouttojb[24]),
.OFJ(arfanouttojb[25]),
.OFK(arfanouttojb[26]),
.OFL(arfanouttojb[27]),
.OFM(arfanouttojb[28]),
.OFN(arfanouttojb[29]),
.OFO(arfanouttojb[30]),
.OFP(arfanouttojb[31]),
.OGA(artoam[0]),
.OGB(artoam[1]),
.OGC(artoam[2]),
.OGD(artoam[3]),
.OGE(artoam[4]),
.OGF(artoam[5]),
.OGG(artoam[6]),
.OGH(artoam[7]),
.OGI(artoam[8]),
.OGJ(artoam[9]),
.OGK(artoam[10]),
.OGL(artoam[11]),
.OGM(artoam[12]),
.OGN(artoam[13]),
.OGO(artoam[14]),
.OGP(artoam[15]),
.OHA(artoam[16]),
.OHB(artoam[17]),
.OHC(artoam[18]),
.OHD(artoam[19]),
.OHE(artoam[20]),
.OHF(artoam[21]),
.OHG(artoam[22]),
.OHH(artoam[23]),
.OHI(artoam[24]),
.OHJ(artoam[25]),
.OHK(artoam[26]),
.OHL(artoam[27]),
.OHM(artoam[28]),
.OHN(artoam[29]),
.OHO(artoam[30]),
.OHP(artoam[31]),
.OIA(shftcnt[0]),
.OIB(shftcnt[1]),
.OIC(shftcnt[2]),
.OID(shftcnt[3]),
.OIE(shftcnt[4]),
.OIF(shftcnt[5]),
.OIG(shftcnt[6]),
.OIH(shftovfl[0]),
.OIJ(shftovfl[2]),
.OJA(vectlentoam[0]),
.OJB(vectlentoam[1]),
.OJC(vectlentoam[2]),
.OJD(vectlentoam[3]),
.OJE(vectlentoam[4]),
.OJF(vectlentoam[5]),
.OKA(arzerotesta),
.OKB(arzerotestb),
.OKC(arsigntest),
.OMA(ensignbit[0]),
.OMB(ensignbit[1]),
.OMC(ensignbit[2]),
.OMD(ensignbit[3]),
.OME(ensignbit[4]),
.OMF(ensignbit[5]),
.OMG(ensignbit[6]),
.OMH(ensignbit[7]));
  
ea ea0 (
.IAA(pregtoea[0]),
.IAB(pregtoea[1]),
.IAC(pregtoea[2]),
.IAD(pregtoea[3]),
.IAE(pregtoea[4]),
.IAF(pregtoea[5]),
.IAG(pregtoea[6]),
.IAH(pregtoea[7]),
.IAI(pregtoea[8]),
.IAJ(pregtoea[9]),
.IAK(pregtoea[10]),
.IAL(pregtoea[11]),
.IAM(pregtoea[12]),
.IAN(pregtoea[13]),
.IAO(pregtoea[14]),
.IAP(pregtoea[15]),
.IBA(pregtoea[16]),
.IBB(pregtoea[17]),
.IBC(pregtoea[18]),
.IBD(pregtoea[19]),
.IBE(pregtoea[20]),
.IBF(pregtoea[21]),
.IBG(pregtoea[22]),
.IBH(pregtoea[23]),
.IBI(pregtoea[24]),
.IBJ(pregtoea[25]),
.IBK(pregtoea[26]),
.IBL(pregtoea[27]),
.IBM(pregtoea[28]),
.IBN(pregtoea[29]),
.IBO(pregtoea[30]),
.IBP(pregtoea[31]),
.ICA(flooptoea[0]),
.ICB(flooptoea[1]),
.ICC(flooptoea[2]),
.ICD(flooptoea[3]),
.ICE(flooptoea[4]),
.ICF(flooptoea[5]),
.ICG(flooptoea[6]),
.ICH(flooptoea[7]),
.ICI(flooptoea[8]),
.ICJ(flooptoea[9]),
.ICK(flooptoea[10]),
.ICL(flooptoea[11]),
.ICM(flooptoea[12]),
.ICN(flooptoea[13]),
.ICO(flooptoea[14]),
.ICP(flooptoea[15]),
.ICQ(flooptoea[16]),
.ICR(flooptoea[17]),
.ICS(flooptoea[18]),
.ICT(flooptoea[19]),
.IDA(jkdatatoea[0]),
.IDB(jkdatatoea[1]),
.IDC(jkdatatoea[2]),
.IDD(jkdatatoea[3]),
.IDE(jkdatatoea[4]),
.IDF(jkdatatoea[5]),
.IEA(setsematoea),
.IEB(clrsematoea),
.IEC(idletoea),
.IED(exittoea),
.IEE(),
.IEF(cmrangeerrortoea),
.IEG(hiwaterenable),
.IFA(fprangeerrfc),
.IFB(fprangeerrme),
.IFC(),
.IFD(raparityerror),
.IGA(kadeadstart),
.IHA(modechcnt[0]),
.IHB(modechcnt[1]),
.IHC(modechcnt[2]),
.IIA(lmbeginref),
.IIB(lmwritemode),
.IIC(lmadvancevec),
.IJA(lmbanktoea[0]),
.IJB(lmbanktoea[1]),
.IJC(lmbanktoea[2]),
.IJD(lmbanktoea[3]),
.IKA(lmaddrtoea[0]),
.IKB(lmaddrtoea[1]),
.IKC(lmaddrtoea[2]),
.IKD(lmaddrtoea[3]),
.IKE(lmaddrtoea[4]),
.IKF(lmaddrtoea[5]),
.IKG(lmaddrtoea[6]),
.IKH(lmaddrtoea[7]),
.IKI(lmaddrtoea[8]),
.IKJ(lmaddrtoea[9]),
.IKK(lmaddrtoea[10]),
.IKL(lmaddrtoea[11]),
.ILA(lmparityea[0]),
.ILB(lmparityea[1]),
.ILC(lmparityea[2]),
.ILD(lmparityea[3]),
.ILE(lmparityea[4]),
.ILF(lmparityea[5]),
.ILG(lmparityea[6]),
.ILH(lmparityea[7]),
.IMA(lmparityeafrvr[0]),
.IMB(lmparityeafrvr[1]),
.IMC(lmparityeafrvr[2]),
.IMD(lmparityeafrvr[3]),
.IME(lmparityeafrvr[4]),
.IMF(lmparityeafrvr[5]),
.IMG(lmparityeafrvr[6]),
.IMH(lmparityeafrvr[7]),
.IXA(eaclock),
.IZZ (sysclock),
.OHA(newpregtoif[0]),
.OHB(newpregtoif[1]),
.OHC(newpregtoif[2]),
.OHD(newpregtoif[3]),
.OHE(newpregtoif[4]),
.OHF(newpregtoif[5]),
.OHG(newpregtoif[6]),
.OHH(newpregtoif[7]),
.OHI(newpregtoif[8]),
.OHJ(newpregtoif[9]),
.OHK(newpregtoif[10]),
.OHL(newpregtoif[11]),
.OHM(newpregtoif[12]),
.OHN(newpregtoif[13]),
.OHO(newpregtoif[14]),
.OHP(newpregtoif[15]),
.OIA(newpregtoif[16]),
.OIB(newpregtoif[17]),
.OIC(newpregtoif[18]),
.OID(newpregtoif[19]),
.OIE(newpregtoif[20]),
.OIF(newpregtoif[21]),
.OIG(newpregtoif[22]),
.OIH(newpregtoif[23]),
.OII(newpregtoif[24]),
.OIJ(newpregtoif[25]),
.OIK(newpregtoif[26]),
.OIL(newpregtoif[27]),
.OIM(newpregtoif[28]),
.OIN(newpregtoif[29]),
.OIO(newpregtoif[30]),
.OIP(newpregtoif[31]),
.OJA(deadstrtja),
.OJB(deadstartjb),
.OJC(deadstartjc1),
.OJD(deadstartjc2),
.OJE(deadstarteb),
.OJF(deadstartqb),
.OJG(deadstartvl),
.OJH(deadstarttc),
.OJI(deadstartie),
.OJJ(deadstartif),
.OJK(deadstartra),
.OJL(deadstartie1),
.OKA(flooptoeb[0]),
.OKB(flooptoeb[1]),
.OKC(flooptoeb[2]),
.OKD(flooptoeb[3]),
.OKE(flooptoeb[4]),
.OKF(flooptoeb[5]),
.OKG(flooptoeb[6]),
.OKH(flooptoeb[7]),
.OKI(flooptoeb[8]),
.OKJ(flooptoeb[9]),
.OKK(flooptoeb[10]),
.OKL(flooptoeb[11]),
.OKM(flooptoeb[12]),
.OKN(flooptoeb[13]),
.OKO(flooptoeb[14]),
.OKP(flooptoeb[15]),
.OKQ(flooptoeb[16]),
.OKR(flooptoeb[17]),
.OKS(flooptoeb[18]),
.OKT(flooptoeb[19]),
.OLA(semaphoreptr[0]),
.OLB(semaphoreptr[1]),
.OLC(semaphoreptr[2]),
.OMA(interrupttoif),
.OMB(enterpfromea),
.OMC(enterbafromea),
.OMD(enterlafromea),
.OME(enablecmtoif),
.OMF(stackmodetoif),
.ONA(enablefmrangeerr),
.ONB(enablefarangeerr),
.OOA(enablecmrangetest));
   

  
eb eb0 (
.IAA(commemtoeb[0]),
.IAB(commemtoeb[1]),
.IAC(commemtoeb[2]),
.IAD(commemtoeb[3]),
.IAE(commemtoeb[4]),
.IAF(commemtoeb[5]),
.IAG(commemtoeb[6]),
.IAH(commemtoeb[7]),
.IAI(commemtoeb[8]),
.IAJ(commemtoeb[9]),
.IAK(commemtoeb[10]),
.IAL(commemtoeb[11]),
.IAM(commemtoeb[12]),
.IAN(commemtoeb[13]),
.IAO(commemtoeb[14]),
.IAP(commemtoeb[15]),
.IBA(commemtoeb[16]),
.IBB(commemtoeb[17]),
.IBC(commemtoeb[18]),
.IBD(commemtoeb[19]),
.IBE(commemtoeb[20]),
.IBF(commemtoeb[21]),
.IBG(commemtoeb[22]),
.IBH(commemtoeb[23]),
.IBI(commemtoeb[24]),
.IBJ(commemtoeb[25]),
.IBK(commemtoeb[26]),
.IBL(commemtoeb[27]),
.IBM(commemtoeb[28]),
.IBN(commemtoeb[29]),
.IBO(commemtoeb[30]),
.IBP(commemtoeb[31]),
.ICA(commemtoeb[32]),
.ICB(commemtoeb[33]),
.ICC(commemtoeb[34]),
.ICD(commemtoeb[35]),
.ICE(commemtoeb[36]),
.ICF(commemtoeb[37]),
.ICG(commemtoeb[38]),
.ICH(commemtoeb[39]),
.ICI(commemtoeb[40]),
.ICJ(commemtoeb[41]),
.ICK(commemtoeb[42]),
.ICL(commemtoeb[43]),
.ICM(commemtoeb[44]),
.ICN(commemtoeb[45]),
.ICO(commemtoeb[46]),
.ICP(commemtoeb[47]),
.IDA(commemtoeb[48]),
.IDB(commemtoeb[49]),
.IDC(commemtoeb[50]),
.IDD(commemtoeb[51]),
.IDE(commemtoeb[52]),
.IDF(commemtoeb[53]),
.IDG(commemtoeb[54]),
.IDH(commemtoeb[55]),
.IDI(commemtoeb[56]),
.IDJ(commemtoeb[57]),
.IDK(commemtoeb[58]),
.IDL(commemtoeb[59]),
.IDM(commemtoeb[60]),
.IDN(commemtoeb[61]),
.IDO(commemtoeb[62]),
.IDP(commemtoeb[63]),
.IEA(erroraddr[0]),
.IEB(erroraddr[1]),
.IEC(erroraddr[2]),
.IED(erroraddr[3]),
.IEE(erroraddr[4]),
.IEF(erroraddr[5]),
.IEG(erroraddr[6]),
.IEH(erroraddr[7]),
.IEI(erroraddr[8]),
.IEJ(erroraddr[9]),
.IEK(erroraddr[10]),
.IEL(erroraddr[11]),
.IEM(erroraddr[12]),
.IEN(erroraddr[13]),
.IEO(erroraddr[14]),
.IEP(erroraddr[15]),
.IFA(erroraddr[16]),
.IFB(erroraddr[17]),
.IFC(erroraddr[18]),
.IFD(erroraddr[19]),
.IFE(erroraddr[20]),
.IFFF(erroraddr[21]),
.IFG(erroraddr[22]),
.IFH(erroraddr[23]),
.IFI(erroraddr[24]),
.IFJ(erroraddr[25]),
.IFK(erroraddr[26]),
.IFL(erroraddr[27]),
.IFM(erroraddr[28]),
.IFN(erroraddr[29]),
.IFO(erroraddr[30]),
.IFP(erroraddr[31]),
.IGA(syndrome[0]),
.IGB(syndrome[1]),
.IGC(syndrome[2]),
.IGD(syndrome[3]),
.IGE(syndrome[4]),
.IGF(syndrome[5]),
.IGG(syndrome[6]),
.IGH(syndrome[7]),
.IHA(fetcharrivaltoeb[0]),
.IHB(fetcharrivaltoeb[1]),
.IHC(fetcharrivaltoeb[2]),
.IIA(singlebiterror),
.IIB(doublebiterror),
.IJA(gowritetoeb),
.IJB(endsequencetoeb),
.IKA(flooptoeb[0]),
.IKB(flooptoeb[1]),
.IKC(flooptoeb[2]),
.IKD(flooptoeb[3]),
.IKE(flooptoeb[4]),
.IKF(flooptoeb[5]),
.IKG(flooptoeb[6]),
.IKH(flooptoeb[7]),
.IKI(flooptoeb[8]),
.IKJ(flooptoeb[9]),
.IKK(flooptoeb[10]),
.IKL(flooptoeb[11]),
.IKM(flooptoeb[12]),
.IKN(flooptoeb[13]),
.IKO(flooptoeb[14]),
.IKP(flooptoeb[15]),
.IKQ(flooptoeb[16]),
.IKR(flooptoeb[17]),
.IKS(flooptoeb[18]),
.IKT(flooptoeb[19]),
.IMA(deadstarteb),
.INA(nxtcpublockref),
.INB(nxtcpup1blockref),
.INC(nxtcpup2blockref),
.IND(refreshenable),
.INE(gatewdfromib),
.IZZ (sysclock),
.OAA(ebdatatb[0]),
.OAB(ebdatatb[1]),
.OAC(ebdatatb[2]),
.OAD(ebdatatb[3]),
.OAE(ebdatatb[4]),
.OAF(ebdatatb[5]),
.OAG(ebdatatb[6]),
.OAH(ebdatatb[7]),
.OAI(ebdatatb[8]),
.OAJ(ebdatatb[9]),
.OAK(ebdatatb[10]),
.OAL(ebdatatb[11]),
.OAM(ebdatatb[12]),
.OAN(ebdatatb[13]),
.OAO(ebdatatb[14]),
.OAP(ebdatatb[15]),
.OBA(ebdatatb[16]),
.OBB(ebdatatb[17]),
.OBC(ebdatatb[18]),
.OBD(ebdatatb[19]),
.OBE(ebdatatb[20]),
.OBF(ebdatatb[21]),
.OBG(ebdatatb[22]),
.OBH(ebdatatb[23]),
.OBI(ebdatatb[24]),
.OBJ(ebdatatb[25]),
.OBK(ebdatatb[26]),
.OBL(ebdatatb[27]),
.OBM(ebdatatb[28]),
.OBN(ebdatatb[29]),
.OBO(ebdatatb[30]),
.OBP(ebdatatb[31]),
.OCA(ebdatatb[32]),
.OCB(ebdatatb[33]),
.OCC(ebdatatb[34]),
.OCD(ebdatatb[35]),
.OCE(ebdatatb[36]),
.OCF(ebdatatb[37]),
.OCG(ebdatatb[38]),
.OCH(ebdatatb[39]),
.OCI(ebdatatb[40]),
.OCJ(ebdatatb[41]),
.OCK(ebdatatb[42]),
.OCL(ebdatatb[43]),
.OCM(ebdatatb[44]),
.OCN(ebdatatb[45]),
.OCO(ebdatatb[46]),
.OCP(ebdatatb[47]),
.ODA(ebdatatb[48]),
.ODB(ebdatatb[49]),
.ODC(ebdatatb[50]),
.ODD(ebdatatb[51]),
.ODE(ebdatatb[52]),
.ODF(ebdatatb[53]),
.ODG(ebdatatb[54]),
.ODH(ebdatatb[55]),
.ODI(ebdatatb[56]),
.ODJ(ebdatatb[57]),
.ODK(ebdatatb[58]),
.ODL(ebdatatb[59]),
.ODM(ebdatatb[60]),
.ODN(ebdatatb[61]),
.ODO(ebdatatb[62]),
.ODP(ebdatatb[63]),
.OEA(ebaddrtotf[0]),
.OEB(ebaddrtotf[1]),
.OEC(ebaddrtotf[2]),
.OED(ebaddrtotf[3]),
.OEE(ebaddrtotf[4]),
.OEF(ebaddrtotf[5]),
.OEG(ebaddrtotf[6]),
.OEH(ebaddrtotf[7]),
.OEI(ebaddrtotf[8]),
.OEJ(ebaddrtotf[9]),
.OEK(ebaddrtotf[10]),
.OEL(ebaddrtotf[11]),
.OEM(ebaddrtotf[12]),
.OEN(ebaddrtotf[13]),
.OEO(ebaddrtotf[14]),
.OEP(ebaddrtotf[15]),
.OFA(ebaddrtotf[16]),
.OFB(ebaddrtotf[17]),
.OFC(ebaddrtotf[18]),
.OFD(ebaddrtotf[19]),
.OFE(ebaddrtotf[20]),
.OFF(ebaddrtotf[21]),
.OFG(ebaddrtotf[22]),
.OFH(ebaddrtotf[23]),
.OFI(ebaddrtotf[24]),
.OFJ(ebaddrtotf[25]),
.OFK(ebaddrtotf[26]),
.OFL(ebaddrtotf[27]),
.OFM(ebaddrtotf[28]),
.OFN(ebaddrtotf[29]),
.OFO(ebaddrtotf[30]),
.OFP(ebaddrtotf[31]),
.OGA(iolentoif[0]),
.OGB(iolentoif[1]),
.OGC(iolentoif[2]),
.OGD(iolentoif[3]),
.OGE(iolentoif[4]),
.OGF(iolentoif[5]),
.OHA(exterreftoif),
.OHB(readmodetoif),
.OHC(blockreftonext),
.OHD(blockreftonextp1),
.OHE(blockreftonextp2),
.OHF(blockreftonextp3),
.OHG(refreshtotf),
.OKA(floopfrmeb[0]),
.OKB(floopfrmeb[1]),
.OKC(floopfrmeb[2]),
.OKD(floopfrmeb[3]),
.OKE(floopfrmeb[4]),
.OKF(floopfrmeb[5]),
.OKG(floopfrmeb[6]),
.OKH(floopfrmeb[7]),
.OKI(floopfrmeb[8]),
.OKJ(floopfrmeb[9]),
.OKK(floopfrmeb[10]),
.OKL(floopfrmeb[11]),
.OKM(floopfrmeb[12]),
.OKN(floopfrmeb[13]),
.OKO(floopfrmeb[14]),
.OKP(floopfrmeb[15]),
.OKQ(floopfrmeb[16]),
.OKR(floopfrmeb[17]),
.OKS(floopfrmeb[18]),
.OKT(floopfrmeb[19]),
.OLA(functiondcdlights[0]),
.OLB(functiondcdlights[1]),
.OLC(functiondcdlights[2]),
.OLD(functiondcdlights[3]),
.OLE(functiondcdlights[4]),
.OLF(functiondcdlights[5]),
.OLG(functiondcdlights[6]),
.OLH(functiondcdlights[7]));


  
fa fa0 (
.IAA(vrtofak[0]),
.IAB(vrtofak[1]),
.IAC(vrtofak[2]),
.IAD(vrtofak[3]),
.IAE(vrtofak[4]),
.IAF(vrtofak[5]),
.IAG(vrtofak[6]),
.IAH(vrtofak[7]),
.IAI(vrtofak[8]),
.IAJ(vrtofak[9]),
.IAK(vrtofak[10]),
.IAL(vrtofak[11]),
.IAM(vrtofak[12]),
.IAN(vrtofak[13]),
.IAO(vrtofak[14]),
.IAP(vrtofak[15]),
.IBA(vrtofak[16]),
.IBB(vrtofak[17]),
.IBC(vrtofak[18]),
.IBD(vrtofak[19]),
.IBE(vrtofak[20]),
.IBF(vrtofak[21]),
.IBG(vrtofak[22]),
.IBH(vrtofak[23]),
.IBI(vrtofak[24]),
.IBJ(vrtofak[25]),
.IBK(vrtofak[26]),
.IBL(vrtofak[27]),
.IBM(vrtofak[28]),
.IBN(vrtofak[29]),
.IBO(vrtofak[30]),
.IBP(vrtofak[31]),
.ICA(vrtofak[32]),
.ICB(vrtofak[33]),
.ICC(vrtofak[34]),
.ICD(vrtofak[35]),
.ICE(vrtofak[36]),
.ICF(vrtofak[37]),
.ICG(vrtofak[38]),
.ICH(vrtofak[39]),
.ICI(vrtofak[40]),
.ICJ(vrtofak[41]),
.ICK(vrtofak[42]),
.ICL(vrtofak[43]),
.ICM(vrtofak[44]),
.ICN(vrtofak[45]),
.ICO(vrtofak[46]),
.ICP(vrtofak[47]),
.IDA(vrtofak[48]),
.IDB(vrtofak[49]),
.IDC(vrtofak[50]),
.IDD(vrtofak[51]),
.IDE(vrtofak[52]),
.IDF(vrtofak[53]),
.IDG(vrtofak[54]),
.IDH(vrtofak[55]),
.IDI(vrtofak[56]),
.IDJ(vrtofak[57]),
.IDK(vrtofak[58]),
.IDL(vrtofak[59]),
.IDM(vrtofak[60]),
.IDN(vrtofak[61]),
.IDO(vrtofak[62]),
.IDP(vrtofak[63]),
.IEA(vrtofaj[0]),
.IEB(vrtofaj[1]),
.IEC(vrtofaj[2]),
.IED(vrtofaj[3]),
.IEE(vrtofaj[4]),
.IEF(vrtofaj[5]),
.IEG(vrtofaj[6]),
.IEH(vrtofaj[7]),
.IEI(vrtofaj[8]),
.IEJ(vrtofaj[9]),
.IEK(vrtofaj[10]),
.IEL(vrtofaj[11]),
.IEM(vrtofaj[12]),
.IEN(vrtofaj[13]),
.IEO(vrtofaj[14]),
.IEP(vrtofaj[15]),
.IFA(vrtofaj[16]),
.IFB(vrtofaj[17]),
.IFC(vrtofaj[18]),
.IFD(vrtofaj[19]),
.IFE(vrtofaj[20]),
.IFFF(vrtofaj[21]),
.IFG(vrtofaj[22]),
.IFH(vrtofaj[23]),
.IFI(vrtofaj[24]),
.IFJ(vrtofaj[25]),
.IFK(vrtofaj[26]),
.IFL(vrtofaj[27]),
.IFM(vrtofaj[28]),
.IFN(vrtofaj[29]),
.IFO(vrtofaj[30]),
.IFP(vrtofaj[31]),
.IGA(vrtofaj[32]),
.IGB(vrtofaj[33]),
.IGC(vrtofaj[34]),
.IGD(vrtofaj[35]),
.IGE(vrtofaj[36]),
.IGF(vrtofaj[37]),
.IGG(vrtofaj[38]),
.IGH(vrtofaj[39]),
.IGI(vrtofaj[40]),
.IGJ(vrtofaj[41]),
.IGK(vrtofaj[42]),
.IGL(vrtofaj[43]),
.IGM(vrtofaj[44]),
.IGN(vrtofaj[45]),
.IGO(vrtofaj[46]),
.IGP(vrtofaj[47]),
.IHA(vrtofaj[48]),
.IHB(vrtofaj[49]),
.IHC(vrtofaj[50]),
.IHD(vrtofaj[51]),
.IHE(vrtofaj[52]),
.IHF(vrtofaj[53]),
.IHG(vrtofaj[54]),
.IHH(vrtofaj[55]),
.IHI(vrtofaj[56]),
.IHJ(vrtofaj[57]),
.IHK(vrtofaj[58]),
.IHL(vrtofaj[59]),
.IHM(vrtofaj[60]),
.IHN(vrtofaj[61]),
.IHO(vrtofaj[62]),
.IHP(vrtofaj[63]),
.IJA(jafacnt[0]),
.IJB(jafacnt[1]),
.IJC(jafacnt[2]),
.IJD(jafacnt[3]),
.IJE(jafacnt[4]),
.IKA(vectorlencntl),
.ILA(enablefarangeerr),
.IZZ (sysclock),
.OAA(shftcoef[0]),
.OAB(shftcoef[1]),
.OAC(shftcoef[2]),
.OAD(shftcoef[3]),
.OAE(shftcoef[4]),
.OAF(shftcoef[5]),
.OAG(shftcoef[6]),
.OAH(shftcoef[7]),
.OAI(shftcoef[8]),
.OAJ(shftcoef[9]),
.OAK(shftcoef[10]),
.OAL(shftcoef[11]),
.OAM(shftcoef[12]),
.OAN(shftcoef[13]),
.OAO(shftcoef[14]),
.OAP(shftcoef[15]),
.OAR(shftcoeflo),
.OBA(shftcoef[16]),
.OBB(shftcoef[17]),
.OBC(shftcoef[18]),
.OBD(shftcoef[19]),
.OBE(shftcoef[20]),
.OBF(shftcoef[21]),
.OBG(shftcoef[22]),
.OBH(shftcoef[23]),
.OBI(shftcoef[24]),
.OBJ(shftcoef[25]),
.OBK(shftcoef[26]),
.OBL(shftcoef[27]),
.OBM(shftcoef[28]),
.OBN(shftcoef[29]),
.OBO(shftcoef[30]),
.OBP(shftcoef[31]),
.OCA(shftcoef[32]),
.OCB(shftcoef[33]),
.OCC(shftcoef[34]),
.OCD(shftcoef[35]),
.OCE(shftcoef[36]),
.OCF(shftcoef[37]),
.OCG(shftcoef[38]),
.OCH(shftcoef[39]),
.OCI(shftcoef[40]),
.OCJ(shftcoef[41]),
.OCK(shftcoef[42]),
.OCL(shftcoef[43]),
.OCM(shftcoef[44]),
.OCN(shftcoef[45]),
.OCO(shftcoef[46]),
.OCP(shftcoef[47]),
.ODA(coeftofb[0]),
.ODB(coeftofb[1]),
.ODC(coeftofb[2]),
.ODD(coeftofb[3]),
.ODE(coeftofb[4]),
.ODF(coeftofb[5]),
.ODG(coeftofb[6]),
.ODH(coeftofb[7]),
.ODI(coeftofb[8]),
.ODJ(coeftofb[9]),
.ODK(coeftofb[10]),
.ODL(coeftofb[11]),
.ODM(coeftofb[12]),
.ODN(coeftofb[13]),
.ODO(coeftofb[14]),
.ODP(coeftofb[15]),
.OEA(coeftofb[16]),
.OEB(coeftofb[17]),
.OEC(coeftofb[18]),
.OED(coeftofb[19]),
.OEE(coeftofb[20]),
.OEF(coeftofb[21]),
.OEG(coeftofb[22]),
.OEH(coeftofb[23]),
.OEI(coeftofb[24]),
.OEJ(coeftofb[25]),
.OEK(coeftofb[26]),
.OEL(coeftofb[27]),
.OEM(coeftofb[28]),
.OEN(coeftofb[29]),
.OEO(coeftofb[30]),
.OEP(coeftofb[31]),
.OFA(coeftofb[32]),
.OFB(coeftofb[33]),
.OFC(coeftofb[34]),
.OFD(coeftofb[35]),
.OFE(coeftofb[36]),
.OFF(coeftofb[37]),
.OFG(coeftofb[38]),
.OFH(coeftofb[39]),
.OFI(coeftofb[40]),
.OFJ(coeftofb[41]),
.OFK(coeftofb[42]),
.OFL(coeftofb[43]),
.OFM(coeftofb[44]),
.OFN(coeftofb[45]),
.OFO(coeftofb[46]),
.OFP(coeftofb[47]),
.OGA(exptofc[0]),
.OGB(exptofc[1]),
.OGC(exptofc[2]),
.OGD(exptofc[3]),
.OGE(exptofc[4]),
.OGF(exptofc[5]),
.OGG(exptofc[6]),
.OGH(exptofc[7]),
.OGI(exptofc[8]),
.OGJ(exptofc[9]),
.OGK(exptofc[10]),
.OGL(exptofc[11]),
.OGM(exptofc[12]),
.OGN(exptofc[13]),
.OGO(exptofc[14]),
.OGP(exptofc[15]),
.OHA(fbsubtractmode),
.OIA(constoverflfc),
.OJA(fbgoadd),
.OJB(gocons122174),
.OJC(gocons123175),
.OKA(enablerangerrfc));

  
fb fb0 (
.IAA(shftcoef[0]),
.IAB(shftcoef[1]),
.IAC(shftcoef[2]),
.IAD(shftcoef[3]),
.IAE(shftcoef[4]),
.IAF(shftcoef[5]),
.IAG(shftcoef[6]),
.IAH(shftcoef[7]),
.IAI(shftcoef[8]),
.IAJ(shftcoef[9]),
.IAK(shftcoef[10]),
.IAL(shftcoef[11]),
.IAM(shftcoef[12]),
.IAN(shftcoef[13]),
.IAO(shftcoef[14]),
.IAP(shftcoef[15]),
.IAR(shftcoeflo),
.IBA(shftcoef[16]),
.IBB(shftcoef[17]),
.IBC(shftcoef[18]),
.IBD(shftcoef[19]),
.IBE(shftcoef[20]),
.IBF(shftcoef[21]),
.IBG(shftcoef[22]),
.IBH(shftcoef[23]),
.IBI(shftcoef[24]),
.IBJ(shftcoef[25]),
.IBK(shftcoef[26]),
.IBL(shftcoef[27]),
.IBM(shftcoef[28]),
.IBN(shftcoef[29]),
.IBO(shftcoef[30]),
.IBP(shftcoef[31]),
.ICA(shftcoef[32]),
.ICB(shftcoef[33]),
.ICC(shftcoef[34]),
.ICD(shftcoef[35]),
.ICE(shftcoef[36]),
.ICF(shftcoef[37]),
.ICG(shftcoef[38]),
.ICH(shftcoef[39]),
.ICI(shftcoef[40]),
.ICJ(shftcoef[41]),
.ICK(shftcoef[42]),
.ICL(shftcoef[43]),
.ICM(shftcoef[44]),
.ICN(shftcoef[45]),
.ICO(shftcoef[46]),
.ICP(shftcoef[47]),
.IDA(coeftofb[0]),
.IDB(coeftofb[1]),
.IDC(coeftofb[2]),
.IDD(coeftofb[3]),
.IDE(coeftofb[4]),
.IDF(coeftofb[5]),
.IDG(coeftofb[6]),
.IDH(coeftofb[7]),
.IDI(coeftofb[8]),
.IDJ(coeftofb[9]),
.IDK(coeftofb[10]),
.IDL(coeftofb[11]),
.IDM(coeftofb[12]),
.IDN(coeftofb[13]),
.IDO(coeftofb[14]),
.IDP(coeftofb[15]),
.IEA(coeftofb[16]),
.IEB(coeftofb[17]),
.IEC(coeftofb[18]),
.IED(coeftofb[19]),
.IEE(coeftofb[20]),
.IEF(coeftofb[21]),
.IEG(coeftofb[22]),
.IEH(coeftofb[23]),
.IEI(coeftofb[24]),
.IEJ(coeftofb[25]),
.IEK(coeftofb[26]),
.IEL(coeftofb[27]),
.IEM(coeftofb[28]),
.IEN(coeftofb[29]),
.IEO(coeftofb[30]),
.IEP(coeftofb[31]),
.IFA(coeftofb[32]),
.IFB(coeftofb[33]),
.IFC(coeftofb[34]),
.IFD(coeftofb[35]),
.IFE(coeftofb[36]),
.IFFF(coeftofb[37]),
.IFG(coeftofb[38]),
.IFH(coeftofb[39]),
.IFI(coeftofb[40]),
.IFJ(coeftofb[41]),
.IFK(coeftofb[42]),
.IFL(coeftofb[43]),
.IFM(coeftofb[44]),
.IFN(coeftofb[45]),
.IFO(coeftofb[46]),
.IFP(coeftofb[47]),
.IJA(fbsubtractmode),
.IJB(fbgoadd),
.IZZ (sysclock),
.OAA(signtofc[0]),
.OAB(signtofc[1]),
.OAC(signtofc[2]),
.OAD(signtofc[3]),
.OAE(signtofc[4]),
.OAF(signtofc[5]),
.OAG(signtofc[6]),
.OAH(signtofc[7]),
.OAI(signtofc[8]),
.OAJ(signtofc[9]),
.OAK(signtofc[10]),
.OAL(signtofc[11]),
.OAM(signtofc[12]),
.OAN(signtofc[13]),
.OAO(signtofc[14]),
.OAP(signtofc[15]),
.OBA(signtofc[16]),
.OBB(signtofc[17]),
.OBC(signtofc[18]),
.OBD(signtofc[19]),
.OBE(signtofc[20]),
.OBF(signtofc[21]),
.OBG(signtofc[22]),
.OBH(signtofc[23]),
.OBI(signtofc[24]),
.OBJ(signtofc[25]),
.OBK(signtofc[26]),
.OBL(signtofc[27]),
.OBM(signtofc[28]),
.OBN(signtofc[29]),
.OBO(signtofc[30]),
.OBP(signtofc[31]),
.OCA(signtofc[32]),
.OCB(signtofc[33]),
.OCC(signtofc[34]),
.OCD(signtofc[35]),
.OCE(signtofc[36]),
.OCF(signtofc[37]),
.OCG(signtofc[38]),
.OCH(signtofc[39]),
.OCI(signtofc[40]),
.OCJ(signtofc[41]),
.OCK(signtofc[42]),
.OCL(signtofc[43]),
.OCM(signtofc[44]),
.OCN(signtofc[45]),
.OCO(signtofc[46]),
.OCP(signtofc[47]),
.ODA( normalizecnt[5]),
.ODB( normalizecnt[4]),
.ODC( normalizecnt[3]),
.ODD( normalizecnt[2]),
.ODE( normalizecnt12),
.OEA(sect0tofc[0]),
.OEB(sect0tofc[1]),
.OFA(sect1tofc[0]),
.OFB(sect1tofc[1]),
.OGA(sect2tofc[0]),
.OGB(sect2tofc[1]),
.OHA(togglesign),
.OHB(shifteqminus1),
.OIA(cunderflowtofc),
.OJA(goaddtofc),
.OJB(unlikesigns));

  
fc fc0 (
.IAA(signtofc[0]),
.IAB(signtofc[1]),
.IAC(signtofc[2]),
.IAD(signtofc[3]),
.IAE(signtofc[4]),
.IAF(signtofc[5]),
.IAG(signtofc[6]),
.IAH(signtofc[7]),
.IAI(signtofc[8]),
.IAJ(signtofc[9]),
.IAK(signtofc[10]),
.IAL(signtofc[11]),
.IAM(signtofc[12]),
.IAN(signtofc[13]),
.IAO(signtofc[14]),
.IAP(signtofc[15]),
.IBA(signtofc[16]),
.IBB(signtofc[17]),
.IBC(signtofc[18]),
.IBD(signtofc[19]),
.IBE(signtofc[20]),
.IBF(signtofc[21]),
.IBG(signtofc[22]),
.IBH(signtofc[23]),
.IBI(signtofc[24]),
.IBJ(signtofc[25]),
.IBK(signtofc[26]),
.IBL(signtofc[27]),
.IBM(signtofc[28]),
.IBN(signtofc[29]),
.IBO(signtofc[30]),
.IBP(signtofc[31]),
.ICA(signtofc[32]),
.ICB(signtofc[33]),
.ICC(signtofc[34]),
.ICD(signtofc[35]),
.ICE(signtofc[36]),
.ICF(signtofc[37]),
.ICG(signtofc[38]),
.ICH(signtofc[39]),
.ICI(signtofc[40]),
.ICJ(signtofc[41]),
.ICK(signtofc[42]),
.ICL(signtofc[43]),
.ICM(signtofc[44]),
.ICN(signtofc[45]),
.ICO(signtofc[46]),
.ICP(signtofc[47]),
.IDA(exptofc[0]),
.IDB(exptofc[1]),
.IDC(exptofc[2]),
.IDD(exptofc[3]),
.IDE(exptofc[4]),
.IDF(exptofc[5]),
.IDG(exptofc[6]),
.IDH(exptofc[7]),
.IDI(exptofc[8]),
.IDJ(exptofc[9]),
.IDK(exptofc[10]),
.IDL(exptofc[11]),
.IDM(exptofc[12]),
.IDN(exptofc[13]),
.IDO(exptofc[14]),
.IDP(exptofc[15]),
.IEA(sect2tofc[0]),
.IEB(sect2tofc[1]),
.IEC(sect1tofc[0]),
.IED(sect1tofc[1]),
.IEE(sect0tofc[0]),
.IEF(sect0tofc[1]),
.IEG( normalizecnt[2]),
.IEH( normalizecnt[3]),
.IEI( normalizecnt[4]),
.IEJ( normalizecnt[5]),
.IEK( normalizecnt12),
.IHA(togglesign),
.IHB(shifteqminus1),
.IIA(cunderflowtofc),
.IIB(constoverflfc),
.IJA(goaddtofc),
.IJB(gocons122174),
.IJC(gocons123175),
.IJD(unlikesigns),
.IKA(enablerangerrfc),
.IZZ (sysclock),
.OAA(fctovr[0]),
.OAB(fctovr[1]),
.OAC(fctovr[2]),
.OAD(fctovr[3]),
.OAE(fctovr[4]),
.OAF(fctovr[5]),
.OAG(fctovr[6]),
.OAH(fctovr[7]),
.OAI(fctovr[8]),
.OAJ(fctovr[9]),
.OAK(fctovr[10]),
.OAL(fctovr[11]),
.OAM(fctovr[12]),
.OAN(fctovr[13]),
.OAO(fctovr[14]),
.OAP(fctovr[15]),
.OBA(fctovr[16]),
.OBB(fctovr[17]),
.OBC(fctovr[18]),
.OBD(fctovr[19]),
.OBE(fctovr[20]),
.OBF(fctovr[21]),
.OBG(fctovr[22]),
.OBH(fctovr[23]),
.OBI(fctovr[24]),
.OBJ(fctovr[25]),
.OBK(fctovr[26]),
.OBL(fctovr[27]),
.OBM(fctovr[28]),
.OBN(fctovr[29]),
.OBO(fctovr[30]),
.OBP(fctovr[31]),
.OCA(fctovr[32]),
.OCB(fctovr[33]),
.OCC(fctovr[34]),
.OCD(fctovr[35]),
.OCE(fctovr[36]),
.OCF(fctovr[37]),
.OCG(fctovr[38]),
.OCH(fctovr[39]),
.OCI(fctovr[40]),
.OCJ(fctovr[41]),
.OCK(fctovr[42]),
.OCL(fctovr[43]),
.OCM(fctovr[44]),
.OCN(fctovr[45]),
.OCO(fctovr[46]),
.OCP(fctovr[47]),
.ODA(fctovr[48]),
.ODB(fctovr[49]),
.ODC(fctovr[50]),
.ODD(fctovr[51]),
.ODE(fctovr[52]),
.ODF(fctovr[53]),
.ODG(fctovr[54]),
.ODH(fctovr[55]),
.ODI(fctovr[56]),
.ODJ(fctovr[57]),
.ODK(fctovr[58]),
.ODL(fctovr[59]),
.ODM(fctovr[60]),
.ODN(fctovr[61]),
.ODO(fctovr[62]),
.ODP(fctovr[63]),
.OEA(fprangeerrfc));
  
ga ga0 (
.IAA(scdatatoga[0]),
.IAB(scdatatoga[1]),
.IAC(scdatatoga[2]),
.IAD(scdatatoga[3]),
.IAE(scdatatoga[4]),
.IAF(scdatatoga[5]),
.IAG(scdatatoga[6]),
.IAH(scdatatoga[7]),
.IAI(scdatatoga[8]),
.IAJ(scdatatoga[9]),
.IAK(scdatatoga[10]),
.IAL(scdatatoga[11]),
.IAM(scdatatoga[12]),
.IAN(scdatatoga[13]),
.IAO(scdatatoga[14]),
.IAP(scdatatoga[15]),
.IBA(scdatatoga[16]),
.IBB(scdatatoga[17]),
.IBC(scdatatoga[18]),
.IBD(scdatatoga[19]),
.IBE(scdatatoga[20]),
.IBF(scdatatoga[21]),
.IBG(scdatatoga[22]),
.IBH(scdatatoga[23]),
.IBI(scdatatoga[24]),
.IBJ(scdatatoga[25]),
.IBK(scdatatoga[26]),
.IBL(scdatatoga[27]),
.IBM(scdatatoga[28]),
.IBN(scdatatoga[29]),
.IBO(scdatatoga[30]),
.IBP(scdatatoga[31]),
.ICA(scdatatoga[32]),
.ICB(scdatatoga[33]),
.ICC(scdatatoga[34]),
.ICD(scdatatoga[35]),
.ICE(scdatatoga[36]),
.ICF(scdatatoga[37]),
.ICG(scdatatoga[38]),
.ICH(scdatatoga[39]),
.ICI(scdatatoga[40]),
.ICJ(scdatatoga[41]),
.ICK(scdatatoga[42]),
.ICL(scdatatoga[43]),
.ICM(scdatatoga[44]),
.ICN(scdatatoga[45]),
.ICO(scdatatoga[46]),
.ICP(scdatatoga[47]),
.IDA(scdatatoga[48]),
.IDB(scdatatoga[49]),
.IDC(scdatatoga[50]),
.IDD(scdatatoga[51]),
.IDE(scdatatoga[52]),
.IDF(scdatatoga[53]),
.IDG(scdatatoga[54]),
.IDH(scdatatoga[55]),
.IDI(scdatatoga[56]),
.IDJ(scdatatoga[57]),
.IDK(scdatatoga[58]),
.IDL(scdatatoga[59]),
.IDM(scdatatoga[60]),
.IDN(scdatatoga[61]),
.IDO(scdatatoga[62]),
.IDP(scdatatoga[63]),
.IGA(jagacnt[0]),
.IPB(jagacnt[1]),
.IPC(jagacnt[2]),
.IPD(jagacnt[3]),
.IZZ (sysclock),
.OAA(gatovr[0]),
.OAB(gatovr[1]),
.OAC(gatovr[2]),
.OAD(gatovr[3]),
.OAE(gatovr[4]),
.OAF(gatovr[5]),
.OAG(gatovr[6]),
.OAH(gatovr[7]),
.OAI(gatovr[8]),
.OAJ(gatovr[9]),
.OAK(gatovr[10]),
.OAL(gatovr[11]),
.OAM(gatovr[12]),
.OAN(gatovr[13]),
.OAO(gatovr[14]),
.OAP(gatovr[15]),
.OBA(gatovr[16]),
.OBB(gatovr[17]),
.OBC(gatovr[18]),
.OBD(gatovr[19]),
.OBE(gatovr[20]),
.OBF(gatovr[21]),
.OBG(gatovr[22]),
.OBH(gatovr[23]),
.OBI(gatovr[24]),
.OBJ(gatovr[25]),
.OBK(gatovr[26]),
.OBL(gatovr[27]),
.OBM(gatovr[28]),
.OBN(gatovr[29]),
.OBO(gatovr[30]),
.OBP(gatovr[31]),
.OCA(gatovr[32]),
.OCB(gatovr[33]),
.OCC(gatovr[34]),
.OCD(gatovr[35]),
.OCE(gatovr[36]),
.OCF(gatovr[37]),
.OCG(gatovr[38]),
.OCH(gatovr[39]),
.OCI(gatovr[40]),
.OCJ(gatovr[41]),
.OCK(gatovr[42]),
.OCL(gatovr[43]),
.OCM(gatovr[44]),
.OCN(gatovr[45]),
.OCO(gatovr[46]),
.OCP(gatovr[47]),
.ODA(gatovr[48]),
.ODB(gatovr[49]),
.ODC(gatovr[50]),
.ODD(gatovr[51]),
.ODE(gatovr[52]),
.ODF(gatovr[53]),
.ODG(gatovr[54]),
.ODH(gatovr[55]),
.ODI(gatovr[56]),
.ODJ(gatovr[57]),
.ODK(gatovr[58]),
.ODL(gatovr[59]),
.ODM(gatovr[60]),
.ODN(gatovr[61]),
.ODO(gatovr[62]),
.ODP(gatovr[63]));


gb gb0 (
.IAA(shftcnt[0]),
.IAB(shftcnt[1]),
.IAC(shftcnt[2]),
.IAD(shftcnt[3]),
.IAE(shftcnt[4]),
.IAF(shftcnt[5]),
.IAG(shftcnt[6]),
.IAH(shftovfl[0]),
.IAI(shftovfl[1]),
.IAJ(shftovfl[2]),
.IIA(shdatatogb[0]),
.IIB(shdatatogb[1]),
.IIC(shdatatogb[2]),
.IID(shdatatogb[3]),
.IIE(shdatatogb[4]),
.IIF(shdatatogb[5]),
.IIG(shdatatogb[6]),
.IIH(shdatatogb[7]),
.III(shdatatogb[8]),
.IIJ(shdatatogb[9]),
.IIK(shdatatogb[10]),
.IIL(shdatatogb[11]),
.IIM(shdatatogb[12]),
.IIN(shdatatogb[13]),
.IIO(shdatatogb[14]),
.IIP(shdatatogb[15]),
.IJA(shdatatogb[16]),
.IJB(shdatatogb[17]),
.IJC(shdatatogb[18]),
.IJD(shdatatogb[19]),
.IJE(shdatatogb[20]),
.IJF(shdatatogb[21]),
.IJG(shdatatogb[22]),
.IJH(shdatatogb[23]),
.IJI(shdatatogb[24]),
.IJJ(shdatatogb[25]),
.IJK(shdatatogb[26]),
.IJL(shdatatogb[27]),
.IJM(shdatatogb[28]),
.IJN(shdatatogb[29]),
.IJO(shdatatogb[30]),
.IJP(shdatatogb[31]),
.IKA(shdatatogb[32]),
.IKB(shdatatogb[33]),
.IKC(shdatatogb[34]),
.IKD(shdatatogb[35]),
.IKE(shdatatogb[36]),
.IKF(shdatatogb[37]),
.IKG(shdatatogb[38]),
.IKH(shdatatogb[39]),
.IKI(shdatatogb[40]),
.IKJ(shdatatogb[41]),
.IKK(shdatatogb[42]),
.IKL(shdatatogb[43]),
.IKM(shdatatogb[44]),
.IKN(shdatatogb[45]),
.IKO(shdatatogb[46]),
.IKP(shdatatogb[47]),
.ILA(shdatatogb[48]),
.ILB(shdatatogb[49]),
.ILC(shdatatogb[50]),
.ILD(shdatatogb[51]),
.ILE(shdatatogb[52]),
.ILF(shdatatogb[53]),
.ILG(shdatatogb[54]),
.ILH(shdatatogb[55]),
.ILI(shdatatogb[56]),
.ILJ(shdatatogb[57]),
.ILK(shdatatogb[58]),
.ILL(shdatatogb[59]),
.ILM(shdatatogb[60]),
.ILN(shdatatogb[61]),
.ILO(shdatatogb[62]),
.ILP(shdatatogb[63]),
.INA(jagbcnt[0]),
.INB(jagbcnt[1]),
.INC(jagbcnt[2]),
.IND(jagbcnt[3]),
.INE(jagbcnt[4]),
.INF(jagbcnt[5]),
.IOA(shftcontogb[0]),
.IOB(shftcontogb[1]),
.IOC(shftcontogb[2]),
.IRA(akshtogb[0]), 
.IRB(akshtogb[1]),
.IRC(akshtogb[2]),
.IRD(akshtogb[3]),
.IRE(akshtogb[4]),
.IRF(akshtogb[5]),
.IRG(akshtogb[6]),
.IRH(akshtogb[7]),
.IRI(akshtogb[8]),
.IRJ(akshtogb[9]),
.IRK(akshtogb[10]),
.IRL(akshtogb[11]),
.IRM(akshtogb[12]),
.IRN(akshtogb[13]),
.IRO(akshtogb[14]),
.IRP(akshtogb[15]),
.IZZ (sysclock),
.OAA(gbtovr[0]),
.OAB(gbtovr[1]),
.OAC(gbtovr[2]),
.OAD(gbtovr[3]),
.OAE(gbtovr[4]),
.OAF(gbtovr[5]),
.OAG(gbtovr[6]),
.OAH(gbtovr[7]),
.OBA(gbtovr[8]),
.OBB(gbtovr[9]),
.OBC(gbtovr[10]),
.OBD(gbtovr[11]),
.OBE(gbtovr[12]),
.OBF(gbtovr[13]),
.OBG(gbtovr[14]),
.OBH(gbtovr[15]),
.OCA(gbtovr[16]),
.OCB(gbtovr[17]),
.OCC(gbtovr[18]),
.OCD(gbtovr[19]),
.OCE(gbtovr[20]),
.OCF(gbtovr[21]),
.OCG(gbtovr[22]),
.OCH(gbtovr[23]),
.ODA(gbtovr[24]),
.ODB(gbtovr[25]),
.ODC(gbtovr[26]),
.ODD(gbtovr[27]),
.ODE(gbtovr[28]),
.ODF(gbtovr[29]),
.ODG(gbtovr[30]),
.ODH(gbtovr[31]),
.OEA(gbtovr[32]),
.OEB(gbtovr[33]),
.OEC(gbtovr[34]),
.OED(gbtovr[35]),
.OEE(gbtovr[36]),
.OEF(gbtovr[37]),
.OEG(gbtovr[38]),
.OEH(gbtovr[39]),
.OFA(gbtovr[40]),
.OFB(gbtovr[41]),
.OFC(gbtovr[42]),
.OFD(gbtovr[43]),
.OFE(gbtovr[44]),
.OFF(gbtovr[45]),
.OFG(gbtovr[46]),
.OFH(gbtovr[47]),
.OGA(gbtovr[48]),
.OGB(gbtovr[49]),
.OGC(gbtovr[50]),
.OGD(gbtovr[51]),
.OGE(gbtovr[52]),
.OGF(gbtovr[53]),
.OGG(gbtovr[54]),
.OGH(gbtovr[55]),
.OHA(gbtovr[56]),
.OHB(gbtovr[57]),
.OHC(gbtovr[58]),
.OHD(gbtovr[59]),
.OHE(gbtovr[60]),
.OHF(gbtovr[61]),
.OHG(gbtovr[62]),
.OHH(gbtovr[63]),
.OKA(shtambtovb[0]),
.OKB(shtambtovb[1]),
.OKC(shtambtovb[2]),
.OKD(shtambtovb[3]),
.OKE(shtambtovb[4]),
.OKF(shtambtovb[5]),
.OKG(shtambtovb[6]),
.OKH(shtovflvb),
.ORA(akshtovr[0]),
.ORB(akshtovr[1]),
.ORC(akshtovr[2]),
.ORD(akshtovr[3]),
.ORE(akshtovr[4]),
.ORF(akshtovr[5]),
.ORG(akshtovr[6]),
.ORH(akshtovr[7]),
.ORI(akshtovr[8]),
.ORJ(akshtovr[9]),
.ORK(akshtovr[10]),
.ORL(akshtovr[11]),
.ORM(akshtovr[12]),
.ORN(akshtovr[13]),
.ORO(akshtovr[14]),
.ORP(akshtovr[15]));

ie ie1 ( 
.IAA(commemtoie[0]),
.IAB(commemtoie[1]),
.IAC(commemtoie[2]),
.IAD(commemtoie[3]),
.IAE(commemtoie[4]),
.IAF(commemtoie[5]),
.IAG(commemtoie[6]),
.IAH(commemtoie[7]),
.IAI(commemtoie[8]),
.IAJ(commemtoie[9]),
.IAK(commemtoie[10]),
.IAL(commemtoie[11]),
.IAM(commemtoie[12]),
.IAN(commemtoie[13]),
.IAO(commemtoie[14]),
.IAP(commemtoie[15]),
.IBA(commemtoie[16]),
.IBB(commemtoie[17]),
.IBC(commemtoie[18]),
.IBD(commemtoie[19]),
.IBE(commemtoie[20]),
.IBF(commemtoie[21]),
.IBG(commemtoie[22]),
.IBH(commemtoie[23]),
.IBI(commemtoie[24]),
.IBJ(commemtoie[25]),
.IBK(commemtoie[26]),
.IBL(commemtoie[27]),
.IBM(commemtoie[28]),
.IBN(commemtoie[29]),
.IBO(commemtoie[30]),
.IBP(commemtoie[31]),
.ICA(commemtoie[32]),
.ICB(commemtoie[33]),
.ICC(commemtoie[34]),
.ICD(commemtoie[35]),
.ICE(commemtoie[36]),
.ICF(commemtoie[37]),
.ICG(commemtoie[38]),
.ICH(commemtoie[39]),
.ICI(commemtoie[40]),
.ICJ(commemtoie[41]),
.ICK(commemtoie[42]),
.ICL(commemtoie[43]),
.ICM(commemtoie[44]),
.ICN(commemtoie[45]),
.ICO(commemtoie[46]),
.ICP(commemtoie[47]),
.IDA(commemtoie[48]),
.IDB(commemtoie[49]),
.IDC(commemtoie[50]),
.IDD(commemtoie[51]),
.IDE(commemtoie[52]),
.IDF(commemtoie[53]),
.IDG(commemtoie[54]),
.IDH(commemtoie[55]),
.IDI(commemtoie[56]),
.IDJ(commemtoie[57]),
.IDK(commemtoie[58]),
.IDL(commemtoie[59]),
.IDM(commemtoie[60]),
.IDN(commemtoie[61]),
.IDO(commemtoie[62]),
.IDP(commemtoie[63]),
.IEA(),
.IEB(),
.IEC(),
.IED(),
.IEE(),
.IEF(),
.IEG(),
.IEH(),
.IEI(),
.IEJ(),
.IFA(),
.IFB(),
.IFC(),
.IFD(),
.IFE(),
.IGA(bankarivfromtf[0]),
.IGB(bankarivfromtf[1]),
.IGC(bankarivfromtf[2]),
.IHA(stkbnd[0]),
.IHB(stkbnd[1]),
.IJA(barreltesttoie),
.IJB(branchpreambletoie),
.IJD(branchintoie),
.IJE(branchouttoie),
.IJF(branchfallthrutoie),
.IJG(clearreadadr1),
.IZZ (sysclock),
.OAA(ibufftoja[0]),
.OAB(ibufftoja[1]),
.OAC(ibufftoja[2]),
.OAD(ibufftoja[3]),
.OAE(ibufftoja[4]),
.OAF(ibufftoja[5]),
.OAG(ibufftoja[6]),
.OAH(ibufftoja[7]),
.OAI(ibufftoja[8]),
.OAJ(ibufftoja[9]),
.OAK(ibufftoja[10]),
.OAL(ibufftoja[11]),
.OAM(ibufftoja[12]),
.OAN(ibufftoja[13]),
.OAO(ibufftoja[14]),
.OAP(ibufftoja[15]),
.OBA(ibufftoja[16]),
.OBB(ibufftoja[17]),
.OBC(ibufftoja[18]),
.OBD(ibufftoja[19]),
.OBE(ibufftoja[20]),
.OBF(ibufftoja[21]),
.OBG(ibufftoja[22]),
.OBH(ibufftoja[23]),
.OBI(ibufftoja[24]),
.OBJ(ibufftoja[25]),
.OBK(ibufftoja[26]),
.OBL(ibufftoja[27]),
.OBM(ibufftoja[28]),
.OBN(ibufftoja[29]),
.OBO(ibufftoja[30]),
.OBP(ibufftoja[31]),
.OCA(ibufftoja[32]),
.OCB(ibufftoja[33]),
.OCC(ibufftoja[34]),
.OCD(ibufftoja[35]),
.OCE(ibufftoja[36]),
.OCF(ibufftoja[37]),
.OCG(ibufftoja[38]),
.OCH(ibufftoja[39]),
.OCI(ibufftoja[40]),
.OCJ(ibufftoja[41]),
.OCK(ibufftoja[42]),
.OCL(ibufftoja[43]),
.OCM(ibufftoja[44]),
.OCN(ibufftoja[45]),
.OCO(ibufftoja[46]),
.OCP(ibufftoja[47]),
.ODA(ibufftoja[48]),
.ODB(ibufftoja[49]),
.ODC(ibufftoja[50]),
.ODD(ibufftoja[51]),
.ODE(ibufftoja[52]),
.ODF(ibufftoja[53]),
.ODG(ibufftoja[54]),
.ODH(ibufftoja[55]),
.ODI(ibufftoja[56]),
.ODJ(ibufftoja[57]),
.ODK(ibufftoja[58]),
.ODL(ibufftoja[59]),
.ODM(ibufftoja[60]),
.ODN(ibufftoja[61]),
.ODO(ibufftoja[62]),
.ODP(ibufftoja[63]),
.OEA(commemtoeb[0]),
.OEB(commemtoeb[1]),
.OEC(commemtoeb[2]),
.OED(commemtoeb[3]),
.OEE(commemtoeb[4]),
.OEF(commemtoeb[5]),
.OEG(commemtoeb[6]),
.OEH(commemtoeb[7]),
.OEI(commemtoeb[8]),
.OEJ(commemtoeb[9]),
.OEK(commemtoeb[10]),
.OEL(commemtoeb[11]),
.OEM(commemtoeb[12]),
.OEN(commemtoeb[13]),
.OEO(commemtoeb[14]),
.OEP(commemtoeb[15]),
.OFA(commemtoeb[16]),
.OFB(commemtoeb[17]),
.OFC(commemtoeb[18]),
.OFD(commemtoeb[19]),
.OFE(commemtoeb[20]),
.OFF(commemtoeb[21]),
.OFG(commemtoeb[22]),
.OFH(commemtoeb[23]),
.OFI(commemtoeb[24]),
.OFJ(commemtoeb[25]),
.OFK(commemtoeb[26]),
.OFL(commemtoeb[27]),
.OFM(commemtoeb[28]),
.OFN(commemtoeb[29]),
.OFO(commemtoeb[30]),
.OFP(commemtoeb[31]),
.OGA(commemtoeb[32]),
.OGB(commemtoeb[33]),
.OGC(commemtoeb[34]),
.OGD(commemtoeb[35]),
.OGE(commemtoeb[36]),
.OGF(commemtoeb[37]),
.OGG(commemtoeb[38]),
.OGH(commemtoeb[39]),
.OGI(commemtoeb[40]),
.OGJ(commemtoeb[41]),
.OGK(commemtoeb[42]),
.OGL(commemtoeb[43]),
.OGM(commemtoeb[44]),
.OGN(commemtoeb[45]),
.OGO(commemtoeb[46]),
.OGP(commemtoeb[47]),
.OHA(commemtoeb[48]),
.OHB(commemtoeb[49]),
.OHC(commemtoeb[50]),
.OHD(commemtoeb[51]),
.OHE(commemtoeb[52]),
.OHF(commemtoeb[53]),
.OHG(commemtoeb[54]),
.OHH(commemtoeb[55]),
.OHI(commemtoeb[56]),
.OHJ(commemtoeb[57]),
.OHK(commemtoeb[58]),
.OHL(commemtoeb[59]),
.OHM(commemtoeb[60]),
.OHN(commemtoeb[61]),
.OHO(commemtoeb[62]),
.OHP(commemtoeb[63]),
.OJA(datareadyja),
.OJB(boundflagtotf),
.OJD(fetchcmletetoif),
.OJF(boundaryflagtoif),
.OKA(ieindlights[0]),
.OKB(ieindlights[1]),
.OKC(ieindlights[2]),
.OKG(ieindlights[6]),
.OKH(ieindlights[7]),
.OKI(ieindlights[8]),
.OKJ(ieindlights[9]),
.OKK(ieindlights[10]),
.OKL(ieindlights[11]),
.OKM(ieindlights[12]),
.OKN(ieindlights[13]),
.OKO(ieindlights[14]),
.OKP(ieindlights[15]),
.OKQ(ieindlights[16]),
.OKR(ieindlights[17]),
.OKS(ieindlights[18]),
.OKT(ieindlights[19]),
.OKU(ieindlights[20]),
.OKV(ieindlights[21]),
.OKW(ieindlights[22]),
.OKX(ieindlights[23]));

  
mif mif0 (
.IAA(artoifviajb[0]),
.IAB(artoifviajb[1]),
.IAC(artoifviajb[2]),
.IAD(artoifviajb[3]),
.IAE(artoifviajb[4]),
.IAF(artoifviajb[5]),
.IAG(artoifviajb[6]),
.IAH(artoifviajb[7]),
.IAI(artoifviajb[8]),
.IAJ(artoifviajb[9]),
.IAK(artoifviajb[10]),
.IAL(artoifviajb[11]),
.IAM(artoifviajb[12]),
.IAN(artoifviajb[13]),
.IAO(artoifviajb[14]),
.IAP(artoifviajb[15]),
.IBA(artoifviajb[16]),
.IBB(artoifviajb[17]),
.IBC(artoifviajb[18]),
.IBD(artoifviajb[19]),
.IBE(artoifviajb[20]),
.IBF(artoifviajb[21]),
.IBG(artoifviajb[22]),
.IBH(artoifviajb[23]),
.IBI(artoifviajb[24]),
.IBJ(artoifviajb[25]),
.IBK(artoifviajb[26]),
.IBL(artoifviajb[27]),
.IBM(artoifviajb[28]),
.IBN(artoifviajb[29]),
.IBO(artoifviajb[30]),
.IBP(artoifviajb[31]),
.ICA(newpregtoif[0]),
.ICB(newpregtoif[1]),
.ICC(newpregtoif[2]),
.ICD(newpregtoif[3]),
.ICE(newpregtoif[4]),
.ICF(newpregtoif[5]),
.ICG(newpregtoif[6]),
.ICH(newpregtoif[7]),
.ICI(newpregtoif[8]),
.ICJ(newpregtoif[9]),
.ICK(newpregtoif[10]),
.ICL(newpregtoif[11]),
.ICM(newpregtoif[12]),
.ICN(newpregtoif[13]),
.ICO(newpregtoif[14]),
.ICP(newpregtoif[15]),
.IDA(newpregtoif[16]),
.IDB(newpregtoif[17]),
.IDC(newpregtoif[18]),
.IDD(newpregtoif[19]),
.IDE(newpregtoif[20]),
.IDF(newpregtoif[21]),
.IDG(newpregtoif[22]),
.IDH(newpregtoif[23]),
.IDI(newpregtoif[24]),
.IDJ(newpregtoif[25]),
.IDK(newpregtoif[26]),
.IDL(newpregtoif[27]),
.IDM(newpregtoif[28]),
.IDN(newpregtoif[29]),
.IDO(newpregtoif[30]),
.IDP(newpregtoif[31]),
.IEA(instpartoif[0]),
.IEB(instpartoif[1]),
.IEC(instpartoif[2]),
.IED(instpartoif[3]),
.IEE(instpartoif[4]),
.IEF(instpartoif[5]),
.IEG(instpartoif[6]),
.IEH(instpartoif[7]),
.IEI(instpartoif[8]),
.IEJ(instpartoif[9]),
.IEK(instpartoif[10]),
.IEL(instpartoif[11]),
.IEM(instpartoif[12]),
.IEN(instpartoif[13]),
.IEO(instpartoif[14]),
.IEP(instpartoif[15]),
.IFA(sregbrdata[0]),
.IFB(sregbrdata[1]),
.IFC(sregbrdata[2]),
.IFD(sregbrdata[3]),
.IFE(sregbrdata[4]),
.IFFF(sregbrdata[5]),
.IFG(sregbrdata[6]),
.IFH(sregbrdata[7]),
.IFI(vasregsign),
.IGA(arzerotesta),
.IGB(arzerotestb),
.IGC(arsigntest),
.IHB(boundaryflagtoif),
.IHC(fetchcompletetoif),
.IJA(goissuetoif[0]),
.IJB(goissuetoif[1]),
.IJC(advanceqif),
.IJD(conflicktchain),
.IKA(semaphorefl_3[0]),
.IKB(semaphorefl_3[1]),
.ILA(semaphorefromea[0]),
.ILB(semaphorefromea[1]),
.ILC(semaphorefromea[2]),
.IMA(deadstarttoif),
.IMB(interrupttoif),
.IMC(enterpfromea),
.IMD(enterbafromea),
.IME(enterlafromea),
.IMF(startfromea),
.IMG(enablecmrangetest),
.INA(phasetoif),
.IOA(quad0bufferbusy),
.IOB(quad1bufferbusy),
.IOC(quad2bufferbusy),
.IOD(quad3bufferbusy),
.IPA(vectlentoif[0]),
.IPB(vectlentoif[1]),
.IPC(vectlentoif[2]),
.IPD(vectlentoif[3]),
.IPE(vectlentoif[4]),
.IPF(vectlentoif[5]),
.IQA(iolentoif[0]),
.IQB(iolentoif[1]),
.IQC(iolentoif[2]),
.IQD(iolentoif[3]),
.IQE(iolentoif[4]),
.IQF(iolentoif[5]),
.IQG(externalseq[0]),
.IQH(externalseq[1]),
.IQI(refreshfromea),
.IZZ (sysclock),
.IZH(ihold),
.OAA(ifaddrtotf[0]),
.OAB(ifaddrtotf[1]),
.OAC(ifaddrtotf[2]),
.OAD(ifaddrtotf[3]),
.OAE(ifaddrtotf[4]),
.OAF(ifaddrtotf[5]),
.OAG(ifaddrtotf[6]),
.OAH(ifaddrtotf[7]),
.OAI(ifaddrtotf[8]),
.OAJ(ifaddrtotf[9]),
.OAK(ifaddrtotf[10]),
.OAL(ifaddrtotf[11]),
.OAM(ifaddrtotf[12]),
.OAN(ifaddrtotf[13]),
.OAO(ifaddrtotf[14]),
.OAP(ifaddrtotf[15]),
.OBA(ifaddrtotf[16]),
.OBB(ifaddrtotf[17]),
.OBC(ifaddrtotf[18]),
.OBD(ifaddrtotf[19]),
.OBE(ifaddrtotf[20]),
.OBF(ifaddrtotf[21]),
.OBG(ifaddrtotf[22]),
.OBH(ifaddrtotf[23]),
.OBI(ifaddrtotf[24]),
.OBJ(ifaddrtotf[25]),
.OBK(ifaddrtotf[26]),
.OBL(ifaddrtotf[27]),
.OBM(ifaddrtotf[28]),
.OBN(ifaddrtotf[29]),
.OBO(ifaddrtotf[30]),
.OBP(ifaddrtotf[31]),
.OCA(pregtoam[0]),
.OCB(pregtoam[1]),
.OCC(pregtoam[2]),
.OCD(pregtoam[3]),
.OCE(pregtoam[4]),
.OCF(pregtoam[5]),
.OCG(pregtoam[6]),
.OCH(pregtoam[7]),
.OCI(pregtoam[8]),
.OCJ(pregtoam[9]),
.OCK(pregtoam[10]),
.OCL(pregtoam[11]),
.OCM(pregtoam[12]),
.OCN(pregtoam[13]),
.OCO(pregtoam[14]),
.OCP(pregtoam[15]),
.ODA(pregtoam[16]),
.ODB(pregtoam[17]),
.ODC(pregtoam[18]),
.ODD(pregtoam[19]),
.ODE(pregtoam[20]),
.ODF(pregtoam[21]),
.ODG(pregtoam[22]),
.ODH(pregtoam[23]),
.ODI(pregtoam[24]),
.ODJ(pregtoam[25]),
.ODK(pregtoam[26]),
.ODL(pregtoam[27]),
.ODM(pregtoam[28]),
.ODN(pregtoam[29]),
.ODO(pregtoam[30]),
.ODP(pregtoam[31]),
.OEA(ifcontroltota[0]),
.OEB(ifcontroltota[1]),
.OEC(ifcontroltota[2]),
.OED(ifcontroltota[3]),
.OEE(ifcontroltota[4]),
.OEF(ifcontroltota[5]),
.OEG(ifcontroltota[6]),
.OEH(ifcontroltota[7]),
.OEI(ifcontroltota[8]),
.OEJ(ifcontroltota[9]),
.OEK(ifcontroltota[10]),
.OEL(ifcontroltota[11]),
.OEM(ifcontroltota[12]),
.OEN(ifcontroltota[13]),
.OEO(ifcontroltota[14]),
.OEP(ifcontroltota[15]),
.OEQ(ifcontroltota[16]),
.OER(ifcontroltota[17]),
.OES(ifcontroltota[18]),
.OET(ifcontroltota[19]),
.OEU(ifcontroltota[20]),
.OEV(ifcontroltota[21]),
.OEW(ifcontroltota[22]),
.OEX(ifcontroltota[23]),
.OEY(ifcontroltota[24]),
.OFA(gosdatatotb),
.OFB(goebdatatotb),
.OFC(retrytotb),
.OGA(artoifviajb[0]),
.OGB(artoifviajb[1]),
.OGC(artoifviajb[2]),
.OGD(artoifviajb[3]),
.OGE(artoifviajb[4]),
.OGF(artoifviajb[5]),
.OGG(artoifviajb[6]),
.OGH(artoifviajb[7]),
.OGI(artoifviajb[8]),
.OGJ(artoifviajb[9]),
.OGK(artoifviajb[10]),
.OGL(artoifviajb[11]),
.OGM(artoifviajb[12]),
.OGN(artoifviajb[13]),
.OGO(artoifviajb[14]),
.OGP(artoifviajb[15]),
.OHA(),
.OHB(),
.OHC(),
.OHD(),
.OHE(),
.OIA(branchpreambletoie),
.OIB(barreltesttoie),
.OIC(branchintoie),
.OID(branchouttoie),
.OIE(branchfallthrutoie),
.OIG(clearreadadr1),
.OJA(parcelptr[0]),
.OJB(parcelptr[1]),
.OJC(memportbusyfromif),
.OJD(holdissuefromif),
.OJE(gobranchfromif),
.OKA(semaphorefl_0[0]),
.OKB(semaphorefl_0[1]),
.OLA(setsematoea),
.OLB(clrsematoea),
.OLC(idletoea),
.OLD(exittoea),
.OLF(),
.OMA(holdadvtojb1),
.OMB(holdadvtojb2),
.OQA(gowritetoeb),
.OQB(endsequencetoeb),
.ORA(jkdatatoea[0]),
.ORB(jkdatatoea[1]),
.ORC(jkdatatoea[2]),
.ORD(jkdatatoea[3]),
.ORE(jkdatatoea[4]),
.ORF(jkdatatoea[5]),
.OTA(ifindlights[0]),
.OTB(ifindlights[1]),
.OTC(ifindlights[2]),
.OTD(ifindlights[3]),
.OTE(ifindlights[4]),
.OTF(ifindlights[5])
);

  
ja ja0 ( 
.IAA(ibufftoja[0]),
.IAB(ibufftoja[1]),
.IAC(ibufftoja[2]),
.IAD(ibufftoja[3]),
.IAE(ibufftoja[4]),
.IAF(ibufftoja[5]),
.IAG(ibufftoja[6]),
.IAH(ibufftoja[7]),
.IAI(ibufftoja[8]),
.IAJ(ibufftoja[9]),
.IAK(ibufftoja[10]),
.IAL(ibufftoja[11]),
.IAM(ibufftoja[12]),
.IAN(ibufftoja[13]),
.IAO(ibufftoja[14]),
.IAP(ibufftoja[15]),
.IBA(ibufftoja[16]),
.IBB(ibufftoja[17]),
.IBC(ibufftoja[18]),
.IBD(ibufftoja[19]),
.IBE(ibufftoja[20]),
.IBF(ibufftoja[21]),
.IBG(ibufftoja[22]),
.IBH(ibufftoja[23]),
.IBI(ibufftoja[24]),
.IBJ(ibufftoja[25]),
.IBK(ibufftoja[26]),
.IBL(ibufftoja[27]),
.IBM(ibufftoja[28]),
.IBN(ibufftoja[29]),
.IBO(ibufftoja[30]),
.IBP(ibufftoja[31]),
.ICA(ibufftoja[32]),
.ICB(ibufftoja[33]),
.ICC(ibufftoja[34]),
.ICD(ibufftoja[35]),
.ICE(ibufftoja[36]),
.ICF(ibufftoja[37]),
.ICG(ibufftoja[38]),
.ICH(ibufftoja[39]),
.ICI(ibufftoja[40]),
.ICJ(ibufftoja[41]),
.ICK(ibufftoja[42]),
.ICL(ibufftoja[43]),
.ICM(ibufftoja[44]),
.ICN(ibufftoja[45]),
.ICO(ibufftoja[46]),
.ICP(ibufftoja[47]),
.IDA(ibufftoja[48]),
.IDB(ibufftoja[49]),
.IDC(ibufftoja[50]),
.IDD(ibufftoja[51]),
.IDE(ibufftoja[52]),
.IDF(ibufftoja[53]),
.IDG(ibufftoja[54]),
.IDH(ibufftoja[55]),
.IDI(ibufftoja[56]),
.IDJ(ibufftoja[57]),
.IDK(ibufftoja[58]),
.IDL(ibufftoja[59]),
.IDM(ibufftoja[60]),
.IDN(ibufftoja[61]),
.IDO(ibufftoja[62]),
.IDP(ibufftoja[63]),
.IEA(vec0rel),
.IEB(vec1rel),
.IEC(vec2rel),
.IED(vec3rel),
.IEE(vec4rel),
.IEF(vec5rel),
.IEG(vec6rel),
.IEH(vec7rel),
.IFA(memdestja[0]),
.IFB(memdestja[1]),
.IFC(memdestja[2]),
.IFD(memdestja[3]),
.IGA(japarcel[0]),
.IGB(japarcel[1]),
.IJA(clrtoja[0]),
.IJB(clrtoja[1]),
.IJC(clrtoja[2]),
.IJD(clrtoja[3]),
.IJE(clrtoja[4]),
.IJJ(membsyja[0]),
.IJK(membsyja[1]),
//.IKA(datareadyja),
.IKA(iedataval),
//.IKB(gobranchfromif),
 .IKB(iedatahold),
.IKC(holdissueja),
.IKQ(deadstrtja),
.ILA(holdissueic),
.IZZ(sysclock),
.IZH(ihold),
.OAA(instpartoif[0]),
.OAB(instpartoif[1]),
.OAC(instpartoif[2]),
.OAD(instpartoif[3]),
.OAE(instpartoif[4]),
.OAF(instpartoif[5]),
.OAG(instpartoif[6]),
.OAH(instpartoif[7]),
.OAI(instpartoif[8]),
.OAJ(instpartoif[9]),
.OAK(instpartoif[10]),
.OAL(instpartoif[11]),
.OAM(instpartoif[12]),
.OAN(instpartoif[13]),
.OAO(instpartoif[14]),
.OAP(instpartoif[15]),
.OBA(instpartojb[0]),
.OBB(instpartojb[1]),
.OBC(instpartojb[2]),
.OBD(instpartojb[3]),
.OBE(instpartojb[4]),
.OBF(instpartojb[5]),
.OBG(instpartojb[6]),
.OBH(instpartojb[7]),
.OBI(instpartojb[8]),
.OBJ(instpartojb[9]),
.OBK(instpartojb[10]),
.OBL(instpartojb[11]),
.OBM(instpartojb[12]),
.OBN(instpartojb[13]),
.OBO(instpartojb[14]),
.OBP(instpartojb[15]),
.OCA(parceltowa[0]),
.OCB(parceltowa[1]),
.OCC(parceltowa[2]),
.OCD(parceltowa[3]),
.OCE(parceltowa[4]),
.OCF(parceltowa[5]),
.OCG(parceltowa[6]),
.OCH(parceltowa[7]),
.OCI(parceltowa[8]),
.OCJ(parceltowa[9]),
.OCK(parceltowa[10]),
.OCL(parceltowa[11]),
.OCM(parceltowa[12]),
.OCN(parceltowa[13]),
.OCO(parceltowa[14]),
.OCP(parceltowa[15]),
.ODA(goissuetoif[0]),
.ODB(goissuetojb[0]),
.ODC(goissuetojc0[0]),
.ODD(goissuetojc1[0]),
.ODE(goissuetowa[0]),
.ODF(goissuetoif[1]),
.ODG(goissuetojb[1]),
.ODH(goissuetojc0[1]),
.ODI(goissuetojc1[1]),
.ODJ(goissuetowa[1]),
.OEA(aregsrctoar[0]),
.OEB(aregsrctoar[1]),
.OEC(aregsrctoar[2]),
.OED(aregsrctoar[3]),
.OEE(aregsrctoar[4]),
.OEF(aregsrctoar[5]),
.OFA(sregsrctoam[0]),
.OFB(sregsrctoam[1]),
.OFC(sregsrctoam[2]),
.OFD(sregsrctoam[3]),
.OFE(sregsrctoam[4]),
.OFF(sregsrctoam[5]),
.OGA(arreadout[0]),
.OGB(arreadout[1]),
.OGC(arreadout[2]),
.OHA(vectorcodeam[0]),
.OHB(vectorcodeam[1]),
.OHC(vectorcodeam[2]),
.OHD(vectorcodeam[3]),
.OHE(vectorcodeam[4]),
.OHF(vectorcodeam[5]),
.OHG(vectorcodeam[6]),
.OIA(advanceqjb),
.OIB(advanceqif),
.OJA(subtracttoar),
.OJB(addtoar),
.OJC(enterltoar),
.OJD(goaddrmul),
.OKA(resumetoie),
.OLA(begvecttojc1[0]),
.OLB(begvecttojc1[1]),
.OLC(begvecttojc1[2]),
.OLD(begvecttojc1[3]),
.OLE(begvecttojc1[4]),
.OLF(begvecttojc1[5]),
.OLG(begvecttojc1[6]),
.OLH(begvecttojc1[7]),
.OMA(vectormode[0]),
.OMB(vectormode[1]),
.ONA(constreadwa),
.ONB(constwritewa),
.OOA(jagbcnt[0]),
.OOB(jagbcnt[1]),
.OOC(jagbcnt[2]),
.OOD(jagbcnt[3]),
.OOE(jagbcnt[4]),
.OOF(jagbcnt[5]),
.OPA(jagacnt[0]),
.OPB(jagacnt[1]),
.OPC(jagacnt[2]),
.OPD(jagacnt[3]),
.OQA(shftcontogb[0]),
.OQB(shftcontogb[1]),
.OQC(shftcontogb[2]),
.ORA(javacntr[0]),
.ORB(javacntr[1]),
.ORC(javacntr[2]),
.ORD(javacntr[3]),
.OSA(javbcntr[0]),
.OSB(javbcntr[1]),
.OSC(javbcntr[2]),
.OSD(javbcntr[3]),
.OSE(javbcntr[4]),
.OTA(javlcnt[0]),
.OTB(javlcnt[1]),
.OTC(javlcnt[2]),
.OTD(javlcnt[3]),
.OTE(javlcnt[4]),
.OTF(javlcnt[5]),
.OTG(javlcnt[6]),
.OUA(jafacnt[0]),
.OUB(jafacnt[1]),
.OUC(jafacnt[2]),
.OUD(jafacnt[3]),
.OUE(jafacnt[4]),
.OVA(jamecnt[0]),
.OVB(jamecnt[1]),
.OVC(jamecnt[2]),
.OVD(jamecnt[3]),
.OVE(jamecnt[4]),
.OVF(jamecnt[5]),
.OWA(gak0),
.OWB(indlightip[1]),
.OWC(indlightip[2]),
.OWD(indlightip[3]),
.OWE(indlightip[4]),
.OWF(indlightip[5]),
.OWG(indlightip[6]),
.OWH(indlightip[7]),
.OWI(indlightip[8]),
.OWJ(gaf0),
.OWK(gaf1),
.OWL(indlightip[11]),
.OWM(indlightip[12]),
.OWN(indlightip[13]),
.OWO(indlightip[14]),
.OWP(indlightip[15]),
.OWQ(indlightadvanceque),
.OWR(indlightlgoissue),
.OWS(indlightrankcfull),
.OWT(indlightrankefull),
.OWU(indlightgateparcel[0]),
.OWV(indlightgateparcel[1]),
.OWW(indlightgateparcel[2]),
.OWX(indlightgateparcel[3]),
.OXA(modechcnt[0]),
.OXB(modechcnt[1]),
.OXC(modechcnt[2]),
.OZA(jclocal[0]),
.OZB(jclocal[1]));


jb jb0( 
.IAA(arfanouttojb[0]),
.IAB(arfanouttojb[1]),
.IAC(arfanouttojb[2]),
.IAD(arfanouttojb[3]),
.IAE(arfanouttojb[4]),
.IAF(arfanouttojb[5]),
.IAG(arfanouttojb[6]),
.IAH(arfanouttojb[7]),
.IAI(arfanouttojb[8]),
.IAJ(arfanouttojb[9]),
.IAK(arfanouttojb[10]),
.IAL(arfanouttojb[11]),
.IAM(arfanouttojb[12]),
.IAN(arfanouttojb[13]),
.IAO(arfanouttojb[14]),
.IAP(arfanouttojb[15]),
.IBA(arfanouttojb[16]),
.IBB(arfanouttojb[17]),
.IBC(arfanouttojb[18]),
.IBD(arfanouttojb[19]),
.IBE(arfanouttojb[20]),
.IBF(arfanouttojb[21]),
.IBG(arfanouttojb[22]),
.IBH(arfanouttojb[23]),
.IBI(arfanouttojb[24]),
.IBJ(arfanouttojb[25]),
.IBK(arfanouttojb[26]),
.IBL(arfanouttojb[27]),
.IBM(arfanouttojb[28]),
.IBN(arfanouttojb[29]),
.IBO(arfanouttojb[30]),
.IBP(arfanouttojb[31]),
.ICA(instpartojb[0]),
.ICB(instpartojb[1]),
.ICC(instpartojb[2]),
.ICD(instpartojb[3]),
.ICE(instpartojb[4]),
.ICF(instpartojb[5]),
.ICG(instpartojb[6]),
.ICH(instpartojb[7]),
.ICI(instpartojb[8]),
.ICJ(instpartojb[9]),
.ICK(instpartojb[10]),
.ICL(instpartojb[11]),
.ICM(instpartojb[12]),
.ICN(instpartojb[13]),
.ICO(instpartojb[14]),
.ICP(instpartojb[15]),
.IDA(vectlentojb[0]),
.IDB(vectlentojb[1]),
.IDC(vectlentojb[2]),
.IDD(vectlentojb[3]),
.IDE(vectlentojb[4]),
.IDF(vectlentojb[5]),
.IEA(goissuetojb[0]),
.IEB(goissuetojb[1]),
.IFA(advanceqjb),
.IGA(phasetojb),
.IHA(deadstartjb),
.IJA(relvitojb),
.IKA(shregdatajb[0]),
.IKB(shregdatajb[1]),
.IKC(shregdatajb[2]),
.IKD(shregdatajb[3]),
.IKE(shregdatajb[4]),
.IKF(shregdatajb[5]),
.IKG(shregdatajb[6]),
.IKH(shregdatajb[7]),
.ILA(tailgatejb),
.IZZ (sysclock),
.IZH(ihold),
.OAA(jbtovr[0]),
.OAB(jbtovr[1]),
.OAC(jbtovr[2]),
.OAD(jbtovr[3]),
.OAE(jbtovr[4]),
.OAF(jbtovr[5]),
.OAG(jbtovr[6]),
.OAH(jbtovr[7]),
.OAI(jbtovr[8]),
.OAJ(jbtovr[9]),
.OAK(jbtovr[10]),
.OAL(jbtovr[11]),
.OAM(jbtovr[12]),
.OAN(jbtovr[13]),
.OAO(jbtovr[14]),
.OAP(jbtovr[15]),
.OBA(jbtovr[16]),
.OBB(jbtovr[17]),
.OBC(jbtovr[18]),
.OBD(jbtovr[19]),
.OBE(jbtovr[20]),
.OBF(jbtovr[21]),
.OBG(jbtovr[22]),
.OBH(jbtovr[23]),
.OBI(jbtovr[24]),
.OBJ(jbtovr[25]),
.OBK(jbtovr[26]),
.OBL(jbtovr[27]),
.OBM(jbtovr[28]),
.OBN(jbtovr[29]),
.OBO(jbtovr[30]),
.OBP(jbtovr[31]),
.OCA(jbtovr[32]),
.OCB(jbtovr[33]),
.OCC(jbtovr[34]),
.OCD(jbtovr[35]),
.OCE(jbtovr[36]),
.OCF(jbtovr[37]),
.OCG(jbtovr[38]),
.OCH(jbtovr[39]),
.OCI(jbtovr[40]),
.OCJ(jbtovr[41]),
.OCK(jbtovr[42]),
.OCL(jbtovr[43]),
.OCM(jbtovr[44]),
.OCN(jbtovr[45]),
.OCO(jbtovr[46]),
.OCP(jbtovr[47]),
.ODA(jbtovr[48]),
.ODB(jbtovr[49]),
.ODC(jbtovr[50]),
.ODD(jbtovr[51]),
.ODE(jbtovr[52]),
.ODF(jbtovr[53]),
.ODG(jbtovr[54]),
.ODH(jbtovr[55]),
.ODI(jbtovr[56]),
.ODJ(jbtovr[57]),
.ODK(jbtovr[58]),
.ODL(jbtovr[59]),
.ODM(jbtovr[60]),
.ODN(jbtovr[61]),
.ODO(jbtovr[62]),
.ODP(jbtovr[63]),
.OEA(jbatoar[0]),
.OEB(jbatoar[1]),
.OEC(jbatoar[2]),
.OED(jbatoar[3]),
.OEE(jbatoar[4]),
.OEF(jbatoar[5]),
.OEG(jbatoar[6]),
.OEH(jbatoar[7]),
.OEI(jbatoar[8]),
.OEJ(jbatoar[9]),
.OEK(jbatoar[10]),
.OEL(jbatoar[11]),
.OEM(jbatoar[12]),
.OEN(jbatoar[13]),
.OEO(jbatoar[14]),
.OEP(jbatoar[15]),
.OFA(jbatoar[16]),
.OFB(jbatoar[17]),
.OFC(jbatoar[18]),
.OFD(jbatoar[19]),
.OFE(jbatoar[20]),
.OFF(jbatoar[21]),
.OFG(jbatoar[22]),
.OFH(jbatoar[23]),
.OFI(jbatoar[24]),
.OFJ(jbatoar[25]),
.OFK(jbatoar[26]),
.OFL(jbatoar[27]),
.OFM(jbatoar[28]),
.OFN(jbatoar[29]),
.OFO(jbatoar[30]),
.OFP(jbatoar[31]),
.OGA(artoifviajb[0]),
.OGB(artoifviajb[1]),
.OGC(artoifviajb[2]),
.OGD(artoifviajb[3]),
.OGE(artoifviajb[4]),
.OGF(artoifviajb[5]),
.OGG(artoifviajb[6]),
.OGH(artoifviajb[7]),
.OGI(artoifviajb[8]),
.OGJ(artoifviajb[9]),
.OGK(artoifviajb[10]),
.OGL(artoifviajb[11]),
.OGM(artoifviajb[12]),
.OGN(artoifviajb[13]),
.OGO(artoifviajb[14]),
.OGP(artoifviajb[15]),
.OHA(artoifviajb[16]),
.OHB(artoifviajb[17]),
.OHC(artoifviajb[18]),
.OHD(artoifviajb[19]),
.OHE(artoifviajb[20]),
.OHF(artoifviajb[21]),
.OHG(artoifviajb[22]),
.OHH(artoifviajb[23]),
.OHI(artoifviajb[24]),
.OHJ(artoifviajb[25]),
.OHK(artoifviajb[26]),
.OHL(artoifviajb[27]),
.OHM(artoifviajb[28]),
.OHN(artoifviajb[29]),
.OHO(artoifviajb[30]),
.OHP(artoifviajb[31]),
.OIA(bwritetojc0[0]),
.OIB(bwritetojc0[1]),
.OIC(bwritetojc0[2]),
.OID(bwritetojc0[3]),
.OIE(bwritetojc1[0]),
.OIF(bwritetojc1[1]),
.OIG(bwritetojc1[2]),
.OIH(bwritetojc1[3]),
.OJA(phasejbtocm[0]),
.OJB(phasejbtocm[1]),
.OJC(phasejbtocm[2]),
.OJD(phasejbtocm[3]),
.OJE(phasejbtonxtjb),
.OJF(phasejbtotm[0]),
.OJG(phasejbtotm[1]),
.OJH(phasejbtotm[2]),
.OJI(phasejbtotm[3]),
.OJJ(phasejbtotm[4]),
.OJK(phasejbtotm[5]),
.OJL(phasejbtoas),
.OKA(clrtoja[0]),
.OKB(clrtoja[1]),
.OKC(clrtoja[2]),
.OKD(clrtoja[3]),
.OKE(clrtoja[4]),
.OKF(membsyja[0]),
.OLA(clearvectorlenvl),
.OLB(vectorenablefromjb),
.OLC(vectorlencntl),
.OLD(mefuenable),
.OLF(vectorshiftenable),
.OMA(jbindlight[0]),
.OMB(jbindlight[1]),
.OMC(jbindlight[2]),
.OMD(jbindlight[3]),
.OMF(jblengthlight[5]),
.ONA(jblengthlight[0]),
.ONB(jblengthlight[1]),
.ONC(jblengthlight[2]),
.OND(jblengthlight[3]),
.ONE(jblengthlight[4]),
.ONF(jblengthlight[5]),
.ORA(enteradtowa),
.ORB(entervrtowa),
.ORC(enterardtowa),
.ORD(advlmadrtowa),
.OSA(artoas[0]),
.OSB(artoas[1]),
.OSC(artoas[2]),
.OSD(artoas[3]),
.OSE(artoas[4]),
.OSF(artoas[5]),
.OSG(artoas[6]),
.OSH(artoas[7]),
.OTA(gosharedreg),
.OUA(shregoddeven),
.OUB(shregtype1),
.OUC(shregtype2));

jc jc0( 
.IAA(goissuetojc0[0]),
.IAB(goissuetojc0[1]),
.IBA(begvecttojc0[0]),
.IBB(begvecttojc0[1]),
.IBC(begvecttojc0[2]),
.IBD(begvecttojc0[3]),
.IBE(jclocal[0]),
.ICA(membackup2),
.ICB(holdadvjc[0]),
.IDA(bwritetojc0[0]),
.IDB(bwritetojc0[1]),
.IDC(bwritetojc0[2]),
.IDD(bwritetojc0[3]),
.IEA(memarivtojc0[0]),
.IEB(memarivtojc0[1]),
.IEC(memarivtojc0[2]),
.IED(memarivtojc0[3]),
.IEE(memarivtojc0[4]),
.IFA(vectlentojc0[0]),
.IFB(vectlentojc0[1]),
.IFC(vectlentojc0[2]),
.IFD(vectlentojc0[3]),
.IFE(vectlentojc0[4]),
.IFFF(vectlentojc0[5]),
.IGA(deadstartjc0),
.IHA(enableiota[0]),
.IHB(reliota[0]),
.IZZ (sysclock),
.OAA(v0addr1[0]),
.OAB(v0addr2[0]),
.OAC(v0addr3[0]),
.OAD(v0addr4[0]),
.OAE(v0addr5[0]),
.OAF(v0addr6[0]),
.OAG(v0addr7[0]),
.OAH(v0addr8[0]),
.OAI(v0addr1[1]),
.OAJ(v0addr2[1]),
.OAK(v0addr3[1]),
.OAL(v0addr4[1]),
.OAM(v0addr5[1]),
.OAN(v0addr6[1]),
.OAO(v0addr7[1]),
.OAP(v0addr8[1]),
.OBA(v0addr1[2]),
.OBB(v0addr2[2]),
.OBC(v0addr3[2]),
.OBD(v0addr4[2]),
.OBE(v0addr5[2]),
.OBF(v0addr6[2]),
.OBG(v0addr7[2]),
.OBH(v0addr8[2]),
.OBI(v0addr1[3]),
.OBJ(v0addr2[3]),
.OBK(v0addr3[3]),
.OBL(v0addr4[3]),
.OBM(v0addr5[3]),
.OBN(v0addr6[3]),
.OBO(v0addr7[3]),
.OBP(v0addr8[3]),
.OCA(v0addr1[4]),
.OCB(v0addr2[4]),
.OCC(v0addr3[4]),
.OCD(v0addr4[4]),
.OCE(v0addr5[4]),
.OCF(v0addr6[4]),
.OCG(v0addr7[4]),
.OCH(v0addr8[4]),
.OCI(v0addr1[5]),
.OCJ(v0addr2[5]),
.OCK(v0addr3[5]),
.OCL(v0addr4[5]),
.OCM(v0addr5[5]),
.OCN(v0addr6[5]),
.OCO(v0addr7[5]),
.OCP(v0addr8[5]),
.ODA(v0vectmode[0]),
.ODB(v0vectmode[1]),
.ODC(v0vectmode[2]),
.ODD(v0vectmode[3]),
.ODE(v0vectmode[4]),
.ODF(v0vectmode[5]),
.ODG(v0vectmode[6]),
.ODH(v0vectmode[7]),
.ODI(v0vectstep[0]),
.ODJ(v0vectstep[1]),
.ODK(v0vectstep[2]),
.ODL(v0vectstep[3]),
.ODM(v0vectstep[4]),
.ODN(v0vectstep[5]),
.ODO(v0vectstep[6]),
.ODP(v0vectstep[7]),
.OEA(v1addr1[0]),
.OEB(v1addr2[0]),
.OEC(v1addr3[0]),
.OED(v1addr4[0]),
.OEE(v1addr5[0]),
.OEF(v1addr6[0]),
.OEG(v1addr7[0]),
.OEH(v1addr8[0]),
.OEI(v1addr1[1]),
.OEJ(v1addr2[1]),
.OEK(v1addr3[1]),
.OEL(v1addr4[1]),
.OEM(v1addr5[1]),
.OEN(v1addr6[1]),
.OEO(v1addr7[1]),
.OEP(v1addr8[1]),
.OFA(v1addr1[2]),
.OFB(v1addr2[2]),
.OFC(v1addr3[2]),
.OFD(v1addr4[2]),
.OFE(v1addr5[2]),
.OFF(v1addr6[2]),
.OFG(v1addr7[2]),
.OFH(v1addr8[2]),
.OFI(v1addr1[3]),
.OFJ(v1addr2[3]),
.OFK(v1addr3[3]),
.OFL(v1addr4[3]),
.OFM(v1addr5[3]),
.OFN(v1addr6[3]),
.OFO(v1addr7[3]),
.OFP(v1addr8[3]),
.OGA(v1addr1[4]),
.OGB(v1addr2[4]),
.OGC(v1addr3[4]),
.OGD(v1addr4[4]),
.OGE(v1addr5[4]),
.OGF(v1addr6[4]),
.OGG(v1addr7[4]),
.OGH(v1addr8[4]),
.OGI(v1addr1[5]),
.OGJ(v1addr2[5]),
.OGK(v1addr3[5]),
.OGL(v1addr4[5]),
.OGM(v1addr5[5]),
.OGN(v1addr6[5]),
.OGO(v1addr7[5]),
.OGP(v1addr8[5]),
.OHA(v1vectmode[0]),
.OHB(v1vectmode[1]),
.OHC(v1vectmode[2]),
.OHD(v1vectmode[3]),
.OHE(v1vectmode[4]),
.OHF(v1vectmode[5]),
.OHG(v1vectmode[6]),
.OHH(v1vectmode[7]),
.OHI(v1vectstep[0]),
.OHJ(v1vectstep[1]),
.OHK(v1vectstep[2]),
.OHL(v1vectstep[3]),
.OHM(v1vectstep[4]),
.OHN(v1vectstep[5]),
.OHO(v1vectstep[6]),
.OHP(v1vectstep[7]),
.OIA(v2addr1[0]),
.OIB(v2addr2[0]),
.OIC(v2addr3[0]),
.OID(v2addr4[0]),
.OIE(v2addr5[0]),
.OIF(v2addr6[0]),
.OIG(v2addr7[0]),
.OIH(v2addr8[0]),
.OII(v2addr1[1]),
.OIJ(v2addr2[1]),
.OIK(v2addr3[1]),
.OIL(v2addr4[1]),
.OIM(v2addr5[1]),
.OIN(v2addr6[1]),
.OIO(v2addr7[1]),
.OIP(v2addr8[1]),
.OJA(v2addr1[2]),
.OJB(v2addr2[2]),
.OJC(v2addr3[2]),
.OJD(v2addr4[2]),
.OJE(v2addr5[2]),
.OJF(v2addr6[2]),
.OJG(v2addr7[2]),
.OJH(v2addr8[2]),
.OJI(v2addr1[3]),
.OJJ(v2addr2[3]),
.OJK(v2addr3[3]),
.OJL(v2addr4[3]),
.OJM(v2addr5[3]),
.OJN(v2addr6[3]),
.OJO(v2addr7[3]),
.OJP(v2addr8[3]),
.OKA(v2addr1[4]),
.OKB(v2addr2[4]),
.OKC(v2addr3[4]),
.OKD(v2addr4[4]),
.OKE(v2addr5[4]),
.OKF(v2addr6[4]),
.OKG(v2addr7[4]),
.OKH(v2addr8[4]),
.OKI(v2addr1[5]),
.OKJ(v2addr2[5]),
.OKK(v2addr3[5]),
.OKL(v2addr4[5]),
.OKM(v2addr5[5]),
.OKN(v2addr6[5]),
.OKO(v2addr7[5]),
.OKP(v2addr8[5]),
.OLA(v2vectmode[0]),
.OLB(v2vectmode[1]),
.OLC(v2vectmode[2]),
.OLD(v2vectmode[3]),
.OLE(v2vectmode[4]),
.OLF(v2vectmode[5]),
.OLG(v2vectmode[6]),
.OLH(v2vectmode[7]),
.OLI(v2vectstep[0]),
.OLJ(v2vectstep[1]),
.OLK(v2vectstep[2]),
.OLL(v2vectstep[3]),
.OLM(v2vectstep[4]),
.OLN(v2vectstep[5]),
.OLO(v2vectstep[6]),
.OLP(v2vectstep[7]),
.OMA(v3addr1[0]),
.OMB(v3addr2[0]),
.OMC(v3addr3[0]),
.OMD(v3addr4[0]),
.OME(v3addr5[0]),
.OMF(v3addr6[0]),
.OMG(v3addr7[0]),
.OMH(v3addr8[0]),
.OMI(v3addr1[1]),
.OMJ(v3addr2[1]),
.OMK(v3addr3[1]),
.OML(v3addr4[1]),
.OMM(v3addr5[1]),
.OMN(v3addr6[1]),
.OMO(v3addr7[1]),
.OMP(v3addr8[1]),
.ONA(v3addr1[2]),
.ONB(v3addr2[2]),
.ONC(v3addr3[2]),
.OND(v3addr4[2]),
.ONE(v3addr5[2]),
.ONF(v3addr6[2]),
.ONG(v3addr7[2]),
.ONH(v3addr8[2]),
.ONI(v3addr1[3]),
.ONJ(v3addr2[3]),
.ONK(v3addr3[3]),
.ONL(v3addr4[3]),
.ONM(v3addr5[3]),
.ONN(v3addr6[3]),
.ONO(v3addr7[3]),
.ONP(v3addr8[3]),
.OOA(v3addr1[4]),
.OOB(v3addr2[4]),
.OOC(v3addr3[4]),
.OOD(v3addr4[4]),
.OOE(v3addr5[4]),
.OOF(v3addr6[4]),
.OOG(v3addr7[4]),
.OOH(v3addr8[4]),
.OOI(v3addr1[5]),
.OOJ(v3addr2[5]),
.OOK(v3addr3[5]),
.OOL(v3addr4[5]),
.OOM(v3addr5[5]),
.OON(v3addr6[5]),
.OOO(v3addr7[5]),
.OOP(v3addr8[5]),
.OPA(v3vectmode[0]),
.OPB(v3vectmode[1]),
.OPC(v3vectmode[2]),
.OPD(v3vectmode[3]),
.OPE(v3vectmode[4]),
.OPF(v3vectmode[5]),
.OPG(v3vectmode[6]),
.OPH(v3vectmode[7]),
.OPI(v3vectstep[0]),
.OPJ(v3vectstep[1]),
.OPK(v3vectstep[2]),
.OPL(v3vectstep[3]),
.OPM(v3vectstep[4]),
.OPN(v3vectstep[5]),
.OPO(v3vectstep[6]),
.OPP(v3vectstep[7]),
.OQA(vec0rel),
.OQB(vec1rel),
.OQC(vec2rel),
.OQD(vec3rel));

  
jc jc1 ( 
.IAA(goissuetojc1[0]),
.IAB(goissuetojc1[1]),
.IBA(begvecttojc1[4]),
.IBB(begvecttojc1[5]),
.IBC(begvecttojc1[6]),
.IBD(begvecttojc1[7]),
.IBE(jclocal[1]),
.ICA(membackup3),
.ICB(holdadvjc[1]),
.IDA(bwritetojc1[0]),
.IDB(bwritetojc1[1]),
.IDC(bwritetojc1[2]),
.IDD(bwritetojc1[3]),
.IEA(memarivtojc1[0]),
.IEB(memarivtojc1[1]),
.IEC(memarivtojc1[2]),
.IED(memarivtojc1[3]),
.IEE(memarivtojc1[4]),
.IFA(vectlentojc1[0]),
.IFB(vectlentojc1[1]),
.IFC(vectlentojc1[2]),
.IFD(vectlentojc1[3]),
.IFE(vectlentojc1[4]),
.IFFF(vectlentojc1[5]),
.IGA(deadstartjc1),
.IHA(enableiota[1]),
.IHB(reliota[1]),
.IZZ (sysclock),
.OAA(v4addr1[0]),
.OAB(v4addr2[0]),
.OAC(v4addr3[0]),
.OAD(v4addr4[0]),
.OAE(v4addr5[0]),
.OAF(v4addr6[0]),
.OAG(v4addr7[0]),
.OAH(v4addr8[0]),
.OAI(v4addr1[1]),
.OAJ(v4addr2[1]),
.OAK(v4addr3[1]),
.OAL(v4addr4[1]),
.OAM(v4addr5[1]),
.OAN(v4addr6[1]),
.OAO(v4addr7[1]),
.OAP(v4addr8[1]),
.OBA(v4addr1[2]),
.OBB(v4addr2[2]),
.OBC(v4addr3[2]),
.OBD(v4addr4[2]),
.OBE(v4addr5[2]),
.OBF(v4addr6[2]),
.OBG(v4addr7[2]),
.OBH(v4addr8[2]),
.OBI(v4addr1[3]),
.OBJ(v4addr2[3]),
.OBK(v4addr3[3]),
.OBL(v4addr4[3]),
.OBM(v4addr5[3]),
.OBN(v4addr6[3]),
.OBO(v4addr7[3]),
.OBP(v4addr8[3]),
.OCA(v4addr1[4]),
.OCB(v4addr2[4]),
.OCC(v4addr3[4]),
.OCD(v4addr4[4]),
.OCE(v4addr5[4]),
.OCF(v4addr6[4]),
.OCG(v4addr7[4]),
.OCH(v4addr8[4]),
.OCI(v4addr1[5]),
.OCJ(v4addr2[5]),
.OCK(v4addr3[5]),
.OCL(v4addr4[5]),
.OCM(v4addr5[5]),
.OCN(v4addr6[5]),
.OCO(v4addr7[5]),
.OCP(v4addr8[5]),
.ODA(v4vectmode[0]),
.ODB(v4vectmode[1]),
.ODC(v4vectmode[2]),
.ODD(v4vectmode[3]),
.ODE(v4vectmode[4]),
.ODF(v4vectmode[5]),
.ODG(v4vectmode[6]),
.ODH(v4vectmode[7]),
.ODI(v4vectstep[0]),
.ODJ(v4vectstep[1]),
.ODK(v4vectstep[2]),
.ODL(v4vectstep[3]),
.ODM(v4vectstep[4]),
.ODN(v4vectstep[5]),
.ODO(v4vectstep[6]),
.ODP(v4vectstep[7]),
.OEA(v5addr1[0]),
.OEB(v5addr2[0]),
.OEC(v5addr3[0]),
.OED(v5addr4[0]),
.OEE(v5addr5[0]),
.OEF(v5addr6[0]),
.OEG(v5addr7[0]),
.OEH(v5addr8[0]),
.OEI(v5addr1[1]),
.OEJ(v5addr2[1]),
.OEK(v5addr3[1]),
.OEL(v5addr4[1]),
.OEM(v5addr5[1]),
.OEN(v5addr6[1]),
.OEO(v5addr7[1]),
.OEP(v5addr8[1]),
.OFA(v5addr1[2]),
.OFB(v5addr2[2]),
.OFC(v5addr3[2]),
.OFD(v5addr4[2]),
.OFE(v5addr5[2]),
.OFF(v5addr6[2]),
.OFG(v5addr7[2]),
.OFH(v5addr8[2]),
.OFI(v5addr1[3]),
.OFJ(v5addr2[3]),
.OFK(v5addr3[3]),
.OFL(v5addr4[3]),
.OFM(v5addr5[3]),
.OFN(v5addr6[3]),
.OFO(v5addr7[3]),
.OFP(v5addr8[3]),
.OGA(v5addr1[4]),
.OGB(v5addr2[4]),
.OGC(v5addr3[4]),
.OGD(v5addr4[4]),
.OGE(v5addr5[4]),
.OGF(v5addr6[4]),
.OGG(v5addr7[4]),
.OGH(v5addr8[4]),
.OGI(v5addr1[5]),
.OGJ(v5addr2[5]),
.OGK(v5addr3[5]),
.OGL(v5addr4[5]),
.OGM(v5addr5[5]),
.OGN(v5addr6[5]),
.OGO(v5addr7[5]),
.OGP(v5addr8[5]),
.OHA(v5vectmode[0]),
.OHB(v5vectmode[1]),
.OHC(v5vectmode[2]),
.OHD(v5vectmode[3]),
.OHE(v5vectmode[4]),
.OHF(v5vectmode[5]),
.OHG(v5vectmode[6]),
.OHH(v5vectmode[7]),
.OHI(v5vectstep[0]),
.OHJ(v5vectstep[1]),
.OHK(v5vectstep[2]),
.OHL(v5vectstep[3]),
.OHM(v5vectstep[4]),
.OHN(v5vectstep[5]),
.OHO(v5vectstep[6]),
.OHP(v5vectstep[7]),
.OIA(v6addr1[0]),
.OIB(v6addr2[0]),
.OIC(v6addr3[0]),
.OID(v6addr4[0]),
.OIE(v6addr5[0]),
.OIF(v6addr6[0]),
.OIG(v6addr7[0]),
.OIH(v6addr8[0]),
.OII(v6addr1[1]),
.OIJ(v6addr2[1]),
.OIK(v6addr3[1]),
.OIL(v6addr4[1]),
.OIM(v6addr5[1]),
.OIN(v6addr6[1]),
.OIO(v6addr7[1]),
.OIP(v6addr8[1]),
.OJA(v6addr1[2]),
.OJB(v6addr2[2]),
.OJC(v6addr3[2]),
.OJD(v6addr4[2]),
.OJE(v6addr5[2]),
.OJF(v6addr6[2]),
.OJG(v6addr7[2]),
.OJH(v6addr8[2]),
.OJI(v6addr1[3]),
.OJJ(v6addr2[3]),
.OJK(v6addr3[3]),
.OJL(v6addr4[3]),
.OJM(v6addr5[3]),
.OJN(v6addr6[3]),
.OJO(v6addr7[3]),
.OJP(v6addr8[3]),
.OKA(v6addr1[4]),
.OKB(v6addr2[4]),
.OKC(v6addr3[4]),
.OKD(v6addr4[4]),
.OKE(v6addr5[4]),
.OKF(v6addr6[4]),
.OKG(v6addr7[4]),
.OKH(v6addr8[4]),
.OKI(v6addr1[5]),
.OKJ(v6addr2[5]),
.OKK(v6addr3[5]),
.OKL(v6addr4[5]),
.OKM(v6addr5[5]),
.OKN(v6addr6[5]),
.OKO(v6addr7[5]),
.OKP(v6addr8[5]),
.OLA(v6vectmode[0]),
.OLB(v6vectmode[1]),
.OLC(v6vectmode[2]),
.OLD(v6vectmode[3]),
.OLE(v6vectmode[4]),
.OLF(v6vectmode[5]),
.OLG(v6vectmode[6]),
.OLH(v6vectmode[7]),
.OLI(v6vectstep[0]),
.OLJ(v6vectstep[1]),
.OLK(v6vectstep[2]),
.OLL(v6vectstep[3]),
.OLM(v6vectstep[4]),
.OLN(v6vectstep[5]),
.OLO(v6vectstep[6]),
.OLP(v6vectstep[7]),
.OMA(v7addr1[0]),
.OMB(v7addr2[0]),
.OMC(v7addr3[0]),
.OMD(v7addr4[0]),
.OME(v7addr5[0]),
.OMF(v7addr6[0]),
.OMG(v7addr7[0]),
.OMH(v7addr8[0]),
.OMI(v7addr1[1]),
.OMJ(v7addr2[1]),
.OMK(v7addr3[1]),
.OML(v7addr4[1]),
.OMM(v7addr5[1]),
.OMN(v7addr6[1]),
.OMO(v7addr7[1]),
.OMP(v7addr8[1]),
.ONA(v7addr1[2]),
.ONB(v7addr2[2]),
.ONC(v7addr3[2]),
.OND(v7addr4[2]),
.ONE(v7addr5[2]),
.ONF(v7addr6[2]),
.ONG(v7addr7[2]),
.ONH(v7addr8[2]),
.ONI(v7addr1[3]),
.ONJ(v7addr2[3]),
.ONK(v7addr3[3]),
.ONL(v7addr4[3]),
.ONM(v7addr5[3]),
.ONN(v7addr6[3]),
.ONO(v7addr7[3]),
.ONP(v7addr8[3]),
.OOA(v7addr1[4]),
.OOB(v7addr2[4]),
.OOC(v7addr3[4]),
.OOD(v7addr4[4]),
.OOE(v7addr5[4]),
.OOF(v7addr6[4]),
.OOG(v7addr7[4]),
.OOH(v7addr8[4]),
.OOI(v7addr1[5]),
.OOJ(v7addr2[5]),
.OOK(v7addr3[5]),
.OOL(v7addr4[5]),
.OOM(v7addr5[5]),
.OON(v7addr6[5]),
.OOO(v7addr7[5]),
.OOP(v7addr8[5]),
.OPA(v7vectmode[0]),
.OPB(v7vectmode[1]),
.OPC(v7vectmode[2]),
.OPD(v7vectmode[3]),
.OPE(v7vectmode[4]),
.OPF(v7vectmode[5]),
.OPG(v7vectmode[6]),
.OPH(v7vectmode[7]),
.OPI(v7vectstep[0]),
.OPJ(v7vectstep[1]),
.OPK(v7vectstep[2]),
.OPL(v7vectstep[3]),
.OPM(v7vectstep[4]),
.OPN(v7vectstep[5]),
.OPO(v7vectstep[6]),
.OPP(v7vectstep[7]),
.OQA(vec4rel),
.OQB(vec5rel),
.OQC(vec6rel),
.OQD(vec7rel));

ma ma0 (
.IAA(jopfotoma[0]),
.IAB(jopfotoma[1]),
.IAC(jopfotoma[2]),
.IAD(jopfotoma[3]),
.IAE(jopfotoma[4]),
.IAF(jopfotoma[5]),
.IAG(jopfotoma[6]),
.IAH(jopfotoma[7]),
.IAI(jopfotoma[8]),
.IAJ(jopfotoma[9]),
.IAK(jopfotoma[10]),
.IAL(jopfotoma[11]),
.IAM(jopfotoma[12]),
.IAN(jopfotoma[13]),
.IAO(jopfotoma[14]),
.IAP(jopfotoma[15]),
.IBA(kopfotoma[0]),
.IBB(kopfotoma[1]),
.IBC(kopfotoma[2]),
.IBD(kopfotoma[3]),
.IBE(kopfotoma[4]),
.IBF(kopfotoma[5]),
.IBG(kopfotoma[6]),
.IBH(kopfotoma[7]),
.IBI(kopfotoma[8]),
.IBJ(kopfotoma[9]),
.IBK(kopfotoma[10]),
.IBL(kopfotoma[11]),
.IBM(kopfotoma[12]),
.IBN(kopfotoma[13]),
.IBO(kopfotoma[14]),
.IBP(kopfotoma[15]),
.ICA(vrtomulj[16]),
.ICB(vrtomulj[17]),
.ICC(vrtomulj[18]),
.ICD(vrtomulj[19]),
.ICE(vrtomulj[20]),
.ICF(vrtomulj[21]),
.ICG(vrtomulj[22]),
.ICH(vrtomulj[23]),
.ICI(vrtomulj[24]),
.ICJ(vrtomulj[25]),
.ICK(vrtomulj[26]),
.ICL(vrtomulj[27]),
.ICM(vrtomulj[28]),
.ICN(vrtomulj[29]),
.ICO(vrtomulj[30]),
.ICP(vrtomulj[31]),
.IDA(vrtomulk[16]),
.IDB(vrtomulk[17]),
.IDC(vrtomulk[18]),
.IDD(vrtomulk[19]),
.IDE(vrtomulk[20]),
.IDF(vrtomulk[21]),
.IDG(vrtomulk[22]),
.IDH(vrtomulk[23]),
.IDI(vrtomulk[24]),
.IDJ(vrtomulk[25]),
.IDK(vrtomulk[26]),
.IDL(vrtomulk[27]),
.IDM(vrtomulk[28]),
.IDN(vrtomulk[29]),
.IDO(vrtomulk[30]),
.IDP(vrtomulk[31]),
.IEA(lufotoma[0]),
.IEB(lufotoma[1]),
.IEC(lufotoma[2]),
.IED(lufotoma[3]),
.IEE(lufotoma[4]),
.IEF(lufotoma[5]),
.IEG(lufotoma[6]),
.IEH(lufotoma[7]),
.IEI(lufotoma[8]),
.IEJ(lufotoma[9]),
.IEK(jopfotoma[32]),
.IEL(jopfotoma[33]),
.IEM(jopfotoma[34]),
.IEN(jopfotoma[35]),
.IEO(jopfotoma[36]),
.IEP(jopfotoma[37]),
.IEQ(jopfotoma[38]),
.IER(jopfotoma[39]),
.IES(jopfotoma[40]),
.IET(jopfotoma[41]),
.IEU(jopfotoma[42]),
.IEV(jopfotoma[43]),
.IEW(jopfotoma[44]),
.IEX(jopfotoma[45]),
.IEY(jopfotoma[46]),
.IEZ(jopfotoma[47]),
.IFA(kopfotoma[32]),
.IFB(kopfotoma[33]),
.IFC(kopfotoma[34]),
.IFD(kopfotoma[35]),
.IFE(kopfotoma[36]),
.IFFF(kopfotoma[37]),
.IFG(kopfotoma[38]),
.IFH(kopfotoma[39]),
.IFI(kopfotoma[40]),
.IFJ(kopfotoma[41]),
.IFK(kopfotoma[42]),
.IFL(kopfotoma[43]),
.IFM(kopfotoma[44]),
.IFN(kopfotoma[45]),
.IFO(kopfotoma[46]),
.IFP(kopfotoma[47]),
.IGA(magatekdatadel),
.IHA(maholdjdata),
.IKA(magatekdatatoj),
.IMM(mefloatrnd),
.IMR(mereciprnd),
.IMS(mesqrtrnd),
.IRA(masellookup),
.ISA(magatejdata),
.ITA(magatekdata),
.IZZ (sysclock),
.OAA(jopfotoma[16]),
.OAB(jopfotoma[17]),
.OAC(jopfotoma[18]),
.OAD(jopfotoma[19]),
.OAE(jopfotoma[20]),
.OAF(jopfotoma[21]),
.OAG(jopfotoma[22]),
.OAH(jopfotoma[23]),
.OAI(jopfotoma[24]),
.OAJ(jopfotoma[25]),
.OAK(jopfotoma[26]),
.OAL(jopfotoma[27]),
.OAM(jopfotoma[28]),
.OAN(jopfotoma[29]),
.OAO(jopfotoma[30]),
.OAP(jopfotoma[31]),
.OBA(jopfotomc[16]),
.OBB(jopfotomc[17]),
.OBC(jopfotomc[18]),
.OBD(jopfotomc[19]),
.OBE(jopfotomc[20]),
.OBF(jopfotomc[21]),
.OBG(jopfotomc[22]),
.OBH(jopfotomc[23]),
.OBI(jopfotomc[24]),
.OBJ(jopfotomc[25]),
.OBK(jopfotomc[26]),
.OBL(jopfotomc[27]),
.OBM(jopfotomc[28]),
.OBN(jopfotomc[29]),
.OBO(jopfotomc[30]),
.OBP(jopfotomc[31]),
.OCG(jopfotomd[22]),
.OCH(jopfotomd[23]),
.OCI(jopfotomd[24]),
.OCJ(jopfotomd[25]),
.OCK(jopfotomd[26]),
.OCL(jopfotomd[27]),
.OCM(jopfotomd[28]),
.OCN(jopfotomd[29]),
.OCO(jopfotomd[30]),
.OCP(jopfotomd[31]),
.ODA(kopfotoma[16]),
.ODB(kopfotoma[17]),
.ODC(kopfotoma[18]),
.ODD(kopfotoma[19]),
.ODE(kopfotoma[20]),
.ODF(kopfotoma[21]),
.ODG(kopfotoma[22]),
.ODH(kopfotoma[23]),
.ODI(kopfotoma[24]),
.ODJ(kopfotoma[25]),
.ODK(kopfotoma[26]),
.ODL(kopfotoma[27]),
.ODM(kopfotoma[28]),
.ODN(kopfotoma[29]),
.ODO(kopfotoma[30]),
.ODP(kopfotoma[31]),
.OEA(kopfotomc[16]),
.OEB(kopfotomc[17]),
.OEC(kopfotomc[18]),
.OED(kopfotomc[19]),
.OEE(kopfotomc[20]),
.OEF(kopfotomc[21]),
.OEG(kopfotomc[22]),
.OEH(kopfotomc[23]),
.OEI(kopfotomc[24]),
.OEJ(kopfotomc[25]),
.OEK(kopfotomc[26]),
.OEL(kopfotomc[27]),
.OEM(kopfotomc[28]),
.OEN(kopfotomc[29]),
.OEO(kopfotomc[30]),
.OEP(kopfotomc[31]),
.OFG(kopfotomd[22]),
.OFH(kopfotomd[23]),
.OFI(kopfotomd[24]),
.OFJ(kopfotomd[25]),
.OFK(kopfotomd[26]),
.OFL(kopfotomd[27]),
.OFM(kopfotomd[28]),
.OFN(kopfotomd[29]),
.OFO(kopfotomd[30]),
.OFP(kopfotomd[31]),
.OGA(mambflcar[0]),
.OGB(mambflcar[1]),
.OGC(mambflcar[2]),
.OGD(mambflcar[3]),
.OGE(mambflcar[4]),
.OGF(mambflcar[5]),
.OGG(mambflcar[6]),
.OGH(mambflcar[7]),
.OGI(mambflcar[8]),
.OGJ(mambflcar[9]),
.OGK(mambflcar[10]),
.OGL(mambflcar[11]),
.OGM(mambflcar[12]),
.OGN(mambflcar[13]),
.OGO(mambflcar[14]),
.OGP(mambflcar[15]),
.OHA(mambslcar[0]),
.OHB(mambslcar[1]),
.OHC(mambslcar[2]),
.OHD(mambslcar[3]),
.OHE(mambslcar[4]),
.OHF(mambslcar[5]),
.OHG(mambslcar[6]),
.OHH(mambslcar[7]),
.OHI(mambslcar[8]),
.OHJ(mambslcar[9]),
.OHK(mambslcar[10]),
.OIH(mambslcar[11]),
.OII(mambslcar[12]),
.OIJ(mambslcar[13]),
.OKA(mambtlcar[0]),
.OKB(mambtlcar[1]),
.OKC(mambtlcar[2]),
.OKD(mambtlcar[3]),
.OKE(mambtlcar[4]),
.OKF(mambtlcar[5]),
.OLD(mambtlcar[6]),
.OMA(mambftlcar[0]),
.OMB(mambftlcar[1]),
.ONB(mambftlcar[2]),
.OPK(marestomea[0]),
.OPM(marestomea[1]),
.OPO(marestomea[2]),
.OPQ(marestomea[3]),
.OPR(marestomea[4]),
.OQJ(marestomeb[0]),
.OQK(marestomeb[1]),
.OQM(marestomeb[2]),
.OQO(marestomeb[3]),
.OQQ(marestomeb[4]));


mb mb0 ( 
.IBA(jopfotoma[16]),
.IBB(jopfotoma[17]),
.IBC(jopfotoma[18]),
.IBD(jopfotoma[19]),
.IBE(jopfotoma[20]),
.IBF(jopfotoma[21]),
.IBG(jopfotoma[22]),
.IBH(jopfotoma[23]),
.IBI(jopfotoma[24]),
.IBJ(jopfotoma[25]),
.IBK(jopfotoma[26]),
.IBL(jopfotoma[27]),
.IBM(jopfotoma[28]),
.IBN(jopfotoma[29]),
.IBO(jopfotoma[30]),
.IBP(jopfotoma[31]),
.ICA(vrtomulj[0]),
.ICB(vrtomulj[1]),
.ICC(vrtomulj[2]),
.ICD(vrtomulj[3]),
.ICE(vrtomulj[4]),
.ICF(vrtomulj[5]),
.ICG(vrtomulj[6]),
.ICH(vrtomulj[7]),
.ICI(vrtomulj[8]),
.ICJ(vrtomulj[9]),
.ICK(vrtomulj[10]),
.ICL(vrtomulj[11]),
.ICM(vrtomulj[12]),
.ICN(vrtomulj[13]),
.ICO(vrtomulj[14]),
.ICP(vrtomulj[15]),
.IDA(vrtomulk[0]),
.IDB(vrtomulk[1]),
.IDC(vrtomulk[2]),
.IDD(vrtomulk[3]),
.IDE(vrtomulk[4]),
.IDF(vrtomulk[5]),
.IDG(vrtomulk[6]),
.IDH(vrtomulk[7]),
.IDI(vrtomulk[8]),
.IDJ(vrtomulk[9]),
.IDK(vrtomulk[10]),
.IDL(vrtomulk[11]),
.IDM(vrtomulk[12]),
.IDN(vrtomulk[13]),
.IDO(vrtomulk[14]),
.IDP(vrtomulk[15]),
.IEA(lufotomb[0]),
.IEB(lufotomb[1]),
.IEC(lufotomb[2]),
.IED(lufotomb[3]),
.IEE(lufotomb[4]),
.IEF(lufotomb[5]),
.IEG(lufotomb[6]),
.IEH(lufotomb[7]),
.IEI(lufotomb[8]),
.IEJ(lufotomb[9]),
.IEK(jopfotomb[32]),
.IEL(jopfotomb[33]),
.IEM(jopfotomb[34]),
.IEN(jopfotomb[35]),
.IEO(jopfotomb[36]),
.IEP(jopfotomb[37]),
.IEQ(jopfotomb[38]),
.IER(jopfotomb[39]),
.IES(jopfotomb[40]),
.IET(jopfotomb[41]),
.IEU(jopfotomb[42]),
.IEV(jopfotomb[43]),
.IEW(jopfotomb[44]),
.IEX(jopfotomb[45]),
.IEY(jopfotomb[46]),
.IEZ(jopfotomb[47]),
.IFA(kopfotoma[16]),
.IFB(kopfotoma[17]),
.IFC(kopfotoma[18]),
.IFD(kopfotoma[19]),
.IFE(kopfotoma[20]),
.IFFF(kopfotoma[21]),
.IFG(kopfotoma[22]),
.IFH(kopfotoma[23]),
.IFI(kopfotoma[24]),
.IFJ(kopfotoma[25]),
.IFK(kopfotoma[26]),
.IFL(kopfotoma[27]),
.IFM(kopfotoma[28]),
.IFN(kopfotoma[29]),
.IFO(kopfotoma[30]),
.IFP(kopfotoma[31]),
.IGA(kopfotomb[32]),
.IGB(kopfotomb[33]),
.IGC(kopfotomb[34]),
.IGD(kopfotomb[35]),
.IGE(kopfotomb[36]),
.IGF(kopfotomb[37]),
.IGG(kopfotomb[38]),
.IGH(kopfotomb[39]),
.IGI(kopfotomb[40]),
.IGJ(kopfotomb[41]),
.IGK(kopfotomb[42]),
.IGL(kopfotomb[43]),
.IGM(kopfotomb[44]),
.IGN(kopfotomb[45]),
.IGO(kopfotomb[46]),
.IGP(kopfotomb[47]),
.IHA(mbholdjdata),
.IIA(mbgatekdatadel),
.IKA(mbgatekdatatoj),
.ILA(mambflcar[0]),
.ILB(mambflcar[1]),
.ILC(mambflcar[2]),
.ILD(mambflcar[3]),
.ILE(mambflcar[4]),
.ILF(mambflcar[5]),
.ILG(mambflcar[6]),
.ILH(mambflcar[7]),
.ILI(mambflcar[8]),
.ILJ(mambflcar[9]),
.ILK(mambflcar[10]),
.ILL(mambflcar[11]),
.ILM(mambflcar[12]),
.ILN(mambflcar[13]),
.ILO(mambflcar[14]),
.ILP(mambflcar[15]),
.IMA(mambslcar[0]),
.IMB(mambslcar[1]),
.IMC(mambslcar[2]),
.IMD(mambslcar[3]),
.IME(mambslcar[4]),
.IMF(mambslcar[5]),
.IMG(mambslcar[6]),
.IMH(mambslcar[7]),
.IMI(mambslcar[8]),
.IMJ(mambslcar[9]),
.IMK(mambslcar[10]),
.IML(mambslcar[11]),
.IMM(mambslcar[12]),
.IMN(mambslcar[13]),
.INA(mambtlcar[0]),
.INB(mambtlcar[1]),
.INC(mambtlcar[2]),
.IND(mambtlcar[3]),
.INE(mambtlcar[4]),
.INF(mambtlcar[5]),
.ING(mambtlcar[6]),
.IOA(mambftlcar[0]),
.IOB(mambftlcar[1]),
.IOC(mambftlcar[2]),
.IRA(mbsellookup),
.ISA(mbgatejdata),
.ITA(mbgatekdata),
.ITB(mbitercntl),
.IZZ (sysclock),
.OAA(jopfotoma[0]),
.OAB(jopfotoma[1]),
.OAC(jopfotoma[2]),
.OAD(jopfotoma[3]),
.OAE(jopfotoma[4]),
.OAF(jopfotoma[5]),
.OAG(jopfotoma[6]),
.OAH(jopfotoma[7]),
.OAI(jopfotoma[8]),
.OAJ(jopfotoma[9]),
.OAK(jopfotoma[10]),
.OAL(jopfotoma[11]),
.OAM(jopfotoma[12]),
.OAN(jopfotoma[13]),
.OAO(jopfotoma[14]),
.OAP(jopfotoma[15]),
.OBL(jopfotomc[11]),
.OBM(jopfotomc[12]),
.OBN(jopfotomc[13]),
.OBO(jopfotomc[14]),
.OBP(jopfotomc[15]),
.OCA(kopfotoma[0]),
.OCB(kopfotoma[1]),
.OCC(kopfotoma[2]),
.OCD(kopfotoma[3]),
.OCE(kopfotoma[4]),
.OCF(kopfotoma[5]),
.OCG(kopfotoma[6]),
.OCH(kopfotoma[7]),
.OCI(kopfotoma[8]),
.OCJ(kopfotoma[9]),
.OCK(kopfotoma[10]),
.OCL(kopfotoma[11]),
.OCM(kopfotoma[12]),
.OCN(kopfotoma[13]),
.OCO(kopfotoma[14]),
.OCP(kopfotoma[15]),
.ODL(kopfotomc[11]),
.ODM(kopfotomc[12]),
.ODN(kopfotomc[13]),
.ODO(kopfotomc[14]),
.ODP(kopfotomc[15]),
.OGA(mbmcflcar[0]),
.OGB(mbmcflcar[1]),
.OGC(mbmcflcar[2]),
.OGD(mbmcflcar[3]),
.OGE(mbmcflcar[4]),
.OGF(mbmcflcar[5]),
.OGG(mbmcflcar[6]),
.OGH(mbmcflcar[7]),
.OGI(mbmcflcar[8]),
.OGJ(mbmcflcar[9]),
.OGK(mbmcflcar[10]),
.OGL(mbmcflcar[11]),
.OGM(mbmcflcar[12]),
.OHA(mbmcslcar[0]),
.OHB(mbmcslcar[1]),
.OHC(mbmcslcar[2]),
.OHD(mbmcslcar[3]),
.OHE(mbmcslcar[4]),
.OHF(mbmcslcar[5]),
.OHG(mbmcslcar[6]),
.OHH(mbmcslcar[7]),
.OHI(mbmcslcar[8]),
.OHJ(mbmcslcar[9]),
.OIG(mbmcftlcar[0]),
.OIH(mbmcftlcar[1]),
.OKA(mbmctlcar[0]),
.OKB(mbmctlcar[1]),
.OKC(mbmctlcar[2]),
.OKD(mbmctlcar[3]),
.OKE(mbmctlcar[4]),
.OLD(mbmctlcar[5]),
.OMA(mbmcfitlcar[0]),
.OMB(mbmcfitlcar[1]),
.OPA(mbrestomea[0]),
.OPB(mbrestomeb[0]),
.OPC(mbrestomea[1]),
.OPD(mbrestomeb[1]),
.OPE(mbrestomea[2]),
.OPF(mbrestomeb[2]),
.OPG(mbrestomea[3]),
.OPH(mbrestomeb[4]),
.OPI(mbrestomea[4]),
.OPK(mbrestomea[5]),
.OPM(mbrestomea[6]),
.OPO(mbrestomea[7]),
.OPQ(mbrestomea[8]),
.OPR(mbrestomea[9]),
.OQA(mbrestomec[1]),
.OQC(mbrestomec[2]),
.OQE(mbrestomec[3]),
.OQI(mbrestomeb[5]),
.OQK(mbrestomeb[6]),
.OQM(mbrestomeb[7]),
.OQO(mbrestomeb[8]),
.OQQ(mbrestomeb[9]));


mc mc0 ( 
.IAL(jopfotomc[11]),
.IAM(jopfotomc[12]),
.IAN(jopfotomc[13]),
.IAO(jopfotomc[14]),
.IAP(jopfotomc[15]),
.IBA(jopfotomc[16]),
.IBB(jopfotomc[17]),
.IBC(jopfotomc[18]),
.IBD(jopfotomc[19]),
.IBE(jopfotomc[20]),
.IBF(jopfotomc[21]),
.IBG(jopfotomc[22]),
.IBH(jopfotomc[23]),
.IBI(jopfotomc[24]),
.IBJ(jopfotomc[25]),
.IBK(jopfotomc[26]),
.IBL(jopfotomc[27]),
.IBM(jopfotomc[28]),
.IBN(jopfotomc[29]),
.IBO(jopfotomc[30]),
.IBP(jopfotomc[31]),
.ICA(jopfotomc[32]),
.ICB(jopfotomc[33]),
.ICC(jopfotomc[34]),
.ICD(jopfotomc[35]),
.ICE(jopfotomc[36]),
.ICF(jopfotomc[37]),
.ICG(jopfotomc[38]),
.ICH(jopfotomc[39]),
.ICI(jopfotomc[40]),
.ICJ(jopfotomc[41]),
.ICK(jopfotomc[42]),
.ICL(jopfotomc[43]),
.ICM(jopfotomc[44]),
.ICN(jopfotomc[45]),
.ICO(jopfotomc[46]),
.ICP(jopfotomc[47]),
.IDL(kopfotomc[11]),
.IDM(kopfotomc[12]),
.IDN(kopfotomc[13]),
.IDO(kopfotomc[14]),
.IDP(kopfotomc[15]),
.IEA(kopfotomc[16]),
.IEB(kopfotomc[17]),
.IEC(kopfotomc[18]),
.IED(kopfotomc[19]),
.IEE(kopfotomc[20]),
.IEF(kopfotomc[21]),
.IEG(kopfotomc[22]),
.IEH(kopfotomc[23]),
.IEI(kopfotomc[24]),
.IEJ(kopfotomc[25]),
.IEK(kopfotomc[26]),
.IEL(kopfotomc[27]),
.IEM(kopfotomc[28]),
.IEN(kopfotomc[29]),
.IEO(kopfotomc[30]),
.IEP(kopfotomc[31]),
.IFA(kopfotomc[32]),
.IFB(kopfotomc[33]),
.IFC(kopfotomc[34]),
.IFD(kopfotomc[35]),
.IFE(kopfotomc[36]),
.IFFF(kopfotomc[37]),
.IFG(kopfotomc[38]),
.IFH(kopfotomc[39]),
.IFI(kopfotomc[40]),
.IFJ(kopfotomc[41]),
.IFK(kopfotomc[42]),
.IFL(kopfotomc[43]),
.IFM(kopfotomc[44]),
.IFN(kopfotomc[45]),
.IFO(kopfotomc[46]),
.IFP(kopfotomc[47]),
.IGA(lufotomc[22]),
.IGB(lufotomc[23]),
.IGC(lufotomc[24]),
.IGD(lufotomc[25]),
.IGE(lufotomc[26]),
.IGF(lufotomc[27]),
.IGG(lufotomc[28]),
.IGH(lufotomc[29]),
.IGI(lufotomc[30]),
.IGJ(lufotomc[31]),
.ILA(mbmcflcar[0]),
.ILB(mbmcflcar[1]),
.ILC(mbmcflcar[2]),
.ILD(mbmcflcar[3]),
.ILE(mbmcflcar[4]),
.ILF(mbmcflcar[5]),
.ILG(mbmcflcar[6]),
.ILH(mbmcflcar[7]),
.ILI(mbmcflcar[8]),
.ILJ(mbmcflcar[9]),
.ILK(mbmcflcar[10]),
.ILL(mbmcflcar[11]),
.ILM(mbmcflcar[12]),
.IMA(mbmcslcar[0]),
.IMB(mbmcslcar[1]),
.IMC(mbmcslcar[2]),
.IMD(mbmcslcar[3]),
.IME(mbmcslcar[4]),
.IMF(mbmcslcar[5]),
.IMG(mbmcslcar[6]),
.IMH(mbmcslcar[7]),
.IMI(mbmcslcar[8]),
.IMJ(mbmcslcar[9]),
.IMK(mbmcftlcar[0]),
.IML(mbmcftlcar[1]),
.INA(mbmctlcar[0]),
.INB(mbmctlcar[1]),
.INC(mbmctlcar[2]),
.IND(mbmctlcar[3]),
.INE(mbmctlcar[4]),
.INF(mbmctlcar[5]),
.IOA(mbmcfitlcar[0]),
.IOB(mbmcfitlcar[1]),
.IQC(mchardrnd[0]),
.IQD(mchardrnd[1]),
.IQE(mchardrnd[2]),
.IQF(mchardrnd[3]),
.IQG(mchardrnd[4]),
.IQH(mchardrnd[5]),
.IRA(mcsellookup),
.IRB(mcitercntl),
.IRC(),
.IZZ (sysclock),
.OGA(mcmdflcar[0]),
.OGB(mcmdflcar[1]),
.OGC(mcmdflcar[2]),
.OGD(mcmdflcar[3]),
.OGE(mcmdflcar[4]),
.OGF(mcmdflcar[5]),
.OGG(mcmdflcar[6]),
.OGH(mcmdflcar[7]),
.OGI(mcmdflcar[8]),
.OHA(mcmdslcar[0]),
.OHB(mcmdslcar[1]),
.OHC(mcmdslcar[2]),
.OHD(mcmdslcar[3]),
.OHE(mcmdslcar[4]),
.OHF(mcmdslcar[5]),
.OIE(mcmdslcar[6]),
.OIF(mcmdslcar[7]),
.OKA(mcmdtlcar[0]),
.OKB(mcmdtlcar[1]),
.OKC(mcmdtlcar[2]),
.OLC(mcmdtlcar[3]),
.OMA(mcmdftlcar[0]),
.OMB(mcmdftlcar[1]),
.OPA(mcrestomea[10]),
.OPC(mcrestomea[9]),
.OPD(mcrestomeb[9]),
.OPE(mcrestomea[8]),
.OPF(mcrestomeb[8]),
.OPG(mcrestomea[7]),
.OPI(mcrestomea[6]),
.OPK(mcrestomea[5]),
.OPM(mcrestomea[4]),
.OPO(mcrestomea[3]),
.OPQ(mcrestomea[2]),
.OPS(mcrestomea[1]),
.OPU(mcrestomea[0]),
.OQA(mcrestomec[9]),
.OQC(mcrestomec[8]),
.OQD(mcrestomec[7]),
.OQG(mcrestomeb[6]),
.OQI(mcrestomeb[5]),
.OQK(mcrestomeb[4]),
.OQM(mcrestomeb[3]),
.OQO(mcrestomeb[2]),
.OQQ(mcrestomeb[1]),
.OQS(mcrestomeb[0]),
.OQU(mccotwoseven));
  
md md0 ( 
.IAA(lufotomd[0]),
.IAB(lufotomd[1]),
.IAC(lufotomd[2]),
.IAD(lufotomd[3]),
.IAE(lufotomd[4]),
.IAF(lufotomd[5]),
.IAG(lufotomd[6]),
.IAH(lufotomd[7]),
.IAI(lufotomd[8]),
.IAJ(lufotomd[9]),
.IAK(jopfotomd[32]),
.IAL(jopfotomd[33]),
.IAM(jopfotomd[34]),
.IAN(jopfotomd[35]),
.IAO(jopfotomd[36]),
.IAP(jopfotomd[37]),
.IAQ(jopfotomd[38]),
.IAR(jopfotomd[39]),
.IAS(jopfotomd[40]),
.IAT(jopfotomd[41]),
.IAU(jopfotomd[42]),
.IAV(jopfotomd[43]),
.IAW(jopfotomd[44]),
.IAX(jopfotomd[45]),
.IAY(jopfotomd[46]),
.IAZ(jopfotomd[47]),
.IBA(kopfotomd[22]),
.IBB(kopfotomd[23]),
.IBC(kopfotomd[24]),
.IBD(kopfotomd[25]),
.IBE(kopfotomd[26]),
.IBF(kopfotomd[27]),
.IBG(kopfotomd[28]),
.IBH(kopfotomd[29]),
.IBI(kopfotomd[30]),
.IBJ(kopfotomd[31]),
.IBK(kopfotomd[32]),
.IBL(kopfotomd[33]),
.IBM(kopfotomd[34]),
.IBN(kopfotomd[35]),
.IBO(kopfotomd[36]),
.IBP(kopfotomd[37]),
.IBQ(kopfotomd[38]),
.IBR(kopfotomd[39]),
.IBS(kopfotomd[40]),
.IBT(kopfotomd[41]),
.IBU(kopfotomd[42]),
.IBV(kopfotomd[43]),
.IBW(kopfotomd[44]),
.IBX(kopfotomd[45]),
.IBY(kopfotomd[46]),
.IBZ(kopfotomd[47]),
.ICA(jopfotomd[22]),
.ICB(jopfotomd[23]),
.ICC(jopfotomd[24]),
.ICD(jopfotomd[25]),
.ICE(jopfotomd[26]),
.ICF(jopfotomd[27]),
.ICG(jopfotomd[28]),
.ICH(jopfotomd[29]),
.ICI(jopfotomd[30]),
.ICJ(jopfotomd[31]),
.IIA(mditercntl),
.IKA(mdludata[0]),
.IKB(mdludata[1]),
.IKC(mdludata[2]),
.IKD(mdludata[3]),
.IKE(mdludata[4]),
.IKF(mdludata[5]),
.IKG(mdludata[6]),
.IKH(mdludata[7]),
.IKI(mdludata[8]),
.IKJ(mdludata[9]),
.IKK(mdludata[10]),
.IKL(mdludata[11]),
.IKM(mdludata[12]),
.ILA(mcmdflcar[0]),
.ILB(mcmdflcar[1]),
.ILC(mcmdflcar[2]),
.ILD(mcmdflcar[3]),
.ILE(mcmdflcar[4]),
.ILF(mcmdflcar[5]),
.ILG(mcmdflcar[6]),
.ILH(mcmdflcar[7]),
.ILI(mcmdflcar[8]),
.IMA(mcmdslcar[0]),
.IMB(mcmdslcar[1]),
.IMC(mcmdslcar[2]),
.IMD(mcmdslcar[3]),
.IME(mcmdslcar[4]),
.IMF(mcmdslcar[5]),
.IMG(mcmdslcar[6]),
.IMH(mcmdslcar[7]),
.INA(mcmdtlcar[0]),
.INB(mcmdtlcar[1]),
.INC(mcmdtlcar[2]),
.IND(mcmdtlcar[3]),
.IOA(mcmdftlcar[0]),
.IOB(mcmdftlcar[1]),
.IRA(mdsellookup),
.ISA(mdrndbit[0]),
.ISB(mdrndbit[1]),
.ISC(mdrndbit[2]),
.ITA(mdselsqrtsh),
.IZZ (sysclock),
.OAA(mdrestomea[26]),
.OAM(mdrestomeb[25]),
.OBA(mdrestomea[25]),
.OBM(mdrestomeb[24]),
.OCA(mdrestomea[24]),
.OCM(mdrestomeb[23]),
.ODA(mdrestomea[23]),
.OEA(mdrestomea[22]),
.OEB(mdrestomeb[22]),
.OFA(mdrestomea[21]),
.OFB(mdrestomeb[21]),
.OGA(mdrestomea[20]),
.OGB(mdrestomeb[20]),
.OHA(mdrestomea[19]),
.OHB(mdrestomeb[19]),
.OIA(mdrestomea[18]),
.OIB(mdrestomeb[18]),
.OJA(mdrestomea[17]),
.OJB(mdrestomeb[17]),
.OKA(mdrestomea[16]),
.OKB(mdrestomeb[16]),
.OLA(mdrestomea[15]),
.OLB(mdrestomeb[15]),
.OMA(mdrestomea[14]),
.OMB(mdrestomeb[14]),
.ONA(mdrestomea[13]),
.ONB(mdrestomeb[13]),
.OOA(mdrestomea[12]),
.OOB(mdrestomeb[12]),
.OPA(mdrestomea[11]),
.OPB(mdrestomeb[11]),
.OQA(mdrestomea[10]),
.OQB(mdrestomeb[10]),
.ORA(mdrestomea[9]),
.ORB(mdrestomeb[9]),
.OSA(mdrestomea[8]),
.OSB(mdrestomeb[8]),
.OTA(mdrestomea[7]),
.OTB(mdrestomeb[7]),
.OUA(mdrestomea[6]),
.OUB(mdrestomeb[6]),
.OVA(mdrestomea[5]),
.OVB(mdrestomeb[5]),
.OWA(mdrestomea[4]),
.OWB(mdrestomeb[4]),
.OXA(mdrestomea[3]),
.OXB(mdrestomeb[3]),
.OYA(mdrestomea[2]),
.OYB(mdrestomeb[2]),
.OZA(mdrestomea[1]),
.OZB(mdrestomeb[1]),
.OZM(mdrestomea[0]),
.OZN(mdrestomeb[0]));


me me0 ( 
.IAB(),
.IAC(marestomea[0]),
.IAD(marestomea[1]),
.IAE(marestomea[2]),
.IAF(marestomea[3]),
.IAG(mbrestomea[0]),
.IAH(mbrestomea[1]),
.IAI(mbrestomea[2]),
.IAJ(mbrestomea[3]),
.IAK(mbrestomea[4]),
.IAL(mbrestomea[5]),
.IAM(mbrestomea[6]),
.IAN(mbrestomea[7]),
.IAO(mbrestomea[8]),
.IAP(mcrestomea[10]),
.IAQ(mcrestomea[9]),
.IAR(mcrestomea[8]),
.IAS(mcrestomea[7]),
.IAT(mcrestomea[6]),
.IAU(mcrestomea[5]),
.IAV(mcrestomea[4]),
.IAW(mcrestomea[3]),
.IAX(mcrestomea[2]),
.IAY(mcrestomea[1]),
.IAZ(mcrestomea[0]),
.IBA(mdrestomea[26]),
.IBB(mdrestomea[25]),
.IBC(mdrestomea[24]),
.IBD(mdrestomea[23]),
.IBE(mdrestomea[22]),
.IBF(mdrestomea[21]),
.IBG(mdrestomea[20]),
.IBH(mdrestomea[19]),
.IBI(mdrestomea[18]),
.IBJ(mdrestomea[17]),
.IBK(mdrestomea[16]),
.IBL(mdrestomea[15]),
.IBM(mdrestomea[14]),
.IBN(mdrestomea[13]),
.IBO(mdrestomea[12]),
.IBP(mdrestomea[11]),
.IBQ(mdrestomea[10]),
.IBR(mdrestomea[9]),
.IBS(mdrestomea[8]),
.IBT(mdrestomea[7]),
.IBU(mdrestomea[6]),
.IBV(mdrestomea[5]),
.IBW(mdrestomea[4]),
.IBX(mdrestomea[3]),
.IBY(mdrestomea[2]),
.IBZ(mdrestomea[1]),
.ICB(marestomeb[0]),
.ICC(marestomeb[0]),
.ICD(marestomeb[1]),
.ICE(marestomeb[2]),
.ICF(marestomeb[3]),
.ICG(marestomea[4]),
.ICH(mbrestomeb[1]),
.ICI(mbrestomeb[2]),
.ICK(mbrestomeb[4]),
.ICL(mbrestomeb[5]),
.ICM(mbrestomeb[6]),
.ICN(mbrestomeb[7]),
.ICO(mbrestomeb[8]),
.ICP(mbrestomeb[9]),
.ICQ(mcrestomeb[9]),
.ICR(mcrestomec[7]),
.ICS(mcrestomeb[8]),
.ICT(mcrestomeb[6]),
.ICU(mcrestomeb[5]),
.ICV(mcrestomeb[4]),
.ICW(mcrestomeb[3]),
.ICX(mcrestomeb[2]),
.ICY(mcrestomeb[1]),
.ICZ(mcrestomeb[0]),
.IDA(mccotwoseven),
.IDB(mdrestomeb[25]),
.IDC(mdrestomeb[24]),
.IDD(mdrestomeb[23]),
.IDE(mdrestomeb[22]),
.IDF(mdrestomeb[21]),
.IDG(mdrestomeb[20]),
.IDH(mdrestomeb[19]),
.IDI(mdrestomeb[18]),
.IDJ(mdrestomeb[17]),
.IDK(mdrestomeb[16]),
.IDL(mdrestomeb[15]),
.IDM(mdrestomeb[14]),
.IDN(mdrestomeb[13]),
.IDO(mdrestomeb[12]),
.IDP(mdrestomeb[11]),
.IDQ(mdrestomeb[10]),
.IDR(mdrestomeb[9]),
.IDS(mdrestomeb[8]),
.IDT(mdrestomeb[7]),
.IDU(mdrestomeb[6]),
.IDV(mdrestomeb[5]),
.IDW(mdrestomeb[4]),
.IDX(mdrestomeb[3]),
.IDY(mdrestomeb[2]),
.IDZ(mdrestomeb[1]),
.IEF(marestomeb[3]),
.IEG(marestomeb[4]),
.IEH(mbrestomec[1]),
.IEI(mbrestomec[2]),
.IEO(mbrestomea[9]),
.IEP(mbrestomea[9]),
.IEQ(mcrestomec[9]),
.IER(mcrestomec[8]),
.IFFF(mbrestomeb[0]),
.IGA(vrtomulj[48]),
.IGB(vrtomulj[49]),
.IGC(vrtomulj[50]),
.IGD(vrtomulj[51]),
.IGE(vrtomulj[52]),
.IGF(vrtomulj[53]),
.IGG(vrtomulj[54]),
.IGH(vrtomulj[55]),
.IGI(vrtomulj[56]),
.IGJ(vrtomulj[57]),
.IGK(vrtomulj[58]),
.IGL(vrtomulj[59]),
.IGM(vrtomulj[60]),
.IGN(vrtomulj[61]),
.IGO(vrtomulj[62]),
.IGP(vrtomulj[63]),
.IHA(vrtomulk[48]),
.IHB(vrtomulk[49]),
.IHC(vrtomulk[50]),
.IHD(vrtomulk[51]),
.IHE(vrtomulk[52]),
.IHF(vrtomulk[53]),
.IHG(vrtomulk[54]),
.IHH(vrtomulk[55]),
.IHI(vrtomulk[56]),
.IHJ(vrtomulk[57]),
.IHK(vrtomulk[58]),
.IHL(vrtomulk[59]),
.IHM(vrtomulk[60]),
.IHN(vrtomulk[61]),
.IHO(vrtomulk[62]),
.IHP(vrtomulk[63]),
.IUA(mefuenable),
.IUB(enablefmrangeerr),
.IVA(wajamecnt[0]),
.IVB(wajamecnt[1]),
.IVC(wajamecnt[2]),
.IVD(wajamecnt[3]),
.IVE(wajamecnt[4]),
.IVF(wajamecnt[5]),
.IWA(mdrestomea[0]),
.IWB(mdrestomeb[0]),
.IZZ (sysclock),
.OAA(),
.OAB(metovr[0]),
.OAC(metovr[1]),
.OAD(metovr[2]),
.OAE(metovr[3]),
.OAF(metovr[4]),
.OAG(metovr[5]),
.OAH(metovr[6]),
.OAI(metovr[7]),
.OAJ(metovr[8]),
.OAK(metovr[9]),
.OAL(metovr[10]),
.OAM(metovr[11]),
.OAN(metovr[12]),
.OAO(metovr[13]),
.OAP(metovr[14]),
.OAQ(metovr[15]),
.OAR(metovr[16]),
.OAS(metovr[17]),
.OAT(metovr[18]),
.OAU(metovr[19]),
.OAV(metovr[20]),
.OAW(metovr[21]),
.OAX(metovr[22]),
.OBA(metovr[23]),
.OBB(metovr[24]),
.OBC(metovr[25]),
.OBD(metovr[26]),
.OBE(metovr[27]),
.OBF(metovr[28]),
.OBG(metovr[29]),
.OBH(metovr[30]),
.OBI(metovr[31]),
.OBJ(metovr[32]),
.OBK(metovr[33]),
.OBL(metovr[34]),
.OBM(metovr[35]),
.OBN(metovr[36]),
.OBO(metovr[37]),
.OBP(metovr[38]),
.OBQ(metovr[39]),
.OBR(metovr[40]),
.OBS(metovr[41]),
.OBT(metovr[42]),
.OBU(metovr[43]),
.OBV(metovr[44]),
.OBW(metovr[45]),
.OBX(metovr[46]),
.OBY(metovr[47]),
.OCA(metovr[48]),
.OCB(metovr[49]),
.OCC(metovr[50]),
.OCD(metovr[51]),
.OCE(metovr[52]),
.OCF(metovr[53]),
.OCG(metovr[54]),
.OCH(metovr[55]),
.OCI(metovr[56]),
.OCJ(metovr[57]),
.OCK(metovr[58]),
.OCL(metovr[59]),
.OCM(metovr[60]),
.OCN(metovr[61]),
.OCO(metovr[62]),
.OCP(metovr[63]),
.ODA(magatekdata),
.ODB(mbgatekdata),
.ODC(ragatekdata),
.OEA(magatekdatatoj),
.OEB(mbgatekdatatoj),
.OEC(ragatekdatatoj),
.OFA(maholdjdata),
.OFB(mbholdjdata),
.OFC(raholdjdata),
.OGA(magatejdata),
.OGB(mbgatejdata),
.OGC(ragatejdata),
.OHA(magatekdatadel),
.OHB(mbgatekdatadel),
.OHC(ragatekdatadel),
.OIA(mbsellookup),
.OIB(masellookup),
.OIC(mcsellookup),
.OID(mdsellookup),
.OJA(mefloatrnd),
.OJB(mereciprnd),
.OJC(mesqrtrnd),
.OJD(mbitercntl),
.OJE(mcitercntl),
.OJF(mditercntl),
.OKA(mdselsqrtsh),
.OLA(fprangeerrme),
.OMA(),
.OMB(ragaterecip),
.OMC(raselrecip),
.OMD(ragatesqrthardround));

ra ra0 (
.IAA(vrtomulj[32]),
.IAB(vrtomulj[33]),
.IAC(vrtomulj[34]),
.IAD(vrtomulj[35]),
.IAE(vrtomulj[36]),
.IAF(vrtomulj[37]),
.IAG(vrtomulj[38]),
.IAH(vrtomulj[39]),
.IAI(vrtomulj[40]),
.IAJ(vrtomulj[41]),
.IAK(vrtomulj[42]),
.IAL(vrtomulj[43]),
.IAM(vrtomulj[44]),
.IAN(vrtomulj[45]),
.IAO(vrtomulj[46]),
.IAP(vrtomulj[47]),
.ICA(vrtomulk[32]),
.ICB(vrtomulk[33]),
.ICC(vrtomulk[34]),
.ICD(vrtomulk[35]),
.ICE(vrtomulk[36]),
.ICF(vrtomulk[37]),
.ICG(vrtomulk[38]),
.ICH(vrtomulk[39]),
.ICI(vrtomulk[40]),
.ICJ(vrtomulk[41]),
.ICK(vrtomulk[42]),
.ICL(vrtomulk[43]),
.ICM(vrtomulk[44]),
.ICN(vrtomulk[45]),
.ICO(vrtomulk[46]),
.ICP(vrtomulk[47]),
.IGA(luoddevenadd),
.IJA(ragatesqrthardround),
.IKA(deadstartra),
.ILA(kaconsoletora[0]),
.ILB(kaconsoletora[1]),
.ILC(kaconsoletora[2]),
.ILD(kaconsoletora[3]),
.ILE(kaconsoletora[4]),
.ILF(kaconsoletora[5]),
.ILG(kaconsoletora[6]),
.ILH(kaconsoletora[7]),
.ILI(raloadbyte),
.IPA(ragatekdata),
.IPB(ragatekdatadel),
.IQA(ragatejdata),
.IQB(raholdjdata),
.IQC(ragatekdatatoj),
.IRA(raselrecip),
.IRB(ragaterecip),
.ISA(ragatesqrt),
.IZZ (sysclock),
.OAA(lufotoma[0]),
.OAB(lufotoma[1]),
.OAC(lufotoma[2]),
.OAD(lufotoma[3]),
.OAE(lufotoma[4]),
.OAF(lufotoma[5]),
.OAG(lufotoma[6]),
.OAH(lufotoma[7]),
.OAI(lufotoma[8]),
.OAJ(lufotoma[9]),
.OAK(jopfotoma[32]),
.OAL(jopfotoma[33]),
.OAM(jopfotoma[34]),
.OAN(jopfotoma[35]),
.OAO(jopfotoma[36]),
.OAP(jopfotoma[37]),
.OAQ(jopfotoma[38]),
.OAR(jopfotoma[39]),
.OAS(jopfotoma[40]),
.OAT(jopfotoma[41]),
.OAU(jopfotoma[42]),
.OAV(jopfotoma[43]),
.OAW(jopfotoma[44]),
.OAX(jopfotoma[45]),
.OAY(jopfotoma[46]),
.OAZ(jopfotoma[47]),
.OBA(lufotomb[0]),
.OBB(lufotomb[1]),
.OBC(lufotomb[2]),
.OBD(lufotomb[3]),
.OBE(lufotomb[4]),
.OBF(lufotomb[5]),
.OBG(lufotomb[6]),
.OBH(lufotomb[7]),
.OBI(lufotomb[8]),
.OBJ(lufotomb[9]),
.OBK(jopfotomb[32]),
.OBL(jopfotomb[33]),
.OBM(jopfotomb[34]),
.OBN(jopfotomb[35]),
.OBO(jopfotomb[36]),
.OBP(jopfotomb[37]),
.OBQ(jopfotomb[38]),
.OBR(jopfotomb[39]),
.OBS(jopfotomb[40]),
.OBT(jopfotomb[41]),
.OBU(jopfotomb[42]),
.OBV(jopfotomb[43]),
.OBW(jopfotomb[44]),
.OBX(jopfotomb[45]),
.OBY(jopfotomb[46]),
.OBZ(jopfotomb[47]),
.OCA(lufotomc[22]),
.OCB(lufotomc[23]),
.OCC(lufotomc[24]),
.OCD(lufotomc[25]),
.OCE(lufotomc[26]),
.OCF(lufotomc[27]),
.OCG(lufotomc[28]),
.OCH(lufotomc[29]),
.OCI(lufotomc[30]),
.OCJ(lufotomc[31]),
.OCK(jopfotomc[32]),
.OCL(jopfotomc[33]),
.OCM(jopfotomc[34]),
.OCN(jopfotomc[35]),
.OCO(jopfotomc[36]),
.OCP(jopfotomc[37]),
.OCQ(jopfotomc[38]),
.OCR(jopfotomc[39]),
.OCS(jopfotomc[40]),
.OCT(jopfotomc[41]),
.OCU(jopfotomc[42]),
.OCV(jopfotomc[43]),
.OCW(jopfotomc[44]),
.OCX(jopfotomc[45]),
.OCY(jopfotomc[46]),
.OCZ(jopfotomc[47]),
.ODA(lufotomd[0]),
.ODB(lufotomd[1]),
.ODC(lufotomd[2]),
.ODD(lufotomd[3]),
.ODE(lufotomd[4]),
.ODF(lufotomd[5]),
.ODG(lufotomd[6]),
.ODH(lufotomd[7]),
.ODI(lufotomd[8]),
.ODJ(lufotomd[9]),
.ODK(jopfotomd[32]),
.ODL(jopfotomd[33]),
.ODM(jopfotomd[34]),
.ODN(jopfotomd[35]),
.ODO(jopfotomd[36]),
.ODP(jopfotomd[37]),
.ODQ(jopfotomd[38]),
.ODR(jopfotomd[39]),
.ODS(jopfotomd[40]),
.ODT(jopfotomd[41]),
.ODU(jopfotomd[42]),
.ODV(jopfotomd[43]),
.ODW(jopfotomd[44]),
.ODX(jopfotomd[45]),
.ODY(jopfotomd[46]),
.ODZ(jopfotomd[47]),
.OEA(kopfotoma[32]),
.OEB(kopfotoma[33]),
.OEC(kopfotoma[34]),
.OED(kopfotoma[35]),
.OEE(kopfotoma[36]),
.OEF(kopfotoma[37]),
.OEG(kopfotoma[38]),
.OEH(kopfotoma[39]),
.OEI(kopfotoma[40]),
.OEJ(kopfotoma[41]),
.OEK(kopfotoma[42]),
.OEL(kopfotoma[43]),
.OEM(kopfotoma[44]),
.OEN(kopfotoma[45]),
.OEO(kopfotoma[46]),
.OEP(kopfotoma[47]),
.OFA(kopfotomb[32]),
.OFB(kopfotomb[33]),
.OFC(kopfotomb[34]),
.OFD(kopfotomb[35]),
.OFE(kopfotomb[36]),
.OFF(kopfotomb[37]),
.OFG(kopfotomb[38]),
.OFH(kopfotomb[39]),
.OFI(kopfotomb[40]),
.OFJ(kopfotomb[41]),
.OFK(kopfotomb[42]),
.OFL(kopfotomb[43]),
.OFM(kopfotomb[44]),
.OFN(kopfotomb[45]),
.OFO(kopfotomb[46]),
.OFP(kopfotomb[47]),
.OGA(kopfotomc[32]),
.OGB(kopfotomc[33]),
.OGC(kopfotomc[34]),
.OGD(kopfotomc[35]),
.OGE(kopfotomc[36]),
.OGF(kopfotomc[37]),
.OGG(kopfotomc[38]),
.OGH(kopfotomc[39]),
.OGI(kopfotomc[40]),
.OGJ(kopfotomc[41]),
.OGK(kopfotomc[42]),
.OGL(kopfotomc[43]),
.OGM(kopfotomc[44]),
.OGN(kopfotomc[45]),
.OGO(kopfotomc[46]),
.OGP(kopfotomc[47]),
.OHA(kopfotomd[32]),
.OHB(kopfotomd[33]),
.OHC(kopfotomd[34]),
.OHD(kopfotomd[35]),
.OHE(kopfotomd[36]),
.OHF(kopfotomd[37]),
.OHG(kopfotomd[38]),
.OHH(kopfotomd[39]),
.OHI(kopfotomd[40]),
.OHJ(kopfotomd[41]),
.OHK(kopfotomd[42]),
.OHL(kopfotomd[43]),
.OHM(kopfotomd[44]),
.OHN(kopfotomd[45]),
.OHO(kopfotomd[46]),
.OHP(kopfotomd[47]),
.OIA(mdludata[0]),
.OIB(mdludata[1]),
.OIC(mdludata[2]),
.OID(mdludata[3]),
.OIE(mdludata[4]),
.OIF(mdludata[5]),
.OIG(mdludata[6]),
.OIH(mdludata[7]),
.OII(mdludata[8]),
.OIJ(mdludata[9]),
.OIK(mdludata[10]),
.OIL(mdludata[11]),
.OIM(mdludata[12]),
.OJA(rafourtyeight),
.OKA(rarndbit[0]),
.OKB(rarndbit[1]),
.OKC(mchardrnd[0]),
.OKD(mchardrnd[1]),
.OKE(mchardrnd[2]),
.OKF(mchardrnd[3]),
.OKG(mchardrnd[4]),
.OLA(consoletonextra[0]),
.OLB(consoletonextra[1]),
.OLC(consoletonextra[2]),
.OLD(consoletonextra[3]),
.OLE(consoletonextra[4]),
.OLF(consoletonextra[5]),
.OLG(consoletonextra[6]),
.OLH(consoletonextra[7]),
.OLI(raloadbytenext),
.OMA(radeadstartnext),
.ONA(raparityerror));


tb tb0 (
.IAA(vrtocm[0]),
.IAB(vrtocm[1]),
.IAC(vrtocm[2]),
.IAD(vrtocm[3]),
.IAE(vrtocm[4]),
.IAF(vrtocm[5]),
.IAG(vrtocm[6]),
.IAH(vrtocm[7]),
.IAI(vrtocm[8]),
.IAJ(vrtocm[9]),
.IAK(vrtocm[10]),
.IAL(vrtocm[11]),
.IAM(vrtocm[12]),
.IAN(vrtocm[13]),
.IAO(vrtocm[14]),
.IAP(vrtocm[15]),
.IBA(vrtocm[16]),
.IBB(vrtocm[17]),
.IBC(vrtocm[18]),
.IBD(vrtocm[19]),
.IBE(vrtocm[20]),
.IBF(vrtocm[21]),
.IBG(vrtocm[22]),
.IBH(vrtocm[23]),
.IBI(vrtocm[24]),
.IBJ(vrtocm[25]),
.IBK(vrtocm[26]),
.IBL(vrtocm[27]),
.IBM(vrtocm[28]),
.IBN(vrtocm[29]),
.IBO(vrtocm[30]),
.IBP(vrtocm[31]),
.ICA(vrtocm[32]),
.ICB(vrtocm[33]),
.ICC(vrtocm[34]),
.ICD(vrtocm[35]),
.ICE(vrtocm[36]),
.ICF(vrtocm[37]),
.ICG(vrtocm[38]),
.ICH(vrtocm[39]),
.ICI(vrtocm[40]),
.ICJ(vrtocm[41]),
.ICK(vrtocm[42]),
.ICL(vrtocm[43]),
.ICM(vrtocm[44]),
.ICN(vrtocm[45]),
.ICO(vrtocm[46]),
.ICP(vrtocm[47]),
.IDA(vrtocm[48]),
.IDB(vrtocm[49]),
.IDC(vrtocm[50]),
.IDD(vrtocm[51]),
.IDE(vrtocm[52]),
.IDF(vrtocm[53]),
.IDG(vrtocm[54]),
.IDH(vrtocm[55]),
.IDI(vrtocm[56]),
.IDJ(vrtocm[57]),
.IDK(vrtocm[58]),
.IDL(vrtocm[59]),
.IDM(vrtocm[60]),
.IDN(vrtocm[61]),
.IDO(vrtocm[62]),
.IDP(vrtocm[63]),
.IEA(ebdatatb[0]),
.IEB(ebdatatb[1]),
.IEC(ebdatatb[2]),
.IED(ebdatatb[3]),
.IEE(ebdatatb[4]),
.IEF(ebdatatb[5]),
.IEG(ebdatatb[6]),
.IEH(ebdatatb[7]),
.IEI(ebdatatb[8]),
.IEJ(ebdatatb[9]),
.IEK(ebdatatb[10]),
.IEL(ebdatatb[11]),
.IEM(ebdatatb[12]),
.IEN(ebdatatb[13]),
.IEO(ebdatatb[14]),
.IEP(ebdatatb[15]),
.IFA(ebdatatb[16]),
.IFB(ebdatatb[17]),
.IFC(ebdatatb[18]),
.IFD(ebdatatb[19]),
.IFE(ebdatatb[20]),
.IFFF(ebdatatb[21]),
.IFG(ebdatatb[22]),
.IFH(ebdatatb[23]),
.IFI(ebdatatb[24]),
.IFJ(ebdatatb[25]),
.IFK(ebdatatb[26]),
.IFL(ebdatatb[27]),
.IFM(ebdatatb[28]),
.IFN(ebdatatb[29]),
.IFO(ebdatatb[30]),
.IFP(ebdatatb[31]),
.IGA(ebdatatb[32]),
.IGB(ebdatatb[33]),
.IGC(ebdatatb[34]),
.IGD(ebdatatb[35]),
.IGE(ebdatatb[36]),
.IGF(ebdatatb[37]),
.IGG(ebdatatb[38]),
.IGH(ebdatatb[39]),
.IGI(ebdatatb[40]),
.IGJ(ebdatatb[41]),
.IGK(ebdatatb[42]),
.IGL(ebdatatb[43]),
.IGM(ebdatatb[44]),
.IGN(ebdatatb[45]),
.IGO(ebdatatb[46]),
.IGP(ebdatatb[47]),
.IHA(ebdatatb[48]),
.IHB(ebdatatb[49]),
.IHC(ebdatatb[50]),
.IHD(ebdatatb[51]),
.IHE(ebdatatb[52]),
.IHF(ebdatatb[53]),
.IHG(ebdatatb[54]),
.IHH(ebdatatb[55]),
.IHI(ebdatatb[56]),
.IHJ(ebdatatb[57]),
.IHK(ebdatatb[58]),
.IHL(ebdatatb[59]),
.IHM(ebdatatb[60]),
.IHN(ebdatatb[61]),
.IHO(ebdatatb[62]),
.IHP(ebdatatb[63]),
.IIA(bp0mergetb1[0]),
.IIB(bp1mergetb1[0]),
.IIC(bp2mergetb1[0]),
.IID(bp3mergetb1[0]),
.IIE(bp0mergetb1[1]),
.IIF(bp1mergetb1[1]),
.IIG(bp2mergetb1[1]),
.IIH(bp3mergetb1[1]),
.III(bp0mergetb1[2]),
.IIJ(bp1mergetb1[2]),
.IIK(bp2mergetb1[2]),
.IIL(bp3mergetb1[2]),
.IIM(bp0mergetb1[3]),
.IIN(bp1mergetb1[3]),
.IIO(bp2mergetb1[3]),
.IIP(bp3mergetb1[3]),
.IIQ(bp0mergetb1[4]),
.IIR(bp1mergetb1[4]),
.IIS(bp2mergetb1[4]),
.IIT(bp3mergetb1[4]),
.IJA(ltwaystation[0]),
.IJB(ltwaystation[1]),
.IJC(ltwaystation[2]),
.IJD(ltwaystation[3]),
.IJE(ltwaystation[4]),
.IJF(ltwaystation[5]),
.IJG(ltwaystation[6]),
.IJH(ltwaystation[7]),
.IJI(ltwaystation[8]),
.IJJ(ltwaystation[9]),
.IJK(ltwaystation[10]),
.IJL(ltwaystation[11]),
.IJM(ltwaystation[12]),
.IJN(ltwaystation[13]),
.IJO(ltwaystation[14]),
.IJP(ltwaystation[15]),
.IKA(gosdatatotb),
.IKB(selextdata),
.IKC(recyclebd),
//.IKD(pkgphasetb),
.IKD(phasejbtotm[1]),
.IZZ (sysclock),
.OAA(p0pktdata[0]),
.OAB(p0pktdata[1]),
.OAC(p0pktdata[2]),
.OAD(p0pktdata[3]),
.OAE(p0pktdata[4]),
.OAF(p0pktdata[5]),
.OAG(p0pktdata[6]),
.OAH(p0pktdata[7]),
.OAI(p0pktdata[8]),
.OAJ(p0pktdata[9]),
.OAK(p0pktdata[10]),
.OAL(p0pktdata[11]),
.OAM(p0pktdata[12]),
.OAN(p0pktdata[13]),
.OAO(p0pktdata[14]),
.OAP(p0pktdata[15]),
.OAQ(p0pktdata[16]),
.OAR(p0pktdata[17]),
.OAS(p0pktdata[18]),
.OAT(p0pktdata[19]),
.OAU(p0pktdata[20]),
.OAV(p0pktdata[21]),
.OAW(p0pktdata[22]),
.OAX(p0pktdata[23]),
.OBA(p1pktdata[0]),
.OBB(p1pktdata[1]),
.OBC(p1pktdata[2]),
.OBD(p1pktdata[3]),
.OBE(p1pktdata[4]),
.OBF(p1pktdata[5]),
.OBG(p1pktdata[6]),
.OBH(p1pktdata[7]),
.OBI(p1pktdata[8]),
.OBJ(p1pktdata[9]),
.OBK(p1pktdata[10]),
.OBL(p1pktdata[11]),
.OBM(p1pktdata[12]),
.OBN(p1pktdata[13]),
.OBO(p1pktdata[14]),
.OBP(p1pktdata[15]),
.OBQ(p1pktdata[16]),
.OBR(p1pktdata[17]),
.OBS(p1pktdata[18]),
.OBT(p1pktdata[19]),
.OBU(p1pktdata[20]),
.OBV(p1pktdata[21]),
.OBW(p1pktdata[22]),
.OBX(p1pktdata[23]),
.OCA(p2pktdata[0]),
.OCB(p2pktdata[1]),
.OCC(p2pktdata[2]),
.OCD(p2pktdata[3]),
.OCE(p2pktdata[4]),
.OCF(p2pktdata[5]),
.OCG(p2pktdata[6]),
.OCH(p2pktdata[7]),
.OCI(p2pktdata[8]),
.OCJ(p2pktdata[9]),
.OCK(p2pktdata[10]),
.OCL(p2pktdata[11]),
.OCM(p2pktdata[12]),
.OCN(p2pktdata[13]),
.OCO(p2pktdata[14]),
.OCP(p2pktdata[15]),
.OCQ(p2pktdata[16]),
.OCR(p2pktdata[17]),
.OCS(p2pktdata[18]),
.OCT(p2pktdata[19]),
.OCU(p2pktdata[20]),
.OCV(p2pktdata[21]),
.OCW(p2pktdata[22]),
.OCX(p2pktdata[23]),
.ODA(p3pktdata[0]),
.ODB(p3pktdata[1]),
.ODC(p3pktdata[2]),
.ODD(p3pktdata[3]),
.ODE(p3pktdata[4]),
.ODF(p3pktdata[5]),
.ODG(p3pktdata[6]),
.ODH(p3pktdata[7]),
.ODI(p3pktdata[8]),
.ODJ(p3pktdata[9]),
.ODK(p3pktdata[10]),
.ODL(p3pktdata[11]),
.ODM(p3pktdata[12]),
.ODN(p3pktdata[13]),
.ODO(p3pktdata[14]),
.ODP(p3pktdata[15]),
.ODQ(p3pktdata[16]),
.ODR(p3pktdata[17]),
.ODS(p3pktdata[18]),
.ODT(p3pktdata[19]),
.ODU(p3pktdata[20]),
.ODV(p3pktdata[21]),
.ODW(p3pktdata[22]),
.ODX(p3pktdata[23]),
.OFA(bankptrtoqb[0]),
.OFB(bankptrtoqb[1]),
.OFC(bankptrtoqb[2]),
.OFD(bankptrtoqb[3]),
.OFE(bankptrtoqb[4])
);


tc tc0 (
.IAA(p0pktdata[0]),
.IAB(p0pktdata[1]),
.IAC(p0pktdata[2]),
.IAD(p0pktdata[3]),
.IAE(p0pktdata[4]),
.IAF(p0pktdata[5]),
.IAG(p0pktdata[6]),
.IAH(p0pktdata[7]),
.IAI(p0pktdata[8]),
.IAJ(p0pktdata[9]),
.IAK(p0pktdata[10]),
.IAL(p0pktdata[11]),
.IAM(p0pktdata[12]),
.IAN(p0pktdata[13]),
.IAO(p0pktdata[14]),
.IAP(p0pktdata[15]),
.IAQ(p0pktdata[16]),
.IAR(p0pktdata[17]),
.IAS(p0pktdata[18]),
.IAT(p0pktdata[19]),
.IAU(p0pktdata[20]),
.IAV(p0pktdata[21]),
.IAW(p0pktdata[22]),
.IAX(p0pktdata[23]),
.IBA(p1pktdata[0]),
.IBB(p1pktdata[1]),
.IBC(p1pktdata[2]),
.IBD(p1pktdata[3]),
.IBE(p1pktdata[4]),
.IBF(p1pktdata[5]),
.IBG(p1pktdata[6]),
.IBH(p1pktdata[7]),
.IBI(p1pktdata[8]),
.IBJ(p1pktdata[9]),
.IBK(p1pktdata[10]),
.IBL(p1pktdata[11]),
.IBM(p1pktdata[12]),
.IBN(p1pktdata[13]),
.IBO(p1pktdata[14]),
.IBP(p1pktdata[15]),
.IBQ(p1pktdata[16]),
.IBR(p1pktdata[17]),
.IBS(p1pktdata[18]),
.IBT(p1pktdata[19]),
.IBU(p1pktdata[20]),
.IBV(p1pktdata[21]),
.IBW(p1pktdata[22]),
.IBX(p1pktdata[23]),
.ICA(p2pktdata[0]),
.ICB(p2pktdata[1]),
.ICC(p2pktdata[2]),
.ICD(p2pktdata[3]),
.ICE(p2pktdata[4]),
.ICF(p2pktdata[5]),
.ICG(p2pktdata[6]),
.ICH(p2pktdata[7]),
.ICI(p2pktdata[8]),
.ICJ(p2pktdata[9]),
.ICK(p2pktdata[10]),
.ICL(p2pktdata[11]),
.ICM(p2pktdata[12]),
.ICN(p2pktdata[13]),
.ICO(p2pktdata[14]),
.ICP(p2pktdata[15]),
.ICQ(p2pktdata[16]),
.ICR(p2pktdata[17]),
.ICS(p2pktdata[18]),
.ICT(p2pktdata[19]),
.ICU(p2pktdata[20]),
.ICV(p2pktdata[21]),
.ICW(p2pktdata[22]),
.ICX(p2pktdata[23]),
.IDA(p3pktdata[0]),
.IDB(p3pktdata[1]),
.IDC(p3pktdata[2]),
.IDD(p3pktdata[3]),
.IDE(p3pktdata[4]),
.IDF(p3pktdata[5]),
.IDG(p3pktdata[6]),
.IDH(p3pktdata[7]),
.IDI(p3pktdata[8]),
.IDJ(p3pktdata[9]),
.IDK(p3pktdata[10]),
.IDL(p3pktdata[11]),
.IDM(p3pktdata[12]),
.IDN(p3pktdata[13]),
.IDO(p3pktdata[14]),
.IDP(p3pktdata[15]),
.IDQ(p3pktdata[16]),
.IDR(p3pktdata[17]),
.IDS(p3pktdata[18]),
.IDT(p3pktdata[19]),
.IDU(p3pktdata[20]),
.IDV(p3pktdata[21]),
.IDW(p3pktdata[22]),
.IDX(p3pktdata[23]),
.IEA(addrtotc[0]),
.IEB(addrtotc[1]),
.IEC(addrtotc[2]),
.IED(addrtotc[3]),
.IEE(addrtotc[4]),
.IEF(addrtotc[5]),
.IEG(addrtotc[6]),
.IEH(addrtotc[7]),
.IEI(addrtotc[8]),
.IEJ(addrtotc[9]),
.IEK(addrtotc[10]),
.IEL(addrtotc[11]),
.IEM(addrtotc[12]),
.IEN(addrtotc[13]),
.IEO(addrtotc[14]),
.IEP(addrtotc[15]),
.IEQ(addrtotc[16]),
.IER(addrtotc[17]),
.IES(addrtotc[18]),
.IET(addrtotc[19]),
.IEU(addrtotc[20]),
.IEV(addrtotc[21]),
.IEW(addrtotc[22]),
.IEX(addrtotc[23]),
.IFA(goquadrant[0]),
.IFB(goquadrant[1]),
.IFC(goquadrant[2]),
.IFD(goquadrant[3]),
.IGA(qd0release[0]),
.IGB(qd0release[1]),
.IGC(qd1release[0]),
.IGD(qd1release[1]),
.IGE(qd2release[0]),
.IGF(qd2release[1]),
.IGG(qd3release[0]),
.IGH(qd3release[1]),
.IHA(phasejbtotm[2]),
.IHC(deadstartfromea),
.IHD(backupfromtf),
.IZZ (sysclock),
.OAA(quad0packet[0]),
.OAB(quad0packet[1]),
.OAC(quad0packet[2]),
.OAD(quad0packet[3]),
.OAE(quad0packet[4]),
.OAF(quad0packet[5]),
.OAG(quad0packet[6]),
.OAH(quad0packet[7]),
.OAI(quad0packet[8]),
.OAJ(quad0packet[9]),
.OAK(quad0packet[10]),
.OAL(quad0packet[11]),
.OAM(quad0packet[12]),
.OAN(quad0packet[13]),
.OAO(quad0packet[14]),
.OAP(quad0packet[15]),
.OAQ(quad0packet[16]),
.OAR(quad0packet[17]),
.OAS(quad0packet[18]),
.OAT(quad0packet[19]),
.OAU(quad0packet[20]),
.OAV(quad0packet[21]),
.OAW(quad0packet[22]),
.OAX(quad0packet[23]),
.OBA(quad1packet[0]),
.OBB(quad1packet[1]),
.OBC(quad1packet[2]),
.OBD(quad1packet[3]),
.OBE(quad1packet[4]),
.OBF(quad1packet[5]),
.OBG(quad1packet[6]),
.OBH(quad1packet[7]),
.OBI(quad1packet[8]),
.OBJ(quad1packet[9]),
.OBK(quad1packet[10]),
.OBL(quad1packet[11]),
.OBM(quad1packet[12]),
.OBN(quad1packet[13]),
.OBO(quad1packet[14]),
.OBP(quad1packet[15]),
.OBQ(quad1packet[16]),
.OBR(quad1packet[17]),
.OBS(quad1packet[18]),
.OBT(quad1packet[19]),
.OBU(quad1packet[20]),
.OBV(quad1packet[21]),
.OBW(quad1packet[22]),
.OBX(quad1packet[23]),
.OCA(quad2packet[0]),
.OCB(quad2packet[1]),
.OCC(quad2packet[2]),
.OCD(quad2packet[3]),
.OCE(quad2packet[4]),
.OCF(quad2packet[5]),
.OCG(quad2packet[6]),
.OCH(quad2packet[7]),
.OCI(quad2packet[8]),
.OCJ(quad2packet[9]),
.OCK(quad2packet[10]),
.OCL(quad2packet[11]),
.OCM(quad2packet[12]),
.OCN(quad2packet[13]),
.OCO(quad2packet[14]),
.OCP(quad2packet[15]),
.OCQ(quad2packet[16]),
.OCR(quad2packet[17]),
.OCS(quad2packet[18]),
.OCT(quad2packet[19]),
.OCU(quad2packet[20]),
.OCV(quad2packet[21]),
.OCW(quad2packet[22]),
.OCX(quad2packet[23]),
.ODA(quad3packet[0]),
.ODB(quad3packet[1]),
.ODC(quad3packet[2]),
.ODD(quad3packet[3]),
.ODE(quad3packet[4]),
.ODF(quad3packet[5]),
.ODG(quad3packet[6]),
.ODH(quad3packet[7]),
.ODI(quad3packet[8]),
.ODJ(quad3packet[9]),
.ODK(quad3packet[10]),
.ODL(quad3packet[11]),
.ODM(quad3packet[12]),
.ODN(quad3packet[13]),
.ODO(quad3packet[14]),
.ODP(quad3packet[15]),
.ODQ(quad3packet[16]),
.ODR(quad3packet[17]),
.ODS(quad3packet[18]),
.ODT(quad3packet[19]),
.ODU(quad3packet[20]),
.ODV(quad3packet[21]),
.ODW(quad3packet[22]),
.ODX(quad3packet[23]));



  
td td0( 
.IAA(quad0memparcel[0]),
.IAB(quad0memparcel[1]),
.IAC(quad0memparcel[2]),
.IAD(quad0memparcel[3]),
.IAE(quad0memparcel[4]),
.IAF(quad0memparcel[5]),
.IAG(quad0memparcel[6]),
.IAH(quad0memparcel[7]),
.IAI(quad0memparcel[8]),
.IAJ(quad0memparcel[9]),
.IAK(quad0memparcel[10]),
.IAL(quad0memparcel[11]),
.IAM(quad0memparcel[12]),
.IAN(quad0memparcel[13]),
.IAO(quad0memparcel[14]),
.IAP(quad0memparcel[15]),
.IAQ(quad0memparcel[16]),
.IAR(quad0memparcel[17]),
.IAS(quad0memparcel[18]),
.IAT(quad0memparcel[19]),
.IAU(quad0memparcel[20]),
.IAV(quad0memparcel[21]),
.IAW(quad0memparcel[22]),
.IAX(quad0memparcel[23]),
.IBA(quad1memparcel[0]),
.IBB(quad1memparcel[1]),
.IBC(quad1memparcel[2]),
.IBD(quad1memparcel[3]),
.IBE(quad1memparcel[4]),
.IBF(quad1memparcel[5]),
.IBG(quad1memparcel[6]),
.IBH(quad1memparcel[7]),
.IBI(quad1memparcel[8]),
.IBJ(quad1memparcel[9]),
.IBK(quad1memparcel[10]),
.IBL(quad1memparcel[11]),
.IBM(quad1memparcel[12]),
.IBN(quad1memparcel[13]),
.IBO(quad1memparcel[14]),
.IBP(quad1memparcel[15]),
.IBQ(quad1memparcel[16]),
.IBR(quad1memparcel[17]),
.IBS(quad1memparcel[18]),
.IBT(quad1memparcel[19]),
.IBU(quad1memparcel[20]),
.IBV(quad1memparcel[21]),
.IBW(quad1memparcel[22]),
.IBX(quad1memparcel[23]),
.ICA(quad2memparcel[0]),
.ICB(quad2memparcel[1]),
.ICC(quad2memparcel[2]),
.ICD(quad2memparcel[3]),
.ICE(quad2memparcel[4]),
.ICF(quad2memparcel[5]),
.ICG(quad2memparcel[6]),
.ICH(quad2memparcel[7]),
.ICI(quad2memparcel[8]),
.ICJ(quad2memparcel[9]),
.ICK(quad2memparcel[10]),
.ICL(quad2memparcel[11]),
.ICM(quad2memparcel[12]),
.ICN(quad2memparcel[13]),
.ICO(quad2memparcel[14]),
.ICP(quad2memparcel[15]),
.ICQ(quad2memparcel[16]),
.ICR(quad2memparcel[17]),
.ICS(quad2memparcel[18]),
.ICT(quad2memparcel[19]),
.ICU(quad2memparcel[20]),
.ICV(quad2memparcel[21]),
.ICW(quad2memparcel[22]),
.ICX(quad2memparcel[23]),
.IDA(quad1memparcel[0]),
.IDB(quad1memparcel[1]),
.IDC(quad1memparcel[2]),
.IDD(quad1memparcel[3]),
.IDE(quad1memparcel[4]),
.IDF(quad1memparcel[5]),
.IDG(quad1memparcel[6]),
.IDH(quad1memparcel[7]),
.IDI(quad1memparcel[8]),
.IDJ(quad1memparcel[9]),
.IDK(quad1memparcel[10]),
.IDL(quad1memparcel[11]),
.IDM(quad1memparcel[12]),
.IDN(quad1memparcel[13]),
.IDO(quad1memparcel[14]),
.IDP(quad1memparcel[15]),
.IDQ(quad1memparcel[16]),
.IDR(quad1memparcel[17]),
.IDS(quad1memparcel[18]),
.IDT(quad1memparcel[19]),
.IDU(quad1memparcel[20]),
.IDV(quad1memparcel[21]),
.IDW(quad1memparcel[22]),
.IDX(quad1memparcel[23]),
.IEA(quad0memdest[0]),
.IEB(quad0memdest[1]),
.IEC(quad0memdest[2]),
.IED(quad0memdest[3]),
.IEE(quad0memdest[4]),
.IEF(quad0memdest[5]),
.IFA(quad1memdest[0]),
.IFB(quad1memdest[1]),
.IFC(quad1memdest[2]),
.IFD(quad1memdest[3]),
.IFE(quad1memdest[4]),
.IFFF(quad1memdest[5]),
.IGA(quad2memdest[0]),
.IGB(quad2memdest[1]),
.IGC(quad2memdest[2]),
.IGD(quad2memdest[3]),
.IGE(quad2memdest[4]),
.IGF(quad2memdest[5]),
.IHA(quad3memdest[0]),
.IHB(quad3memdest[1]),
.IHC(quad3memdest[2]),
.IHD(quad3memdest[3]),
.IHE(quad3memdest[4]),
.IHF(quad3memdest[5]),
.IIA(phasetotd),
.IJA(enablesecded),
.IZZ (sysclock),
.OAA(commemtoie[0]),
.OAB(commemtoie[1]),
.OAC(commemtoie[2]),
.OAD(commemtoie[3]),
.OAE(commemtoie[4]),
.OAF(commemtoie[5]),
.OAG(commemtoie[6]),
.OAH(commemtoie[7]),
.OAI(commemtoie[8]),
.OAJ(commemtoie[9]),
.OAK(commemtoie[10]),
.OAL(commemtoie[11]),
.OAM(commemtoie[12]),
.OAN(commemtoie[13]),
.OAO(commemtoie[14]),
.OAP(commemtoie[15]),
.OBA(commemtoie[16]),
.OBB(commemtoie[17]),
.OBC(commemtoie[18]),
.OBD(commemtoie[19]),
.OBE(commemtoie[20]),
.OBF(commemtoie[21]),
.OBG(commemtoie[22]),
.OBH(commemtoie[23]),
.OBI(commemtoie[24]),
.OBJ(commemtoie[25]),
.OBK(commemtoie[26]),
.OBL(commemtoie[27]),
.OBM(commemtoie[28]),
.OBN(commemtoie[29]),
.OBO(commemtoie[30]),
.OBP(commemtoie[31]),
.OCA(commemtoie[32]),
.OCB(commemtoie[33]),
.OCC(commemtoie[34]),
.OCD(commemtoie[35]),
.OCE(commemtoie[36]),
.OCF(commemtoie[37]),
.OCG(commemtoie[38]),
.OCH(commemtoie[39]),
.OCI(commemtoie[40]),
.OCJ(commemtoie[41]),
.OCK(commemtoie[42]),
.OCL(commemtoie[43]),
.OCM(commemtoie[44]),
.OCN(commemtoie[45]),
.OCO(commemtoie[46]),
.OCP(commemtoie[47]),
.ODA(commemtoie[48]),
.ODB(commemtoie[49]),
.ODC(commemtoie[50]),
.ODD(commemtoie[51]),
.ODE(commemtoie[52]),
.ODF(commemtoie[53]),
.ODG(commemtoie[54]),
.ODH(commemtoie[55]),
.ODI(commemtoie[56]),
.ODJ(commemtoie[57]),
.ODK(commemtoie[58]),
.ODL(commemtoie[59]),
.ODM(commemtoie[60]),
.ODN(commemtoie[61]),
.ODO(commemtoie[62]),
.ODP(commemtoie[63]),
.OEA(commemtovr[0]),
.OEB(commemtovr[1]),
.OEC(commemtovr[2]),
.OED(commemtovr[3]),
.OEE(commemtovr[4]),
.OEF(commemtovr[5]),
.OEG(commemtovr[6]),
.OEH(commemtovr[7]),
.OEI(commemtovr[8]),
.OEJ(commemtovr[9]),
.OEK(commemtovr[10]),
.OEL(commemtovr[11]),
.OEM(commemtovr[12]),
.OEN(commemtovr[13]),
.OEO(commemtovr[14]),
.OEP(commemtovr[15]),
.OFA(commemtovr[16]),
.OFB(commemtovr[17]),
.OFC(commemtovr[18]),
.OFD(commemtovr[19]),
.OFE(commemtovr[20]),
.OFF(commemtovr[21]),
.OFG(commemtovr[22]),
.OFH(commemtovr[23]),
.OFI(commemtovr[24]),
.OFJ(commemtovr[25]),
.OFK(commemtovr[26]),
.OFL(commemtovr[27]),
.OFM(commemtovr[28]),
.OFN(commemtovr[29]),
.OFO(commemtovr[30]),
.OFP(commemtovr[31]),
.OGA(commemtovr[32]),
.OGB(commemtovr[33]),
.OGC(commemtovr[34]),
.OGD(commemtovr[35]),
.OGE(commemtovr[36]),
.OGF(commemtovr[37]),
.OGG(commemtovr[38]),
.OGH(commemtovr[39]),
.OGI(commemtovr[40]),
.OGJ(commemtovr[41]),
.OGK(commemtovr[42]),
.OGL(commemtovr[43]),
.OGM(commemtovr[44]),
.OGN(commemtovr[45]),
.OGO(commemtovr[46]),
.OGP(commemtovr[47]),
.OHA(commemtovr[48]),
.OHB(commemtovr[49]),
.OHC(commemtovr[50]),
.OHD(commemtovr[51]),
.OHE(commemtovr[52]),
.OHF(commemtovr[53]),
.OHG(commemtovr[54]),
.OHH(commemtovr[55]),
.OHI(commemtovr[56]),
.OHJ(commemtovr[57]),
.OHK(commemtovr[58]),
.OHL(commemtovr[59]),
.OHM(commemtovr[60]),
.OHN(commemtovr[61]),
.OHO(commemtovr[62]),
.OHP(commemtovr[63]),
.OIA(syndrome[0]),
.OIB(syndrome[1]),
.OIC(syndrome[2]),
.OID(syndrome[3]),
.OIE(syndrome[4]),
.OIF(syndrome[5]),
.OIG(syndrome[6]),
.OIH(syndrome[7]),
.OJA(singlebiterror),
.OKA(memarivtojc0[0]),
.OKB(memarivtojc0[1]),
.OKC(memarivtojc0[2]),
.OKD(memarivtojc0[3]),
.OKE(memarivtojc0[4]),
.OLA(memarivtojc1[0]),
.OLB(memarivtojc1[1]),
.OLC(memarivtojc1[2]),
.OLD(memarivtojc1[3]),
.OLE(memarivtojc1[4]),
.OMA(memdestja[0]),
.OMB(memdestja[1]),
.OMC(memdestja[2]),
.OMD(memdestja[3]),
.ONA(fetcharrival[0]),
.ONB(fetcharrival[1]),
.ONC(fetcharrival[2]),
.OOA(fetcharrivaltoeb[0]),
.OOB(fetcharrivaltoeb[1]),
.OOC(fetcharrivaltoeb[2]),
.OPA(readparity));



tf tf0 ( 
.IAA(araddrtotf[0]),
.IAB(araddrtotf[1]),
.IAC(araddrtotf[2]),
.IAD(araddrtotf[3]),
.IAE(araddrtotf[4]),
.IAF(araddrtotf[5]),
.IAG(araddrtotf[6]),
.IAH(araddrtotf[7]),
.IAI(araddrtotf[8]),
.IAJ(araddrtotf[9]),
.IAK(araddrtotf[10]),
.IAL(araddrtotf[11]),
.IAM(araddrtotf[12]),
.IAN(araddrtotf[13]),
.IAO(araddrtotf[14]),
.IAP(araddrtotf[15]),
.IBA(araddrtotf[16]),
.IBB(araddrtotf[17]),
.IBC(araddrtotf[18]),
.IBD(araddrtotf[19]),
.IBE(araddrtotf[20]),
.IBF(araddrtotf[21]),
.IBG(araddrtotf[22]),
.IBH(araddrtotf[23]),
.IBI(araddrtotf[24]),
.IBJ(araddrtotf[25]),
.IBK(araddrtotf[26]),
.IBL(araddrtotf[27]),
.IBM(araddrtotf[28]),
.IBN(araddrtotf[29]),
.IBO(araddrtotf[30]),
.IBP(araddrtotf[31]),
.ICA(ebaddrtotf[0]),
.ICB(ebaddrtotf[1]),
.ICC(ebaddrtotf[2]),
.ICD(ebaddrtotf[3]),
.ICE(ebaddrtotf[4]),
.ICF(ebaddrtotf[5]),
.ICG(ebaddrtotf[6]),
.ICH(ebaddrtotf[7]),
.ICI(ebaddrtotf[8]),
.ICJ(ebaddrtotf[9]),
.ICK(ebaddrtotf[10]),
.ICL(ebaddrtotf[11]),
.ICM(ebaddrtotf[12]),
.ICN(ebaddrtotf[13]),
.ICO(ebaddrtotf[14]),
.ICP(ebaddrtotf[15]),
.IDA(ebaddrtotf[16]),
.IDB(ebaddrtotf[17]),
.IDC(ebaddrtotf[18]),
.IDD(ebaddrtotf[19]),
.IDE(ebaddrtotf[20]),
.IDF(ebaddrtotf[21]),
.IDG(ebaddrtotf[22]),
.IDH(ebaddrtotf[23]),
.IDI(ebaddrtotf[24]),
.IDJ(ebaddrtotf[25]),
.IDK(ebaddrtotf[26]),
.IDL(ebaddrtotf[27]),
.IDM(ebaddrtotf[28]),
.IDN(ebaddrtotf[29]),
.IDO(ebaddrtotf[30]),
.IDP(ebaddrtotf[31]),
//.IEA(ifaddrtotf[0]),
//.IEB(ifaddrtotf[1]),
//.IEC(ifaddrtotf[2]),
//.IED(ifaddrtotf[3]),
//.IEE(ifaddrtotf[4]),
//.IEF(ifaddrtotf[5]),
//.IEG(ifaddrtotf[6]),
//.IEH(ifaddrtotf[7]),
//.IEI(ifaddrtotf[8]),
//.IEJ(ifaddrtotf[9]),
//.IEK(ifaddrtotf[10]),
//.IEL(ifaddrtotf[11]),
//.IEM(ifaddrtotf[12]),
//.IEN(ifaddrtotf[13]),
//.IEO(ifaddrtotf[14]),
//.IEP(ifaddrtotf[15]),
//.IFA(ifaddrtotf[16]),
//.IFB(ifaddrtotf[17]),
//.IFC(ifaddrtotf[18]),
//.IFD(ifaddrtotf[19]),
//.IFE(ifaddrtotf[20]),
//.IFFF(ifaddrtotf[21]),
//.IFG(ifaddrtotf[22]),
//.IFH(ifaddrtotf[23]),
//.IFI(ifaddrtotf[24]),
//.IFJ(ifaddrtotf[25]),
//.IFK(ifaddrtotf[26]),
//.IFL(ifaddrtotf[27]),
//.IFM(ifaddrtotf[28]),
//.IFN(ifaddrtotf[29]),
//.IFO(ifaddrtotf[30]),
//.IFP(ifaddrtotf[31]),
.IEA(tfbaseaddr[0]),
.IEB(tfbaseaddr[1]),
.IEC(tfbaseaddr[2]),
.IED(tfbaseaddr[3]),
.IEE(tfbaseaddr[4]),
.IEF(tfbaseaddr[5]),
.IEG(tfbaseaddr[6]),
.IEH(tfbaseaddr[7]),
.IEI(tfbaseaddr[8]),
.IEJ(tfbaseaddr[9]),
.IEK(tfbaseaddr[10]),
.IEL(tfbaseaddr[11]),
.IEM(tfbaseaddr[12]),
.IEN(tfbaseaddr[13]),
.IEO(tfbaseaddr[14]),
.IEP(tfbaseaddr[15]),
.IFA(tfbaseaddr[16]),
.IFB(tfbaseaddr[17]),
.IFC(tfbaseaddr[18]),
.IFD(tfbaseaddr[19]),
.IFE(tfbaseaddr[20]),
.IFFF(tfbaseaddr[21]),
.IFG(tfbaseaddr[22]),
.IFH(tfbaseaddr[23]),
.IFI(tfbaseaddr[24]),
.IFJ(tfbaseaddr[25]),
.IFK(tfbaseaddr[26]),
.IFL(tfbaseaddr[27]),
.IFM(tfbaseaddr[28]),
.IFN(tfbaseaddr[29]),
.IFO(tfbaseaddr[30]),
.IFP(tfbaseaddr[31]),
.IGA(vraddrtotf[0]),
.IGB(vraddrtotf[1]),
.IGC(vraddrtotf[2]),
.IGD(vraddrtotf[3]),
.IGE(vraddrtotf[4]),
.IGF(vraddrtotf[5]),
.IGG(vraddrtotf[6]),
.IGH(vraddrtotf[7]),
.IGI(vraddrtotf[8]),
.IGJ(vraddrtotf[9]),
.IGK(vraddrtotf[10]),
.IGL(vraddrtotf[11]),
.IGM(vraddrtotf[12]),
.IGN(vraddrtotf[13]),
.IGO(vraddrtotf[14]),
.IGP(vraddrtotf[15]),
.IHA(vraddrtotf[16]),
.IHB(vraddrtotf[17]),
.IHC(vraddrtotf[18]),
.IHD(vraddrtotf[19]),
.IHE(vraddrtotf[20]),
.IHF(vraddrtotf[21]),
.IHG(vraddrtotf[22]),
.IHH(vraddrtotf[23]),
.IHI(vraddrtotf[24]),
.IHJ(vraddrtotf[25]),
.IHK(vraddrtotf[26]),
.IHL(vraddrtotf[27]),
.IHM(vraddrtotf[28]),
.IHN(vraddrtotf[29]),
.IHO(vraddrtotf[30]),
.IHP(vraddrtotf[31]),
.IIA(memdestcode[0]),
.IIB(memdestcode[1]),
.IIC(memdestcode[2]),
.IID(memdestcode[3]),
.IIE(memdestcode[4]),
.IIF(memdestcode[5]),
.IJA(qb0quadrela[0]),
.IJB(qb0quadrela[1]),
.IJC(qb1quadrela[0]),
.IJD(qb1quadrela[1]),
.IJE(qb2quadrela[0]),
.IJF(qb2quadrela[1]),
.IJG(qb3quadrela[0]),
.IJH(qb3quadrela[1]),
.IKA(validaddtotf),
.IKB(reproshtdata),
.IKC(enablecmrangetotf),
.IKD(gathertest),
.IKE(phasejbtotm[0]),
.IKF(incrtofirst),
.IKG(artofirstadder),
.IKH(looptofirstaddr),
.IKI(holdtofirstaddr),
.IKJ(vrtosecondadder),
.IKK(carrietosecondaddr),
.IKM(holdtosecondaddr),
.IKN(ioaddrtothirdaddr),
.IKO(incrtothirdaddr),
.IKP(basetothirdaddr),
.IKQ(ardatatoincr),
.IKR(ifinincrement),
.IKS(holdinincrement),
//.IKT(enterbasetf),
.IKT(setbaseaddr),
.IKU(enterlimittf),
.ILA(refreshtotf),
.IZZ (sysclock),
.OAA(packreqq0[0]),
.OAB(packreqq0[1]),
.OAC(packreqq0[2]),
.OAD(packreqq0[3]),
.OAE(packreqq0[4]),
.OAF(packreqq0[5]),
.OAG(packreqq0[6]),
.OAH(packreqq0[7]),
.OAI(packreqq0[8]),
.OAJ(packreqq0[9]),
.OAK(packreqq0[10]),
.OAL(packreqq0[11]),
.OAM(packreqq0[12]),
.OAN(packreqq0[13]),
.OBA(packreqq1[0]),
.OBB(packreqq1[1]),
.OBC(packreqq1[2]),
.OBD(packreqq1[3]),
.OBE(packreqq1[4]),
.OBF(packreqq1[5]),
.OBG(packreqq1[6]),
.OBH(packreqq1[7]),
.OBI(packreqq1[8]),
.OBJ(packreqq1[9]),
.OBK(packreqq1[10]),
.OBL(packreqq1[11]),
.OBM(packreqq1[12]),
.OBN(packreqq1[13]),
.OCA(packreqq2[0]),
.OCB(packreqq2[1]),
.OCC(packreqq2[2]),
.OCD(packreqq2[3]),
.OCE(packreqq2[4]),
.OCF(packreqq2[5]),
.OCG(packreqq2[6]),
.OCH(packreqq2[7]),
.OCI(packreqq2[8]),
.OCJ(packreqq2[9]),
.OCK(packreqq2[10]),
.OCL(packreqq2[11]),
.OCM(packreqq2[12]),
.OCN(packreqq2[13]),
.ODA(packreqq3[0]),
.ODB(packreqq3[1]),
.ODC(packreqq3[2]),
.ODD(packreqq3[3]),
.ODE(packreqq3[4]),
.ODF(packreqq3[5]),
.ODG(packreqq3[6]),
.ODH(packreqq3[7]),
.ODI(packreqq3[8]),
.ODJ(packreqq3[9]),
.ODK(packreqq3[10]),
.ODL(packreqq3[11]),
.ODM(packreqq3[12]),
.ODN(packreqq3[13]),
.OEA(addrtotc[0]),
.OEB(addrtotc[1]),
.OEC(addrtotc[2]),
.OED(addrtotc[3]),
.OEE(addrtotc[4]),
.OEF(addrtotc[5]),
.OEG(addrtotc[6]),
.OEH(addrtotc[7]),
.OEI(addrtotc[8]),
.OEJ(addrtotc[9]),
.OEK(addrtotc[10]),
.OEL(addrtotc[11]),
.OEM(addrtotc[12]),
.OEN(addrtotc[13]),
.OEO(addrtotc[14]),
.OEP(addrtotc[15]),
.OEQ(addrtotc[16]),
.OER(addrtotc[17]),
.OES(addrtotc[18]),
.OET(addrtotc[19]),
.OEU(addrtotc[20]),
.OEV(addrtotc[21]),
.OEW(addrtotc[22]),
.OEX(addrtotc[23]),
.OFA(goquadrant[0]),
.OFB(goquadrant[1]),
.OFC(goquadrant[2]),
.OFD(goquadrant[3]),
.OHA(backupcnd[0]),
.OHB(backupcnd[1]),
.OHC(backupcnd[2]),
.OHD(backupcnd[3]),
.OHE(backupcnd[4]),
.OIA(tfflagtolights[0]),
.OIB(tfflagtolights[1]),
.OIC(tfflagtolights[2]),
.OID(tfflagtolights[3]),
.OIE(tfflagtolights[4]),
.OIF(tfflagtolights[5]),
.OIG(tfflagtolights[6]),
.OIH(tfflagtolights[7]),
.OKA(cmrangeerrortoea),
.OLA(bufferdataqd0),
.OLB(bufferdataqd1),
.OLC(bufferdataqd2),
.OLD(bufferdataqd3));


 
va va0 (
.IAA(vrtovaj[0]),
.IAB(vrtovaj[1]),
.IAC(vrtovaj[2]),
.IAD(vrtovaj[3]),
.IAE(vrtovaj[4]),
.IAF(vrtovaj[5]),
.IAG(vrtovaj[6]),
.IAH(vrtovaj[7]),
.IAI(vrtovaj[8]),
.IAJ(vrtovaj[9]),
.IAK(vrtovaj[10]),
.IAL(vrtovaj[11]),
.IAM(vrtovaj[12]),
.IAN(vrtovaj[13]),
.IAO(vrtovaj[14]),
.IAP(vrtovaj[15]),
.IBA(vrtovaj[16]),
.IBB(vrtovaj[17]),
.IBC(vrtovaj[18]),
.IBD(vrtovaj[19]),
.IBE(vrtovaj[20]),
.IBF(vrtovaj[21]),
.IBG(vrtovaj[22]),
.IBH(vrtovaj[23]),
.IBI(vrtovaj[24]),
.IBJ(vrtovaj[25]),
.IBK(vrtovaj[26]),
.IBL(vrtovaj[27]),
.IBM(vrtovaj[28]),
.IBN(vrtovaj[29]),
.IBO(vrtovaj[30]),
.IBP(vrtovaj[31]),
.ICA(vrtovaj[32]),
.ICB(vrtovaj[33]),
.ICC(vrtovaj[34]),
.ICD(vrtovaj[35]),
.ICE(vrtovaj[36]),
.ICF(vrtovaj[37]),
.ICG(vrtovaj[38]),
.ICH(vrtovaj[39]),
.ICI(vrtovaj[40]),
.ICJ(vrtovaj[41]),
.ICK(vrtovaj[42]),
.ICL(vrtovaj[43]),
.ICM(vrtovaj[44]),
.ICN(vrtovaj[45]),
.ICO(vrtovaj[46]),
.ICP(vrtovaj[47]),
.IDA(vrtovaj[48]),
.IDB(vrtovaj[49]),
.IDC(vrtovaj[50]),
.IDD(vrtovaj[51]),
.IDE(vrtovaj[52]),
.IDF(vrtovaj[53]),
.IDG(vrtovaj[54]),
.IDH(vrtovaj[55]),
.IDI(vrtovaj[56]),
.IDJ(vrtovaj[57]),
.IDK(vrtovaj[58]),
.IDL(vrtovaj[59]),
.IDM(vrtovaj[60]),
.IDN(vrtovaj[61]),
.IDO(vrtovaj[62]),
.IDP(vrtovaj[63]),
.IEA(vrtovak[0]),
.IEB(vrtovak[1]),
.IEC(vrtovak[2]),
.IED(vrtovak[3]),
.IEE(vrtovak[4]),
.IEF(vrtovak[5]),
.IEG(vrtovak[6]),
.IEH(vrtovak[7]),
.IEI(vrtovak[8]),
.IEJ(vrtovak[9]),
.IEK(vrtovak[10]),
.IEL(vrtovak[11]),
.IEM(vrtovak[12]),
.IEN(vrtovak[13]),
.IEO(vrtovak[14]),
.IEP(vrtovak[15]),
.IFA(vrtovak[16]),
.IFB(vrtovak[17]),
.IFC(vrtovak[18]),
.IFD(vrtovak[19]),
.IFE(vrtovak[20]),
.IFFF(vrtovak[21]),
.IFG(vrtovak[22]),
.IFH(vrtovak[23]),
.IFI(vrtovak[24]),
.IFJ(vrtovak[25]),
.IFK(vrtovak[26]),
.IFL(vrtovak[27]),
.IFM(vrtovak[28]),
.IFN(vrtovak[29]),
.IFO(vrtovak[30]),
.IFP(vrtovak[31]),
.IGA(vrtovak[32]),
.IGB(vrtovak[33]),
.IGC(vrtovak[34]),
.IGD(vrtovak[35]),
.IGE(vrtovak[36]),
.IGF(vrtovak[37]),
.IGG(vrtovak[38]),
.IGH(vrtovak[39]),
.IGI(vrtovak[40]),
.IGJ(vrtovak[41]),
.IGK(vrtovak[42]),
.IGL(vrtovak[43]),
.IGM(vrtovak[44]),
.IGN(vrtovak[45]),
.IGO(vrtovak[46]),
.IGP(vrtovak[47]),
.IHA(vrtovak[48]),
.IHB(vrtovak[49]),
.IHC(vrtovak[50]),
.IHD(vrtovak[51]),
.IHE(vrtovak[52]),
.IHF(vrtovak[53]),
.IHG(vrtovak[54]),
.IHH(vrtovak[55]),
.IHI(vrtovak[56]),
.IHJ(vrtovak[57]),
.IHK(vrtovak[58]),
.IHL(vrtovak[59]),
.IHM(vrtovak[60]),
.IHN(vrtovak[61]),
.IHO(vrtovak[62]),
.IHP(vrtovak[63]),
.IMA(),
.IRA(javacntr[0]),
.IRB(javacntr[1]),
.IRC(javacntr[2]),
.IRD(javacntr[3]),
.IZZ (sysclock),
.OAA(vatovb[0]),
.OAB(vatovb[1]),
.OAC(vatovb[2]),
.OAD(vatovb[3]),
.OAE(vatovb[4]),
.OAF(vatovb[5]),
.OAG(vatovb[6]),
.OAH(vatovb[7]),
.OAI(vatovb[8]),
.OAJ(vatovb[9]),
.OAK(vatovb[10]),
.OAL(vatovb[11]),
.OAM(vatovb[12]),
.OAN(vatovb[13]),
.OAO(vatovb[14]),
.OAP(vatovb[15]),
.OBA(vatovb[16]),
.OBB(vatovb[17]),
.OBC(vatovb[18]),
.OBD(vatovb[19]),
.OBE(vatovb[20]),
.OBF(vatovb[21]),
.OBG(vatovb[22]),
.OBH(vatovb[23]),
.OBI(vatovb[24]),
.OBJ(vatovb[25]),
.OBK(vatovb[26]),
.OBL(vatovb[27]),
.OBM(vatovb[28]),
.OBN(vatovb[29]),
.OBO(vatovb[30]),
.OBP(vatovb[31]),
.OCA(vatovb[32]),
.OCB(vatovb[33]),
.OCC(vatovb[34]),
.OCD(vatovb[35]),
.OCE(vatovb[36]),
.OCF(vatovb[37]),
.OCG(vatovb[38]),
.OCH(vatovb[39]),
.OCI(vatovb[40]),
.OCJ(vatovb[41]),
.OCK(vatovb[42]),
.OCL(vatovb[43]),
.OCM(vatovb[44]),
.OCN(vatovb[45]),
.OCO(vatovb[46]),
.OCP(vatovb[47]),
.ODA(vatovb[48]),
.ODB(vatovb[49]),
.ODC(vatovb[50]),
.ODD(vatovb[51]),
.ODE(vatovb[52]),
.ODF(vatovb[53]),
.ODG(vatovb[54]),
.ODH(vatovb[55]),
.ODI(vatovb[56]),
.ODJ(vatovb[57]),
.ODK(vatovb[58]),
.ODL(vatovb[59]),
.ODM(vatovb[60]),
.ODN(vatovb[61]),
.ODO(vatovb[62]),
.ODP(vatovb[63]),
.OEA(relvitojb),
.OEB(reliota[0]),
.OEC(reliota[1]),
.OFA(enableiota[0]),
.OFB(enableiota[1]),
.ONA(gostreamgb));



vb vb0 ( 
.IAA(vrtovb[0]),
.IAB(vrtovb[1]),
.IAC(vrtovb[2]),
.IAD(vrtovb[3]),
.IAE(vrtovb[4]),
.IAF(vrtovb[5]),
.IAG(vrtovb[6]),
.IAH(vrtovb[7]),
.IAI(vrtovb[8]),
.IAJ(vrtovb[9]),
.IAK(vrtovb[10]),
.IAL(vrtovb[11]),
.IAM(vrtovb[12]),
.IAN(vrtovb[13]),
.IAO(vrtovb[14]),
.IAP(vrtovb[15]),
.IBA(vrtovb[16]),
.IBB(vrtovb[17]),
.IBC(vrtovb[18]),
.IBD(vrtovb[19]),
.IBE(vrtovb[20]),
.IBF(vrtovb[21]),
.IBG(vrtovb[22]),
.IBH(vrtovb[23]),
.IBI(vrtovb[24]),
.IBJ(vrtovb[25]),
.IBK(vrtovb[26]),
.IBL(vrtovb[27]),
.IBM(vrtovb[28]),
.IBN(vrtovb[29]),
.IBO(vrtovb[30]),
.IBP(vrtovb[31]),
.ICA(vrtovb[32]),
.ICB(vrtovb[33]),
.ICC(vrtovb[34]),
.ICD(vrtovb[35]),
.ICE(vrtovb[36]),
.ICF(vrtovb[37]),
.ICG(vrtovb[38]),
.ICH(vrtovb[39]),
.ICI(vrtovb[40]),
.ICJ(vrtovb[41]),
.ICK(vrtovb[42]),
.ICL(vrtovb[43]),
.ICM(vrtovb[44]),
.ICN(vrtovb[45]),
.ICO(vrtovb[46]),
.ICP(vrtovb[47]),
.IDA(vrtovb[48]),
.IDB(vrtovb[49]),
.IDC(vrtovb[50]),
.IDD(vrtovb[51]),
.IDE(vrtovb[52]),
.IDF(vrtovb[53]),
.IDG(vrtovb[54]),
.IDH(vrtovb[55]),
.IDI(vrtovb[56]),
.IDJ(vrtovb[57]),
.IDK(vrtovb[58]),
.IDL(vrtovb[59]),
.IDM(vrtovb[60]),
.IDN(vrtovb[61]),
.IDO(vrtovb[62]),
.IDP(vrtovb[63]),
.IEA(vatovb[0]),
.IEB(vatovb[1]),
.IEC(vatovb[2]),
.IED(vatovb[3]),
.IEE(vatovb[4]),
.IEF(vatovb[5]),
.IEG(vatovb[6]),
.IEH(vatovb[7]),
.IEI(vatovb[8]),
.IEJ(vatovb[9]),
.IEK(vatovb[10]),
.IEL(vatovb[11]),
.IEM(vatovb[12]),
.IEN(vatovb[13]),
.IEO(vatovb[14]),
.IEP(vatovb[15]),
.IFA(vatovb[16]),
.IFB(vatovb[17]),
.IFC(vatovb[18]),
.IFD(vatovb[19]),
.IFE(vatovb[20]),
.IFFF(vatovb[21]),
.IFG(vatovb[22]),
.IFH(vatovb[23]),
.IFI(vatovb[24]),
.IFJ(vatovb[25]),
.IFK(vatovb[26]),
.IFL(vatovb[27]),
.IFM(vatovb[28]),
.IFN(vatovb[29]),
.IFO(vatovb[30]),
.IFP(vatovb[31]),
.IGA(vatovb[32]),
.IGB(vatovb[33]),
.IGC(vatovb[34]),
.IGD(vatovb[35]),
.IGE(vatovb[36]),
.IGF(vatovb[37]),
.IGG(vatovb[38]),
.IGH(vatovb[39]),
.IGI(vatovb[40]),
.IGJ(vatovb[41]),
.IGK(vatovb[42]),
.IGL(vatovb[43]),
.IGM(vatovb[44]),
.IGN(vatovb[45]),
.IGO(vatovb[46]),
.IGP(vatovb[47]),
.IHA(vatovb[48]),
.IHB(vatovb[49]),
.IHC(vatovb[50]),
.IHD(vatovb[51]),
.IHE(vatovb[52]),
.IHF(vatovb[53]),
.IHG(vatovb[54]),
.IHH(vatovb[55]),
.IHI(vatovb[56]),
.IHJ(vatovb[57]),
.IHK(vatovb[58]),
.IHL(vatovb[59]),
.IHM(vatovb[60]),
.IHN(vatovb[61]),
.IHO(vatovb[62]),
.IHP(vatovb[63]),
.IIA(shtambtovb[0]),
.IIB(shtambtovb[1]),
.IIC(shtambtovb[2]),
.IID(shtambtovb[3]),
.IIE(shtambtovb[4]),
.IIF(shtambtovb[5]),
.IIG(shtambtovb[6]),
.ISA(javbcntr[0]),
.ISB(javbcntr[1]),
.ISC(javbcntr[2]),
.IZZ (sysclock),
.OAA(vbtovr[0]),
.OAB(vbtovr[1]),
.OAC(vbtovr[2]),
.OAD(vbtovr[3]),
.OAE(vbtovr[4]),
.OAF(vbtovr[5]),
.OAG(vbtovr[6]),
.OAH(vbtovr[7]),
.OAI(vbtovr[8]),
.OAJ(vbtovr[9]),
.OAK(vbtovr[10]),
.OAL(vbtovr[11]),
.OAM(vbtovr[12]),
.OAN(vbtovr[13]),
.OAO(vbtovr[14]),
.OAP(vbtovr[15]),
.OBA(vbtovr[16]),
.OBB(vbtovr[17]),
.OBC(vbtovr[18]),
.OBD(vbtovr[19]),
.OBE(vbtovr[20]),
.OBF(vbtovr[21]),
.OBG(vbtovr[22]),
.OBH(vbtovr[23]),
.OBI(vbtovr[24]),
.OBJ(vbtovr[25]),
.OBK(vbtovr[26]),
.OBL(vbtovr[27]),
.OBM(vbtovr[28]),
.OBN(vbtovr[29]),
.OBO(vbtovr[30]),
.OBP(vbtovr[31]),
.OCA(vbtovr[32]),
.OCB(vbtovr[33]),
.OCC(vbtovr[34]),
.OCD(vbtovr[35]),
.OCE(vbtovr[36]),
.OCF(vbtovr[37]),
.OCG(vbtovr[38]),
.OCH(vbtovr[39]),
.OCI(vbtovr[40]),
.OCJ(vbtovr[41]),
.OCK(vbtovr[42]),
.OCL(vbtovr[43]),
.OCM(vbtovr[44]),
.OCN(vbtovr[45]),
.OCO(vbtovr[46]),
.OCP(vbtovr[47]),
.ODA(vbtovr[48]),
.ODB(vbtovr[49]),
.ODC(vbtovr[50]),
.ODD(vbtovr[51]),
.ODE(vbtovr[52]),
.ODF(vbtovr[53]),
.ODG(vbtovr[54]),
.ODH(vbtovr[55]),
.ODI(vbtovr[56]),
.ODJ(vbtovr[57]),
.ODK(vbtovr[58]),
.ODL(vbtovr[59]),
.ODM(vbtovr[60]),
.ODN(vbtovr[61]),
.ODO(vbtovr[62]),
.ODP(vbtovr[63]));

vl vl0 (
.IAA(scaljtovl[0]),
.IAB(scaljtovl[1]),
.IAC(scaljtovl[2]),
.IAD(scaljtovl[3]),
.IAE(scaljtovl[4]),
.IAF(scaljtovl[5]),
.IAG(scaljtovl[6]),
.IAH(scaljtovl[7]),
.IAI(scaljtovl[8]),
.IAJ(scaljtovl[9]),
.IAK(scaljtovl[10]),
.IAL(scaljtovl[11]),
.IAM(scaljtovl[12]),
.IAN(scaljtovl[13]),
.IAO(scaljtovl[14]),
.IAP(scaljtovl[15]),
.IBA(scaljtovl[16]),
.IBB(scaljtovl[17]),
.IBC(scaljtovl[18]),
.IBD(scaljtovl[19]),
.IBE(scaljtovl[20]),
.IBF(scaljtovl[21]),
.IBG(scaljtovl[22]),
.IBH(scaljtovl[23]),
.IBI(scaljtovl[24]),
.IBJ(scaljtovl[25]),
.IBK(scaljtovl[26]),
.IBL(scaljtovl[27]),
.IBM(scaljtovl[28]),
.IBN(scaljtovl[29]),
.IBO(scaljtovl[30]),
.IBP(scaljtovl[31]),
.ICA(scaljtovl[32]),
.ICB(scaljtovl[33]),
.ICC(scaljtovl[34]),
.ICD(scaljtovl[35]),
.ICE(scaljtovl[36]),
.ICF(scaljtovl[37]),
.ICG(scaljtovl[38]),
.ICH(scaljtovl[39]),
.ICI(scaljtovl[40]),
.ICJ(scaljtovl[41]),
.ICK(scaljtovl[42]),
.ICL(scaljtovl[43]),
.ICM(scaljtovl[44]),
.ICN(scaljtovl[45]),
.ICO(scaljtovl[46]),
.ICP(scaljtovl[47]),
.IDA(scaljtovl[48]),
.IDB(scaljtovl[49]),
.IDC(scaljtovl[50]),
.IDD(scaljtovl[51]),
.IDE(scaljtovl[52]),
.IDF(scaljtovl[53]),
.IDG(scaljtovl[54]),
.IDH(scaljtovl[55]),
.IDI(scaljtovl[56]),
.IDJ(scaljtovl[57]),
.IDK(scaljtovl[58]),
.IDL(scaljtovl[59]),
.IDM(scaljtovl[60]),
.IDN(scaljtovl[61]),
.IDO(scaljtovl[62]),
.IDP(scaljtovl[63]),
.IEA(vrtovlk[0]),
.IEB(vrtovlk[1]),
.IEC(vrtovlk[2]),
.IED(vrtovlk[3]),
.IEE(vrtovlk[4]),
.IEF(vrtovlk[5]),
.IEG(vrtovlk[6]),
.IEH(vrtovlk[7]),
.IEI(vrtovlk[8]),
.IEJ(vrtovlk[9]),
.IEK(vrtovlk[10]),
.IEL(vrtovlk[11]),
.IEM(vrtovlk[12]),
.IEN(vrtovlk[13]),
.IEO(vrtovlk[14]),
.IEP(vrtovlk[15]),
.IFA(vrtovlk[16]),
.IFB(vrtovlk[17]),
.IFC(vrtovlk[18]),
.IFD(vrtovlk[19]),
.IFE(vrtovlk[20]),
.IFFF(vrtovlk[21]),
.IFG(vrtovlk[22]),
.IFH(vrtovlk[23]),
.IFI(vrtovlk[24]),
.IFJ(vrtovlk[25]),
.IFK(vrtovlk[26]),
.IFL(vrtovlk[27]),
.IFM(vrtovlk[28]),
.IFN(vrtovlk[29]),
.IFO(vrtovlk[30]),
.IFP(vrtovlk[31]),
.IGA(vrtovlk[32]),
.IGB(vrtovlk[33]),
.IGC(vrtovlk[34]),
.IGD(vrtovlk[35]),
.IGE(vrtovlk[36]),
.IGF(vrtovlk[37]),
.IGG(vrtovlk[38]),
.IGH(vrtovlk[39]),
.IGI(vrtovlk[40]),
.IGJ(vrtovlk[41]),
.IGK(vrtovlk[42]),
.IGL(vrtovlk[43]),
.IGM(vrtovlk[44]),
.IGN(vrtovlk[45]),
.IGO(vrtovlk[46]),
.IGP(vrtovlk[47]),
.IHA(vrtovlk[48]),
.IHB(vrtovlk[49]),
.IHC(vrtovlk[50]),
.IHD(vrtovlk[51]),
.IHE(vrtovlk[52]),
.IHF(vrtovlk[53]),
.IHG(vrtovlk[54]),
.IHH(vrtovlk[55]),
.IHI(vrtovlk[56]),
.IHJ(vrtovlk[57]),
.IHK(vrtovlk[58]),
.IHL(vrtovlk[59]),
.IHM(vrtovlk[60]),
.IHN(vrtovlk[61]),
.IHO(vrtovlk[62]),
.IHP(vrtovlk[63]),
.IIA(javlcnt[0]),
.IIB(javlcnt[1]),
.IIC(javlcnt[2]),
.IID(javlcnt[3]),
.IIE(javlcnt[4]),
.IIF(javlcnt[5]),
.IIG(javlcnt[6]),
.IJA(vectorenablefromjb),
.IZZ (sysclock),
.IZH (ihold),
.OAA(vltovr[0]),
.OAB(vltovr[1]),
.OAC(vltovr[2]),
.OAD(vltovr[3]),
.OAE(vltovr[4]),
.OAF(vltovr[5]),
.OAG(vltovr[6]),
.OAH(vltovr[7]),
.OAI(vltovr[8]),
.OAJ(vltovr[9]),
.OAK(vltovr[10]),
.OAL(vltovr[11]),
.OAM(vltovr[12]),
.OAN(vltovr[13]),
.OAO(vltovr[14]),
.OAP(vltovr[15]),
.OBA(vltovr[16]),
.OBB(vltovr[17]),
.OBC(vltovr[18]),
.OBD(vltovr[19]),
.OBE(vltovr[20]),
.OBF(vltovr[21]),
.OBG(vltovr[22]),
.OBH(vltovr[23]),
.OBI(vltovr[24]),
.OBJ(vltovr[25]),
.OBK(vltovr[26]),
.OBL(vltovr[27]),
.OBM(vltovr[28]),
.OBN(vltovr[29]),
.OBO(vltovr[30]),
.OBP(vltovr[31]),
.OCA(vltovr[32]),
.OCB(vltovr[33]),
.OCC(vltovr[34]),
.OCD(vltovr[35]),
.OCE(vltovr[36]),
.OCF(vltovr[37]),
.OCG(vltovr[38]),
.OCH(vltovr[39]),
.OCI(vltovr[40]),
.OCJ(vltovr[41]),
.OCK(vltovr[42]),
.OCL(vltovr[43]),
.OCM(vltovr[44]),
.OCN(vltovr[45]),
.OCO(vltovr[46]),
.OCP(vltovr[47]),
.ODA(vltovr[48]),
.ODB(vltovr[49]),
.ODC(vltovr[50]),
.ODD(vltovr[51]),
.ODE(vltovr[52]),
.ODF(vltovr[53]),
.ODG(vltovr[54]),
.ODH(vltovr[55]),
.ODI(vltovr[56]),
.ODJ(vltovr[57]),
.ODK(vltovr[58]),
.ODL(vltovr[59]),
.ODM(vltovr[60]),
.ODN(vltovr[61]),
.ODO(vltovr[62]),
.ODP(vltovr[63]));


vr vr0 ( 
.IAA(v0addr1[0]),
.IAB(v0addr1[1]),
.IAC(v0addr1[2]),
.IAD(v0addr1[3]),
.IAE(v0addr1[4]),
.IAF(v0addr1[5]),
.IAG(v0vectmode[0]),
.IAH(v0vectstep[0]),
.IBA(v1addr1[0]),
.IBB(v1addr1[1]),
.IBC(v1addr1[2]),
.IBD(v1addr1[3]),
.IBE(v1addr1[4]),
.IBF(v1addr1[5]),
.IBG(v1vectmode[0]),
.IBH(v1vectstep[0]),
.ICA(v2addr1[0]),
.ICB(v2addr1[1]),
.ICC(v2addr1[2]),
.ICD(v2addr1[3]),
.ICE(v2addr1[4]),
.ICF(v2addr1[5]),
.ICG(v2vectmode[0]),
.ICH(v2vectstep[0]),
.IDA(v3addr1[0]),
.IDB(v3addr1[1]),
.IDC(v3addr1[2]),
.IDD(v3addr1[3]),
.IDE(v3addr1[4]),
.IDF(v3addr1[5]),
.IDG(v3vectmode[0]),
.IDH(v3vectstep[0]),
.IEA(v4addr1[0]),
.IEB(v4addr1[1]),
.IEC(v4addr1[2]),
.IED(v4addr1[3]),
.IEE(v4addr1[4]),
.IEF(v4addr1[5]),
.IEG(v4vectmode[0]),
.IEH(v4vectstep[0]),
.IFA(v5addr1[0]),
.IFB(v5addr1[1]),
.IFC(v5addr1[2]),
.IFD(v5addr1[3]),
.IFE(v5addr1[4]),
.IFFF(v5addr1[5]),
.IFG(v5vectmode[0]),
.IFH(v5vectstep[0]),
.IGA(v6addr1[0]),
.IGB(v6addr1[1]),
.IGC(v6addr1[2]),
.IGD(v6addr1[3]),
.IGE(v6addr1[4]),
.IGF(v6addr1[5]),
.IGG(v6vectmode[0]),
.IGH(v6vectstep[0]),
.IHA(v7addr1[0]),
.IHB(v7addr1[1]),
.IHC(v7addr1[2]),
.IHD(v7addr1[3]),
.IHE(v7addr1[4]),
.IHF(v7addr1[5]),
.IHG(v7vectmode[0]),
.IHH(v7vectstep[0]),
.IIA(gatovr[0]),
.IIB(gatovr[1]),
.IIC(gatovr[2]),
.IID(gatovr[3]),
.IIE(gatovr[4]),
.IIF(gatovr[5]),
.IIG(gatovr[6]),
.IIH(gatovr[7]),
.IJA(gbtovr[0]),
.IJB(gbtovr[1]),
.IJC(gbtovr[2]),
.IJD(gbtovr[3]),
.IJE(gbtovr[4]),
.IJF(gbtovr[5]),
.IJG(gbtovr[6]),
.IJH(gbtovr[7]),
.IKA(vbtovr[0]),
.IKB(vbtovr[1]),
.IKC(vbtovr[2]),
.IKD(vbtovr[3]),
.IKE(vbtovr[4]),
.IKF(vbtovr[5]),
.IKG(vbtovr[6]),
.IKH(vbtovr[7]),
.IMA(vltovr[0]),
.IMB(vltovr[1]),
.IMC(vltovr[2]),
.IMD(vltovr[3]),
.IME(vltovr[4]),
.IMF(vltovr[5]),
.IMG(vltovr[6]),
.IMH(vltovr[7]),
.INA(fctovr[0]),
.INB(fctovr[1]),
.INC(fctovr[2]),
.IND(fctovr[3]),
.INE(fctovr[4]),
.INF(fctovr[5]),
.ING(fctovr[6]),
.INH(fctovr[7]),
.IOA(metovr[0]),
.IOB(metovr[1]),
.IOC(metovr[2]),
.IOD(metovr[3]),
.IOE(metovr[4]),
.IOF(metovr[5]),
.IOG(metovr[6]),
.IOH(metovr[7]),
.IPA(watovr[0]),
.IPB(watovr[1]),
.IPC(watovr[2]),
.IPD(watovr[3]),
.IPE(watovr[4]),
.IPF(watovr[5]),
.IPG(watovr[6]),
.IPH(watovr[7]),
.IQA(commemtovr[0]),
.IQB(commemtovr[1]),
.IQC(commemtovr[2]),
.IQD(commemtovr[3]),
.IQE(commemtovr[4]),
.IQF(commemtovr[5]),
.IQG(commemtovr[6]),
.IQH(commemtovr[7]),
.IRA(jbtovr[0]),
.IRB(jbtovr[1]),
.IRC(jbtovr[2]),
.IRD(jbtovr[3]),
.IRE(jbtovr[4]),
.IRF(jbtovr[5]),
.IRG(jbtovr[6]),
.IRH(jbtovr[7]),
.ISA(vector1srccode[0]),
.ISB(vector1srccode[1]),
.ISC(vector1srccode[2]),
.ISD(vector1srccode[3]),
.ISE(vector1srccode[4]),
.ISF(vector1srccode[5]),
.ISG(vector1srccode[6]),
.ITA(scaldesttovr0[0]),
.ITB(scaldesttovr0[1]),
.ITC(scaldesttovr0[2]),
.ITD(scaldesttovr0[3]),
.ITE(scaldesttovr0[4]),
.ITF(scaldesttovr0[5]),
.IZZ (sysclock),
.IZH(ihold),
.OAA(scdatatoga[0]),
.OAB(scdatatoga[1]),
.OAC(scdatatoga[2]),
.OAD(scdatatoga[3]),
.OAE(scdatatoga[4]),
.OAF(scdatatoga[5]),
.OAG(scdatatoga[6]),
.OAH(scdatatoga[7]),
.OBA(shdatatogb[0]),
.OBB(shdatatogb[1]),
.OBC(shdatatogb[2]),
.OBD(shdatatogb[3]),
.OBE(shdatatogb[4]),
.OBF(shdatatogb[5]),
.OBG(shdatatogb[6]),
.OBH(shdatatogb[7]),
.OCA(vrtoar[0]),
.OCB(vrtoar[1]),
.OCC(vrtoar[2]),
.OCD(vrtoar[3]),
.OCE(vrtoar[4]),
.OCF(vrtoar[5]),
.OCG(vrtoar[6]),
.OCH(vrtoar[7]),
.ODA(vrtovaj[0]),
.ODB(vrtovaj[1]),
.ODC(vrtovaj[2]),
.ODD(vrtovaj[3]),
.ODE(vrtovaj[4]),
.ODF(vrtovaj[5]),
.ODG(vrtovaj[6]),
.ODH(vrtovaj[7]),
.OEA(vrtovak[0]),
.OEB(vrtovak[1]),
.OEC(vrtovak[2]),
.OED(vrtovak[3]),
.OEE(vrtovak[4]),
.OEF(vrtovak[5]),
.OEG(vrtovak[6]),
.OEH(vrtovak[7]),
.OFA(vrtovb[0]),
.OFB(vrtovb[1]),
.OFC(vrtovb[2]),
.OFD(vrtovb[3]),
.OFE(vrtovb[4]),
.OFF(vrtovb[5]),
.OFG(vrtovb[6]),
.OFH(vrtovb[7]),
.OGA(scaljtovl[0]),
.OGB(scaljtovl[1]),
.OGC(scaljtovl[2]),
.OGD(scaljtovl[3]),
.OGE(scaljtovl[4]),
.OGF(scaljtovl[5]),
.OGG(scaljtovl[6]),
.OGH(scaljtovl[7]),
.OHA(vrtovlk[0]),
.OHB(vrtovlk[1]),
.OHC(vrtovlk[2]),
.OHD(vrtovlk[3]),
.OHE(vrtovlk[4]),
.OHF(vrtovlk[5]),
.OHG(vrtovlk[6]),
.OHH(vrtovlk[7]),
.OIA(vrtofaj[0]),
.OIB(vrtofaj[1]),
.OIC(vrtofaj[2]),
.OID(vrtofaj[3]),
.OIE(vrtofaj[4]),
.OIF(vrtofaj[5]),
.OIG(vrtofaj[6]),
.OIH(vrtofaj[7]),
.OJA(vrtofak[0]),
.OJB(vrtofak[1]),
.OJC(vrtofak[2]),
.OJD(vrtofak[3]),
.OJE(vrtofak[4]),
.OJF(vrtofak[5]),
.OJG(vrtofak[6]),
.OJH(vrtofak[7]),
.OKA(vrtomulj[0]),
.OKB(vrtomulj[1]),
.OKC(vrtomulj[2]),
.OKD(vrtomulj[3]),
.OKE(vrtomulj[4]),
.OKF(vrtomulj[5]),
.OKG(vrtomulj[6]),
.OKH(vrtomulj[7]),
.OLA(vrtomulk[0]),
.OLB(vrtomulk[1]),
.OLC(vrtomulk[2]),
.OLD(vrtomulk[3]),
.OLE(vrtomulk[4]),
.OLF(vrtomulk[5]),
.OLG(vrtomulk[6]),
.OLH(vrtomulk[7]),
.OMA(vrtolm[0]),
.OMB(vrtolm[1]),
.OMC(vrtolm[2]),
.OMD(vrtolm[3]),
.OME(vrtolm[4]),
.OMF(vrtolm[5]),
.OMG(vrtolm[6]),
.OMH(vrtolm[7]),
.ONA(vraddrtotf[0]),
.ONB(vraddrtotf[1]),
.ONC(vraddrtotf[2]),
.OND(vraddrtotf[3]),
.ONE(vraddrtotf[4]),
.ONF(vraddrtotf[5]),
.ONG(vraddrtotf[6]),
.ONH(vraddrtotf[7]),
.OOA(vrtocm[0]),
.OOB(vrtocm[1]),
.OOC(vrtocm[2]),
.OOD(vrtocm[3]),
.OOE(vrtocm[4]),
.OOF(vrtocm[5]),
.OOG(vrtocm[6]),
.OOH(vrtocm[7]),
.OQA(sregbrdata[0]),
.OQB(),
.ORA(lmparityeafrvr[0]));
   



vr vr1 ( 
.IAA(v0addr2[0]),
.IAB(v0addr2[1]),
.IAC(v0addr2[2]),
.IAD(v0addr2[3]),
.IAE(v0addr2[4]),
.IAF(v0addr2[5]),
.IAG(v0vectmode[1]),
.IAH(v0vectstep[1]),
.IBA(v1addr2[0]),
.IBB(v1addr2[1]),
.IBC(v1addr2[2]),
.IBD(v1addr2[3]),
.IBE(v1addr2[4]),
.IBF(v1addr2[5]),
.IBG(v1vectmode[1]),
.IBH(v1vectstep[1]),
.ICA(v2addr2[0]),
.ICB(v2addr2[1]),
.ICC(v2addr2[2]),
.ICD(v2addr2[3]),
.ICE(v2addr2[4]),
.ICF(v2addr2[5]),
.ICG(v2vectmode[1]),
.ICH(v2vectstep[1]),
.IDA(v3addr2[0]),
.IDB(v3addr2[1]),
.IDC(v3addr2[2]),
.IDD(v3addr2[3]),
.IDE(v3addr2[4]),
.IDF(v3addr2[5]),
.IDG(v3vectmode[1]),
.IDH(v3vectstep[1]),
.IEA(v4addr2[0]),
.IEB(v4addr2[1]),
.IEC(v4addr2[2]),
.IED(v4addr2[3]),
.IEE(v4addr2[4]),
.IEF(v4addr2[5]),
.IEG(v4vectmode[1]),
.IEH(v4vectstep[1]),
.IFA(v5addr2[0]),
.IFB(v5addr2[1]),
.IFC(v5addr2[2]),
.IFD(v5addr2[3]),
.IFE(v5addr2[4]),
.IFFF(v5addr2[5]),
.IFG(v5vectmode[1]),
.IFH(v5vectstep[1]),
.IGA(v6addr2[0]),
.IGB(v6addr2[1]),
.IGC(v6addr2[2]),
.IGD(v6addr2[3]),
.IGE(v6addr2[4]),
.IGF(v6addr2[5]),
.IGG(v6vectmode[1]),
.IGH(v6vectstep[1]),
.IHA(v7addr2[0]),
.IHB(v7addr2[1]),
.IHC(v7addr2[2]),
.IHD(v7addr2[3]),
.IHE(v7addr2[4]),
.IHF(v7addr2[5]),
.IHG(v7vectmode[1]),
.IHH(v7vectstep[1]),
.IIA(gatovr[8]),
.IIB(gatovr[9]),
.IIC(gatovr[10]),
.IID(gatovr[11]),
.IIE(gatovr[12]),
.IIF(gatovr[13]),
.IIG(gatovr[14]),
.IIH(gatovr[15]),
.IJA(gbtovr[8]),
.IJB(gbtovr[9]),
.IJC(gbtovr[10]),
.IJD(gbtovr[11]),
.IJE(gbtovr[12]),
.IJF(gbtovr[13]),
.IJG(gbtovr[14]),
.IJH(gbtovr[15]),
.IKA(vbtovr[8]),
.IKB(vbtovr[9]),
.IKC(vbtovr[10]),
.IKD(vbtovr[11]),
.IKE(vbtovr[12]),
.IKF(vbtovr[13]),
.IKG(vbtovr[14]),
.IKH(vbtovr[15]),
.IMA(vltovr[8]),
.IMB(vltovr[9]),
.IMC(vltovr[10]),
.IMD(vltovr[11]),
.IME(vltovr[12]),
.IMF(vltovr[13]),
.IMG(vltovr[14]),
.IMH(vltovr[15]),
.INA(fctovr[8]),
.INB(fctovr[9]),
.INC(fctovr[10]),
.IND(fctovr[11]),
.INE(fctovr[12]),
.INF(fctovr[13]),
.ING(fctovr[14]),
.INH(fctovr[15]),
.IOA(metovr[8]),
.IOB(metovr[9]),
.IOC(metovr[10]),
.IOD(metovr[11]),
.IOE(metovr[12]),
.IOF(metovr[13]),
.IOG(metovr[14]),
.IOH(metovr[15]),
.IPA(watovr[8]),
.IPB(watovr[9]),
.IPC(watovr[10]),
.IPD(watovr[11]),
.IPE(watovr[12]),
.IPF(watovr[13]),
.IPG(watovr[14]),
.IPH(watovr[15]),
.IQA(commemtovr[8]),
.IQB(commemtovr[9]),
.IQC(commemtovr[10]),
.IQD(commemtovr[11]),
.IQE(commemtovr[12]),
.IQF(commemtovr[13]),
.IQG(commemtovr[14]),
.IQH(commemtovr[15]),
.IRA(jbtovr[8]),
.IRB(jbtovr[9]),
.IRC(jbtovr[10]),
.IRD(jbtovr[11]),
.IRE(jbtovr[12]),
.IRF(jbtovr[13]),
.IRG(jbtovr[14]),
.IRH(jbtovr[15]),
.ISA(vector2srccode[0]),
.ISB(vector2srccode[1]),
.ISC(vector2srccode[2]),
.ISD(vector2srccode[3]),
.ISE(vector2srccode[4]),
.ISF(vector2srccode[5]),
.ISG(vector2srccode[6]),
.ITA(scaldesttovr1[0]),
.ITB(scaldesttovr1[1]),
.ITC(scaldesttovr1[2]),
.ITD(scaldesttovr1[3]),
.ITE(scaldesttovr1[4]),
.ITF(scaldesttovr1[5]),
.IZZ (sysclock),
.IZH(ihold),
.OAA(scdatatoga[8]),
.OAB(scdatatoga[9]),
.OAC(scdatatoga[10]),
.OAD(scdatatoga[11]),
.OAE(scdatatoga[12]),
.OAF(scdatatoga[13]),
.OAG(scdatatoga[14]),
.OAH(scdatatoga[15]),
.OBA(shdatatogb[8]),
.OBB(shdatatogb[9]),
.OBC(shdatatogb[10]),
.OBD(shdatatogb[11]),
.OBE(shdatatogb[12]),
.OBF(shdatatogb[13]),
.OBG(shdatatogb[14]),
.OBH(shdatatogb[15]),
.OCA(vrtoar[8]),
.OCB(vrtoar[9]),
.OCC(vrtoar[10]),
.OCD(vrtoar[11]),
.OCE(vrtoar[12]),
.OCF(vrtoar[13]),
.OCG(vrtoar[14]),
.OCH(vrtoar[15]),
.ODA(vrtovaj[8]),
.ODB(vrtovaj[9]),
.ODC(vrtovaj[10]),
.ODD(vrtovaj[11]),
.ODE(vrtovaj[12]),
.ODF(vrtovaj[13]),
.ODG(vrtovaj[14]),
.ODH(vrtovaj[15]),
.OEA(vrtovak[8]),
.OEB(vrtovak[9]),
.OEC(vrtovak[10]),
.OED(vrtovak[11]),
.OEE(vrtovak[12]),
.OEF(vrtovak[13]),
.OEG(vrtovak[14]),
.OEH(vrtovak[15]),
.OFA(vrtovb[8]),
.OFB(vrtovb[9]),
.OFC(vrtovb[10]),
.OFD(vrtovb[11]),
.OFE(vrtovb[12]),
.OFF(vrtovb[13]),
.OFG(vrtovb[14]),
.OFH(vrtovb[15]),
.OGA(scaljtovl[8]),
.OGB(scaljtovl[9]),
.OGC(scaljtovl[10]),
.OGD(scaljtovl[11]),
.OGE(scaljtovl[12]),
.OGF(scaljtovl[13]),
.OGG(scaljtovl[14]),
.OGH(scaljtovl[15]),
.OHA(vrtovlk[8]),
.OHB(vrtovlk[9]),
.OHC(vrtovlk[10]),
.OHD(vrtovlk[11]),
.OHE(vrtovlk[12]),
.OHF(vrtovlk[13]),
.OHG(vrtovlk[14]),
.OHH(vrtovlk[15]),
.OIA(vrtofaj[8]),
.OIB(vrtofaj[9]),
.OIC(vrtofaj[10]),
.OID(vrtofaj[11]),
.OIE(vrtofaj[12]),
.OIF(vrtofaj[13]),
.OIG(vrtofaj[14]),
.OIH(vrtofaj[15]),
.OJA(vrtofak[8]),
.OJB(vrtofak[9]),
.OJC(vrtofak[10]),
.OJD(vrtofak[11]),
.OJE(vrtofak[12]),
.OJF(vrtofak[13]),
.OJG(vrtofak[14]),
.OJH(vrtofak[15]),
.OKA(vrtomulj[8]),
.OKB(vrtomulj[9]),
.OKC(vrtomulj[10]),
.OKD(vrtomulj[11]),
.OKE(vrtomulj[12]),
.OKF(vrtomulj[13]),
.OKG(vrtomulj[14]),
.OKH(vrtomulj[15]),
.OLA(vrtomulk[8]),
.OLB(vrtomulk[9]),
.OLC(vrtomulk[10]),
.OLD(vrtomulk[11]),
.OLE(vrtomulk[12]),
.OLF(vrtomulk[13]),
.OLG(vrtomulk[14]),
.OLH(vrtomulk[15]),
.OMA(vrtolm[8]),
.OMB(vrtolm[9]),
.OMC(vrtolm[10]),
.OMD(vrtolm[11]),
.OME(vrtolm[12]),
.OMF(vrtolm[13]),
.OMG(vrtolm[14]),
.OMH(vrtolm[15]),
.ONA(vraddrtotf[8]),
.ONB(vraddrtotf[9]),
.ONC(vraddrtotf[10]),
.OND(vraddrtotf[11]),
.ONE(vraddrtotf[12]),
.ONF(vraddrtotf[13]),
.ONG(vraddrtotf[14]),
.ONH(vraddrtotf[15]),
.OOA(vrtocm[8]),
.OOB(vrtocm[9]),
.OOC(vrtocm[10]),
.OOD(vrtocm[11]),
.OOE(vrtocm[12]),
.OOF(vrtocm[13]),
.OOG(vrtocm[14]),
.OOH(vrtocm[15]),
.OQA(sregbrdata[1]),
.OQB(),
.ORA(lmparityeafrvr[1]));


vr vr2 (
.IAA(v0addr3[0]),
.IAB(v0addr3[1]),
.IAC(v0addr3[2]),
.IAD(v0addr3[3]),
.IAE(v0addr3[4]),
.IAF(v0addr3[5]),
.IAG(v0vectmode[2]),
.IAH(v0vectstep[2]),
.IBA(v1addr3[0]),
.IBB(v1addr3[1]),
.IBC(v1addr3[2]),
.IBD(v1addr3[3]),
.IBE(v1addr3[4]),
.IBF(v1addr3[5]),
.IBG(v1vectmode[2]),
.IBH(v1vectstep[2]),
.ICA(v2addr3[0]),
.ICB(v2addr3[1]),
.ICC(v2addr3[2]),
.ICD(v2addr3[3]),
.ICE(v2addr3[4]),
.ICF(v2addr3[5]),
.ICG(v2vectmode[2]),
.ICH(v2vectstep[2]),
.IDA(v3addr3[0]),
.IDB(v3addr3[1]),
.IDC(v3addr3[2]),
.IDD(v3addr3[3]),
.IDE(v3addr3[4]),
.IDF(v3addr3[5]),
.IDG(v3vectmode[2]),
.IDH(v3vectstep[2]),
.IEA(v4addr3[0]),
.IEB(v4addr3[1]),
.IEC(v4addr3[2]),
.IED(v4addr3[3]),
.IEE(v4addr3[4]),
.IEF(v4addr3[5]),
.IEG(v4vectmode[2]),
.IEH(v4vectstep[2]),
.IFA(v5addr3[0]),
.IFB(v5addr3[1]),
.IFC(v5addr3[2]),
.IFD(v5addr3[3]),
.IFE(v5addr3[4]),
.IFFF(v5addr3[5]),
.IFG(v5vectmode[2]),
.IFH(v5vectstep[2]),
.IGA(v6addr3[0]),
.IGB(v6addr3[1]),
.IGC(v6addr3[2]),
.IGD(v6addr3[3]),
.IGE(v6addr3[4]),
.IGF(v6addr3[5]),
.IGG(v6vectmode[2]),
.IGH(v6vectstep[2]),
.IHA(v7addr3[0]),
.IHB(v7addr3[1]),
.IHC(v7addr3[2]),
.IHD(v7addr3[3]),
.IHE(v7addr3[4]),
.IHF(v7addr3[5]),
.IHG(v7vectmode[2]),
.IHH(v7vectstep[2]),
.IIA(gatovr[16]),
.IIB(gatovr[17]),
.IIC(gatovr[18]),
.IID(gatovr[19]),
.IIE(gatovr[20]),
.IIF(gatovr[21]),
.IIG(gatovr[22]),
.IIH(gatovr[23]),
.IJA(gbtovr[16]),
.IJB(gbtovr[17]),
.IJC(gbtovr[18]),
.IJD(gbtovr[19]),
.IJE(gbtovr[20]),
.IJF(gbtovr[21]),
.IJG(gbtovr[22]),
.IJH(gbtovr[23]),
.IKA(vbtovr[16]),
.IKB(vbtovr[17]),
.IKC(vbtovr[18]),
.IKD(vbtovr[19]),
.IKE(vbtovr[20]),
.IKF(vbtovr[21]),
.IKG(vbtovr[22]),
.IKH(vbtovr[23]),
.IMA(vltovr[16]),
.IMB(vltovr[17]),
.IMC(vltovr[18]),
.IMD(vltovr[19]),
.IME(vltovr[20]),
.IMF(vltovr[21]),
.IMG(vltovr[22]),
.IMH(vltovr[23]),
.INA(fctovr[16]),
.INB(fctovr[17]),
.INC(fctovr[18]),
.IND(fctovr[19]),
.INE(fctovr[20]),
.INF(fctovr[21]),
.ING(fctovr[22]),
.INH(fctovr[23]),
.IOA(metovr[16]),
.IOB(metovr[17]),
.IOC(metovr[18]),
.IOD(metovr[19]),
.IOE(metovr[20]),
.IOF(metovr[21]),
.IOG(metovr[22]),
.IOH(metovr[23]),
.IPA(watovr[16]),
.IPB(watovr[17]),
.IPC(watovr[18]),
.IPD(watovr[19]),
.IPE(watovr[20]),
.IPF(watovr[21]),
.IPG(watovr[22]),
.IPH(watovr[23]),
.IQA(commemtovr[16]),
.IQB(commemtovr[17]),
.IQC(commemtovr[18]),
.IQD(commemtovr[19]),
.IQE(commemtovr[20]),
.IQF(commemtovr[21]),
.IQG(commemtovr[22]),
.IQH(commemtovr[23]),
.IRA(jbtovr[16]),
.IRB(jbtovr[17]),
.IRC(jbtovr[18]),
.IRD(jbtovr[19]),
.IRE(jbtovr[20]),
.IRF(jbtovr[21]),
.IRG(jbtovr[22]),
.IRH(jbtovr[23]),
.ISA(vector3srccode[0]),
.ISB(vector3srccode[1]),
.ISC(vector3srccode[2]),
.ISD(vector3srccode[3]),
.ISE(vector3srccode[4]),
.ISF(vector3srccode[5]),
.ISG(vector3srccode[6]),
.ITA(scaldesttovr2[0]),
.ITB(scaldesttovr2[1]),
.ITC(scaldesttovr2[2]),
.ITD(scaldesttovr2[3]),
.ITE(scaldesttovr2[4]),
.ITF(scaldesttovr2[5]),
.IZZ (sysclock),
.IZH (ihold),
.OAA(scdatatoga[16]),
.OAB(scdatatoga[17]),
.OAC(scdatatoga[18]),
.OAD(scdatatoga[19]),
.OAE(scdatatoga[20]),
.OAF(scdatatoga[21]),
.OAG(scdatatoga[22]),
.OAH(scdatatoga[23]),
.OBA(shdatatogb[16]),
.OBB(shdatatogb[17]),
.OBC(shdatatogb[18]),
.OBD(shdatatogb[19]),
.OBE(shdatatogb[20]),
.OBF(shdatatogb[21]),
.OBG(shdatatogb[22]),
.OBH(shdatatogb[23]),
.OCA(vrtoar[16]),
.OCB(vrtoar[17]),
.OCC(vrtoar[18]),
.OCD(vrtoar[19]),
.OCE(vrtoar[20]),
.OCF(vrtoar[21]),
.OCG(vrtoar[22]),
.OCH(vrtoar[23]),
.ODA(vrtovaj[16]),
.ODB(vrtovaj[17]),
.ODC(vrtovaj[18]),
.ODD(vrtovaj[19]),
.ODE(vrtovaj[20]),
.ODF(vrtovaj[21]),
.ODG(vrtovaj[22]),
.ODH(vrtovaj[23]),
.OEA(vrtovak[16]),
.OEB(vrtovak[17]),
.OEC(vrtovak[18]),
.OED(vrtovak[19]),
.OEE(vrtovak[20]),
.OEF(vrtovak[21]),
.OEG(vrtovak[22]),
.OEH(vrtovak[23]),
.OFA(vrtovb[16]),
.OFB(vrtovb[17]),
.OFC(vrtovb[18]),
.OFD(vrtovb[19]),
.OFE(vrtovb[20]),
.OFF(vrtovb[21]),
.OFG(vrtovb[22]),
.OFH(vrtovb[23]),
.OGA(scaljtovl[16]),
.OGB(scaljtovl[17]),
.OGC(scaljtovl[18]),
.OGD(scaljtovl[19]),
.OGE(scaljtovl[20]),
.OGF(scaljtovl[21]),
.OGG(scaljtovl[22]),
.OGH(scaljtovl[23]),
.OHA(vrtovlk[16]),
.OHB(vrtovlk[17]),
.OHC(vrtovlk[18]),
.OHD(vrtovlk[19]),
.OHE(vrtovlk[20]),
.OHF(vrtovlk[21]),
.OHG(vrtovlk[22]),
.OHH(vrtovlk[23]),
.OIA(vrtofaj[16]),
.OIB(vrtofaj[17]),
.OIC(vrtofaj[18]),
.OID(vrtofaj[19]),
.OIE(vrtofaj[20]),
.OIF(vrtofaj[21]),
.OIG(vrtofaj[22]),
.OIH(vrtofaj[23]),
.OJA(vrtofak[16]),
.OJB(vrtofak[17]),
.OJC(vrtofak[18]),
.OJD(vrtofak[19]),
.OJE(vrtofak[20]),
.OJF(vrtofak[21]),
.OJG(vrtofak[22]),
.OJH(vrtofak[23]),
.OKA(vrtomulj[16]),
.OKB(vrtomulj[17]),
.OKC(vrtomulj[18]),
.OKD(vrtomulj[19]),
.OKE(vrtomulj[20]),
.OKF(vrtomulj[21]),
.OKG(vrtomulj[22]),
.OKH(vrtomulj[23]),
.OLA(vrtomulk[16]),
.OLB(vrtomulk[17]),
.OLC(vrtomulk[18]),
.OLD(vrtomulk[19]),
.OLE(vrtomulk[20]),
.OLF(vrtomulk[21]),
.OLG(vrtomulk[22]),
.OLH(vrtomulk[23]),
.OMA(vrtolm[16]),
.OMB(vrtolm[17]),
.OMC(vrtolm[18]),
.OMD(vrtolm[19]),
.OME(vrtolm[20]),
.OMF(vrtolm[21]),
.OMG(vrtolm[22]),
.OMH(vrtolm[23]),
.ONA(vraddrtotf[16]),
.ONB(vraddrtotf[17]),
.ONC(vraddrtotf[18]),
.OND(vraddrtotf[19]),
.ONE(vraddrtotf[20]),
.ONF(vraddrtotf[21]),
.ONG(vraddrtotf[22]),
.ONH(vraddrtotf[23]),
.OOA(vrtocm[16]),
.OOB(vrtocm[17]),
.OOC(vrtocm[18]),
.OOD(vrtocm[19]),
.OOE(vrtocm[20]),
.OOF(vrtocm[21]),
.OOG(vrtocm[22]),
.OOH(vrtocm[23]),
.OQA(sregbrdata[2]),
.OQB(),
.ORA(lmparityeafrvr[2]));

  
vr vr3 (
.IAA(v0addr4[0]),
.IAB(v0addr4[1]),
.IAC(v0addr4[2]),
.IAD(v0addr4[3]),
.IAE(v0addr4[4]),
.IAF(v0addr4[5]),
.IAG(v0vectmode[3]),
.IAH(v0vectstep[3]),
.IBA(v1addr4[0]),
.IBB(v1addr4[1]),
.IBC(v1addr4[2]),
.IBD(v1addr4[3]),
.IBE(v1addr4[4]),
.IBF(v1addr4[5]),
.IBG(v1vectmode[3]),
.IBH(v1vectstep[3]),
.ICA(v2addr4[0]),
.ICB(v2addr4[1]),
.ICC(v2addr4[2]),
.ICD(v2addr4[3]),
.ICE(v2addr4[4]),
.ICF(v2addr4[5]),
.ICG(v2vectmode[3]),
.ICH(v2vectstep[3]),
.IDA(v3addr4[0]),
.IDB(v3addr4[1]),
.IDC(v3addr4[2]),
.IDD(v3addr4[3]),
.IDE(v3addr4[4]),
.IDF(v3addr4[5]),
.IDG(v3vectmode[3]),
.IDH(v3vectstep[3]),
.IEA(v4addr4[0]),
.IEB(v4addr4[1]),
.IEC(v4addr4[2]),
.IED(v4addr4[3]),
.IEE(v4addr4[4]),
.IEF(v4addr4[5]),
.IEG(v4vectmode[3]),
.IEH(v4vectstep[3]),
.IFA(v5addr4[0]),
.IFB(v5addr4[1]),
.IFC(v5addr4[2]),
.IFD(v5addr4[3]),
.IFE(v5addr4[4]),
.IFFF(v5addr4[5]),
.IFG(v5vectmode[3]),
.IFH(v5vectstep[3]),
.IGA(v6addr4[0]),
.IGB(v6addr4[1]),
.IGC(v6addr4[2]),
.IGD(v6addr4[3]),
.IGE(v6addr4[4]),
.IGF(v6addr4[5]),
.IGG(v6vectmode[3]),
.IGH(v6vectstep[3]),
.IHA(v7addr4[0]),
.IHB(v7addr4[1]),
.IHC(v7addr4[2]),
.IHD(v7addr4[3]),
.IHE(v7addr4[4]),
.IHF(v7addr4[5]),
.IHG(v7vectmode[3]),
.IHH(v7vectstep[3]),
.IIA(gatovr[24]),
.IIB(gatovr[25]),
.IIC(gatovr[26]),
.IID(gatovr[27]),
.IIE(gatovr[28]),
.IIF(gatovr[29]),
.IIG(gatovr[30]),
.IIH(gatovr[31]),
.IJA(gbtovr[24]),
.IJB(gbtovr[25]),
.IJC(gbtovr[26]),
.IJD(gbtovr[27]),
.IJE(gbtovr[28]),
.IJF(gbtovr[29]),
.IJG(gbtovr[30]),
.IJH(gbtovr[31]),
.IKA(vbtovr[24]),
.IKB(vbtovr[25]),
.IKC(vbtovr[26]),
.IKD(vbtovr[27]),
.IKE(vbtovr[28]),
.IKF(vbtovr[29]),
.IKG(vbtovr[30]),
.IKH(vbtovr[31]),
.IMA(vltovr[24]),
.IMB(vltovr[25]),
.IMC(vltovr[26]),
.IMD(vltovr[27]),
.IME(vltovr[28]),
.IMF(vltovr[29]),
.IMG(vltovr[30]),
.IMH(vltovr[31]),
.INA(fctovr[24]),
.INB(fctovr[25]),
.INC(fctovr[26]),
.IND(fctovr[27]),
.INE(fctovr[28]),
.INF(fctovr[29]),
.ING(fctovr[30]),
.INH(fctovr[31]),
.IOA(metovr[24]),
.IOB(metovr[25]),
.IOC(metovr[26]),
.IOD(metovr[27]),
.IOE(metovr[28]),
.IOF(metovr[29]),
.IOG(metovr[30]),
.IOH(metovr[31]),
.IPA(watovr[24]),
.IPB(watovr[25]),
.IPC(watovr[26]),
.IPD(watovr[27]),
.IPE(watovr[28]),
.IPF(watovr[29]),
.IPG(watovr[30]),
.IPH(watovr[31]),
.IQA(commemtovr[24]),
.IQB(commemtovr[25]),
.IQC(commemtovr[26]),
.IQD(commemtovr[27]),
.IQE(commemtovr[28]),
.IQF(commemtovr[29]),
.IQG(commemtovr[30]),
.IQH(commemtovr[31]),
.IRA(jbtovr[24]),
.IRB(jbtovr[25]),
.IRC(jbtovr[26]),
.IRD(jbtovr[27]),
.IRE(jbtovr[28]),
.IRF(jbtovr[29]),
.IRG(jbtovr[30]),
.IRH(jbtovr[31]),
.ISA(vector4srccode[0]),
.ISB(vector4srccode[1]),
.ISC(vector4srccode[2]),
.ISD(vector4srccode[3]),
.ISE(vector4srccode[4]),
.ISF(vector4srccode[5]),
.ISG(vector4srccode[6]),
.ITA(scaldesttovr3[0]),
.ITB(scaldesttovr3[1]),
.ITC(scaldesttovr3[2]),
.ITD(scaldesttovr3[3]),
.ITE(scaldesttovr3[4]),
.ITF(scaldesttovr3[5]),
.IZZ (sysclock),
.IZH (ihold),
.OAA(scdatatoga[24]),
.OAB(scdatatoga[25]),
.OAC(scdatatoga[26]),
.OAD(scdatatoga[27]),
.OAE(scdatatoga[28]),
.OAF(scdatatoga[29]),
.OAG(scdatatoga[30]),
.OAH(scdatatoga[31]),
.OBA(shdatatogb[24]),
.OBB(shdatatogb[25]),
.OBC(shdatatogb[26]),
.OBD(shdatatogb[27]),
.OBE(shdatatogb[28]),
.OBF(shdatatogb[29]),
.OBG(shdatatogb[30]),
.OBH(shdatatogb[31]),
.OCA(vrtoar[24]),
.OCB(vrtoar[25]),
.OCC(vrtoar[26]),
.OCD(vrtoar[27]),
.OCE(vrtoar[28]),
.OCF(vrtoar[29]),
.OCG(vrtoar[30]),
.OCH(vrtoar[31]),
.ODA(vrtovaj[24]),
.ODB(vrtovaj[25]),
.ODC(vrtovaj[26]),
.ODD(vrtovaj[27]),
.ODE(vrtovaj[28]),
.ODF(vrtovaj[29]),
.ODG(vrtovaj[30]),
.ODH(vrtovaj[31]),
.OEA(vrtovak[24]),
.OEB(vrtovak[25]),
.OEC(vrtovak[26]),
.OED(vrtovak[27]),
.OEE(vrtovak[28]),
.OEF(vrtovak[29]),
.OEG(vrtovak[30]),
.OEH(vrtovak[31]),
.OFA(vrtovb[24]),
.OFB(vrtovb[25]),
.OFC(vrtovb[26]),
.OFD(vrtovb[27]),
.OFE(vrtovb[28]),
.OFF(vrtovb[29]),
.OFG(vrtovb[30]),
.OFH(vrtovb[31]),
.OGA(scaljtovl[24]),
.OGB(scaljtovl[25]),
.OGC(scaljtovl[26]),
.OGD(scaljtovl[27]),
.OGE(scaljtovl[28]),
.OGF(scaljtovl[29]),
.OGG(scaljtovl[30]),
.OGH(scaljtovl[31]),
.OHA(vrtovlk[24]),
.OHB(vrtovlk[25]),
.OHC(vrtovlk[26]),
.OHD(vrtovlk[27]),
.OHE(vrtovlk[28]),
.OHF(vrtovlk[29]),
.OHG(vrtovlk[30]),
.OHH(vrtovlk[31]),
.OIA(vrtofaj[24]),
.OIB(vrtofaj[25]),
.OIC(vrtofaj[26]),
.OID(vrtofaj[27]),
.OIE(vrtofaj[28]),
.OIF(vrtofaj[29]),
.OIG(vrtofaj[30]),
.OIH(vrtofaj[31]),
.OJA(vrtofak[24]),
.OJB(vrtofak[25]),
.OJC(vrtofak[26]),
.OJD(vrtofak[27]),
.OJE(vrtofak[28]),
.OJF(vrtofak[29]),
.OJG(vrtofak[30]),
.OJH(vrtofak[31]),
.OKA(vrtomulj[24]),
.OKB(vrtomulj[25]),
.OKC(vrtomulj[26]),
.OKD(vrtomulj[27]),
.OKE(vrtomulj[28]),
.OKF(vrtomulj[29]),
.OKG(vrtomulj[30]),
.OKH(vrtomulj[31]),
.OLA(vrtomulk[24]),
.OLB(vrtomulk[25]),
.OLC(vrtomulk[26]),
.OLD(vrtomulk[27]),
.OLE(vrtomulk[28]),
.OLF(vrtomulk[29]),
.OLG(vrtomulk[30]),
.OLH(vrtomulk[31]),
.OMA(vrtolm[24]),
.OMB(vrtolm[25]),
.OMC(vrtolm[26]),
.OMD(vrtolm[27]),
.OME(vrtolm[28]),
.OMF(vrtolm[29]),
.OMG(vrtolm[30]),
.OMH(vrtolm[31]),
.ONA(vraddrtotf[24]),
.ONB(vraddrtotf[25]),
.ONC(vraddrtotf[26]),
.OND(vraddrtotf[27]),
.ONE(vraddrtotf[28]),
.ONF(vraddrtotf[29]),
.ONG(vraddrtotf[30]),
.ONH(vraddrtotf[31]),
.OOA(vrtocm[24]),
.OOB(vrtocm[25]),
.OOC(vrtocm[26]),
.OOD(vrtocm[27]),
.OOE(vrtocm[28]),
.OOF(vrtocm[29]),
.OOG(vrtocm[30]),
.OOH(vrtocm[31]),
.OQA(sregbrdata[3]),
.OQB(),
.ORA(lmparityeafrvr[3]));
   



vr vr4 ( 
.IAA(v0addr5[0]),
.IAB(v0addr5[1]),
.IAC(v0addr5[2]),
.IAD(v0addr5[3]),
.IAE(v0addr5[4]),
.IAF(v0addr5[5]),
.IAG(v0vectmode[4]),
.IAH(v0vectstep[4]),
.IBA(v1addr5[0]),
.IBB(v1addr5[1]),
.IBC(v1addr5[2]),
.IBD(v1addr5[3]),
.IBE(v1addr5[4]),
.IBF(v1addr5[5]),
.IBG(v1vectmode[4]),
.IBH(v1vectstep[4]),
.ICA(v2addr5[0]),
.ICB(v2addr5[1]),
.ICC(v2addr5[2]),
.ICD(v2addr5[3]),
.ICE(v2addr5[4]),
.ICF(v2addr5[5]),
.ICG(v2vectmode[4]),
.ICH(v2vectstep[4]),
.IDA(v3addr5[0]),
.IDB(v3addr5[1]),
.IDC(v3addr5[2]),
.IDD(v3addr5[3]),
.IDE(v3addr5[4]),
.IDF(v3addr5[5]),
.IDG(v3vectmode[4]),
.IDH(v3vectstep[4]),
.IEA(v4addr5[0]),
.IEB(v4addr5[1]),
.IEC(v4addr5[2]),
.IED(v4addr5[3]),
.IEE(v4addr5[4]),
.IEF(v4addr5[5]),
.IEG(v4vectmode[4]),
.IEH(v4vectstep[4]),
.IFA(v5addr5[0]),
.IFB(v5addr5[1]),
.IFC(v5addr5[2]),
.IFD(v5addr5[3]),
.IFE(v5addr5[4]),
.IFFF(v5addr5[5]),
.IFG(v5vectmode[4]),
.IFH(v5vectstep[4]),
.IGA(v6addr5[0]),
.IGB(v6addr5[1]),
.IGC(v6addr5[2]),
.IGD(v6addr5[3]),
.IGE(v6addr5[4]),
.IGF(v6addr5[5]),
.IGG(v6vectmode[4]),
.IGH(v6vectstep[4]),
.IHA(v7addr5[0]),
.IHB(v7addr5[1]),
.IHC(v7addr5[2]),
.IHD(v7addr5[3]),
.IHE(v7addr5[4]),
.IHF(v7addr5[5]),
.IHG(v7vectmode[4]),
.IHH(v7vectstep[4]),
.IIA(gatovr[32]),
.IIB(gatovr[33]),
.IIC(gatovr[34]),
.IID(gatovr[35]),
.IIE(gatovr[36]),
.IIF(gatovr[37]),
.IIG(gatovr[38]),
.IIH(gatovr[39]),
.IJA(gbtovr[32]),
.IJB(gbtovr[33]),
.IJC(gbtovr[34]),
.IJD(gbtovr[35]),
.IJE(gbtovr[36]),
.IJF(gbtovr[37]),
.IJG(gbtovr[38]),
.IJH(gbtovr[39]),
.IKA(vbtovr[32]),
.IKB(vbtovr[33]),
.IKC(vbtovr[34]),
.IKD(vbtovr[35]),
.IKE(vbtovr[36]),
.IKF(vbtovr[37]),
.IKG(vbtovr[38]),
.IKH(vbtovr[39]),
.IMA(vltovr[32]),
.IMB(vltovr[33]),
.IMC(vltovr[34]),
.IMD(vltovr[35]),
.IME(vltovr[36]),
.IMF(vltovr[37]),
.IMG(vltovr[38]),
.IMH(vltovr[39]),
.INA(fctovr[32]),
.INB(fctovr[33]),
.INC(fctovr[34]),
.IND(fctovr[35]),
.INE(fctovr[36]),
.INF(fctovr[37]),
.ING(fctovr[38]),
.INH(fctovr[39]),
.IOA(metovr[32]),
.IOB(metovr[33]),
.IOC(metovr[34]),
.IOD(metovr[35]),
.IOE(metovr[36]),
.IOF(metovr[37]),
.IOG(metovr[38]),
.IOH(metovr[39]),
.IPA(watovr[32]),
.IPB(watovr[33]),
.IPC(watovr[34]),
.IPD(watovr[35]),
.IPE(watovr[36]),
.IPF(watovr[37]),
.IPG(watovr[38]),
.IPH(watovr[39]),
.IQA(commemtovr[32]),
.IQB(commemtovr[33]),
.IQC(commemtovr[34]),
.IQD(commemtovr[35]),
.IQE(commemtovr[36]),
.IQF(commemtovr[37]),
.IQG(commemtovr[38]),
.IQH(commemtovr[39]),
.IRA(jbtovr[32]),
.IRB(jbtovr[33]),
.IRC(jbtovr[34]),
.IRD(jbtovr[35]),
.IRE(jbtovr[36]),
.IRF(jbtovr[37]),
.IRG(jbtovr[38]),
.IRH(jbtovr[39]),
.ISA(vector5srccode[0]),
.ISB(vector5srccode[1]),
.ISC(vector5srccode[2]),
.ISD(vector5srccode[3]),
.ISE(vector5srccode[4]),
.ISF(vector5srccode[5]),
.ISG(vector5srccode[6]),
.ITA(scaldesttovr4[0]),
.ITB(scaldesttovr4[1]),
.ITC(scaldesttovr4[2]),
.ITD(scaldesttovr4[3]),
.ITE(scaldesttovr4[4]),
.ITF(scaldesttovr4[5]),
.IZZ (sysclock),
.IZH (ihold),
.OAA(scdatatoga[32]),
.OAB(scdatatoga[33]),
.OAC(scdatatoga[34]),
.OAD(scdatatoga[35]),
.OAE(scdatatoga[36]),
.OAF(scdatatoga[37]),
.OAG(scdatatoga[38]),
.OAH(scdatatoga[39]),
.OBA(shdatatogb[32]),
.OBB(shdatatogb[33]),
.OBC(shdatatogb[34]),
.OBD(shdatatogb[35]),
.OBE(shdatatogb[36]),
.OBF(shdatatogb[37]),
.OBG(shdatatogb[38]),
.OBH(shdatatogb[39]),
.OCA(),
.OCB(),
.OCC(),
.OCD(),
.OCE(),
.OCF(),
.OCG(),
.OCH(),
.ODA(vrtovaj[32]),
.ODB(vrtovaj[33]),
.ODC(vrtovaj[34]),
.ODD(vrtovaj[35]),
.ODE(vrtovaj[36]),
.ODF(vrtovaj[37]),
.ODG(vrtovaj[38]),
.ODH(vrtovaj[39]),
.OEA(vrtovak[32]),
.OEB(vrtovak[33]),
.OEC(vrtovak[34]),
.OED(vrtovak[35]),
.OEE(vrtovak[36]),
.OEF(vrtovak[37]),
.OEG(vrtovak[38]),
.OEH(vrtovak[39]),
.OFA(vrtovb[32]),
.OFB(vrtovb[33]),
.OFC(vrtovb[34]),
.OFD(vrtovb[35]),
.OFE(vrtovb[36]),
.OFF(vrtovb[37]),
.OFG(vrtovb[38]),
.OFH(vrtovb[39]),
.OGA(scaljtovl[32]),
.OGB(scaljtovl[33]),
.OGC(scaljtovl[34]),
.OGD(scaljtovl[35]),
.OGE(scaljtovl[36]),
.OGF(scaljtovl[37]),
.OGG(scaljtovl[38]),
.OGH(scaljtovl[39]),
.OHA(vrtovlk[32]),
.OHB(vrtovlk[33]),
.OHC(vrtovlk[34]),
.OHD(vrtovlk[35]),
.OHE(vrtovlk[36]),
.OHF(vrtovlk[37]),
.OHG(vrtovlk[38]),
.OHH(vrtovlk[39]),
.OIA(vrtofaj[32]),
.OIB(vrtofaj[33]),
.OIC(vrtofaj[34]),
.OID(vrtofaj[35]),
.OIE(vrtofaj[36]),
.OIF(vrtofaj[37]),
.OIG(vrtofaj[38]),
.OIH(vrtofaj[39]),
.OJA(vrtofak[32]),
.OJB(vrtofak[33]),
.OJC(vrtofak[34]),
.OJD(vrtofak[35]),
.OJE(vrtofak[36]),
.OJF(vrtofak[37]),
.OJG(vrtofak[38]),
.OJH(vrtofak[39]),
.OKA(vrtomulj[32]),
.OKB(vrtomulj[33]),
.OKC(vrtomulj[34]),
.OKD(vrtomulj[35]),
.OKE(vrtomulj[36]),
.OKF(vrtomulj[37]),
.OKG(vrtomulj[38]),
.OKH(vrtomulj[39]),
.OLA(vrtomulk[32]),
.OLB(vrtomulk[33]),
.OLC(vrtomulk[34]),
.OLD(vrtomulk[35]),
.OLE(vrtomulk[36]),
.OLF(vrtomulk[37]),
.OLG(vrtomulk[38]),
.OLH(vrtomulk[39]),
.OMA(vrtolm[32]),
.OMB(vrtolm[33]),
.OMC(vrtolm[34]),
.OMD(vrtolm[35]),
.OME(vrtolm[36]),
.OMF(vrtolm[37]),
.OMG(vrtolm[38]),
.OMH(vrtolm[39]),
.ONA(),
.ONB(),
.ONC(),
.OND(),
.ONE(),
.ONF(),
.ONG(),
.ONH(),
.OOA(vrtocm[32]),
.OOB(vrtocm[33]),
.OOC(vrtocm[34]),
.OOD(vrtocm[35]),
.OOE(vrtocm[36]),
.OOF(vrtocm[37]),
.OOG(vrtocm[38]),
.OOH(vrtocm[39]),
.OQA(sregbrdata[4]),
.OQB(),
.ORA(lmparityeafrvr[4]));



vr vr5 ( 
.IAA(v0addr6[0]),
.IAB(v0addr6[1]),
.IAC(v0addr6[2]),
.IAD(v0addr6[3]),
.IAE(v0addr6[4]),
.IAF(v0addr6[5]),
.IAG(v0vectmode[5]),
.IAH(v0vectstep[5]),
.IBA(v1addr6[0]),
.IBB(v1addr6[1]),
.IBC(v1addr6[2]),
.IBD(v1addr6[3]),
.IBE(v1addr6[4]),
.IBF(v1addr6[5]),
.IBG(v1vectmode[5]),
.IBH(v1vectstep[5]),
.ICA(v2addr6[0]),
.ICB(v2addr6[1]),
.ICC(v2addr6[2]),
.ICD(v2addr6[3]),
.ICE(v2addr6[4]),
.ICF(v2addr6[5]),
.ICG(v2vectmode[5]),
.ICH(v2vectstep[5]),
.IDA(v3addr6[0]),
.IDB(v3addr6[1]),
.IDC(v3addr6[2]),
.IDD(v3addr6[3]),
.IDE(v3addr6[4]),
.IDF(v3addr6[5]),
.IDG(v3vectmode[5]),
.IDH(v3vectstep[5]),
.IEA(v4addr6[0]),
.IEB(v4addr6[1]),
.IEC(v4addr6[2]),
.IED(v4addr6[3]),
.IEE(v4addr6[4]),
.IEF(v4addr6[5]),
.IEG(v4vectmode[5]),
.IEH(v4vectstep[5]),
.IFA(v5addr6[0]),
.IFB(v5addr6[1]),
.IFC(v5addr6[2]),
.IFD(v5addr6[3]),
.IFE(v5addr6[4]),
.IFFF(v5addr6[5]),
.IFG(v5vectmode[5]),
.IFH(v5vectstep[5]),
.IGA(v6addr6[0]),
.IGB(v6addr6[1]),
.IGC(v6addr6[2]),
.IGD(v6addr6[3]),
.IGE(v6addr6[4]),
.IGF(v6addr6[5]),
.IGG(v6vectmode[5]),
.IGH(v6vectstep[5]),
.IHA(v7addr6[0]),
.IHB(v7addr6[1]),
.IHC(v7addr6[2]),
.IHD(v7addr6[3]),
.IHE(v7addr6[4]),
.IHF(v7addr6[5]),
.IHG(v7vectmode[5]),
.IHH(v7vectstep[5]),
.IIA(gatovr[40]),
.IIB(gatovr[41]),
.IIC(gatovr[42]),
.IID(gatovr[43]),
.IIE(gatovr[44]),
.IIF(gatovr[45]),
.IIG(gatovr[46]),
.IIH(gatovr[47]),
.IJA(gbtovr[40]),
.IJB(gbtovr[41]),
.IJC(gbtovr[42]),
.IJD(gbtovr[43]),
.IJE(gbtovr[44]),
.IJF(gbtovr[45]),
.IJG(gbtovr[46]),
.IJH(gbtovr[47]),
.IKA(vbtovr[40]),
.IKB(vbtovr[41]),
.IKC(vbtovr[42]),
.IKD(vbtovr[43]),
.IKE(vbtovr[44]),
.IKF(vbtovr[45]),
.IKG(vbtovr[46]),
.IKH(vbtovr[47]),
.IMA(vltovr[40]),
.IMB(vltovr[41]),
.IMC(vltovr[42]),
.IMD(vltovr[43]),
.IME(vltovr[44]),
.IMF(vltovr[45]),
.IMG(vltovr[46]),
.IMH(vltovr[47]),
.INA(fctovr[40]),
.INB(fctovr[41]),
.INC(fctovr[42]),
.IND(fctovr[43]),
.INE(fctovr[44]),
.INF(fctovr[45]),
.ING(fctovr[46]),
.INH(fctovr[47]),
.IOA(metovr[40]),
.IOB(metovr[41]),
.IOC(metovr[42]),
.IOD(metovr[43]),
.IOE(metovr[44]),
.IOF(metovr[45]),
.IOG(metovr[46]),
.IOH(metovr[47]),
.IPA(watovr[40]),
.IPB(watovr[41]),
.IPC(watovr[42]),
.IPD(watovr[43]),
.IPE(watovr[44]),
.IPF(watovr[45]),
.IPG(watovr[46]),
.IPH(watovr[47]),
.IQA(commemtovr[40]),
.IQB(commemtovr[41]),
.IQC(commemtovr[42]),
.IQD(commemtovr[43]),
.IQE(commemtovr[44]),
.IQF(commemtovr[45]),
.IQG(commemtovr[46]),
.IQH(commemtovr[47]),
.IRA(jbtovr[40]),
.IRB(jbtovr[41]),
.IRC(jbtovr[42]),
.IRD(jbtovr[43]),
.IRE(jbtovr[44]),
.IRF(jbtovr[45]),
.IRG(jbtovr[46]),
.IRH(jbtovr[47]),
.ISA(vector6srccode[0]),
.ISB(vector6srccode[1]),
.ISC(vector6srccode[2]),
.ISD(vector6srccode[3]),
.ISE(vector6srccode[4]),
.ISF(vector6srccode[5]),
.ISG(vector6srccode[6]),
.ITA(scaldesttovr5[0]),
.ITB(scaldesttovr5[1]),
.ITC(scaldesttovr5[2]),
.ITD(scaldesttovr5[3]),
.ITE(scaldesttovr5[4]),
.ITF(scaldesttovr5[5]),
.IZZ (sysclock),
.IZH (ihold),
.OAA(scdatatoga[40]),
.OAB(scdatatoga[41]),
.OAC(scdatatoga[42]),
.OAD(scdatatoga[43]),
.OAE(scdatatoga[44]),
.OAF(scdatatoga[45]),
.OAG(scdatatoga[46]),
.OAH(scdatatoga[47]),
.OBA(shdatatogb[40]),
.OBB(shdatatogb[41]),
.OBC(shdatatogb[42]),
.OBD(shdatatogb[43]),
.OBE(shdatatogb[44]),
.OBF(shdatatogb[45]),
.OBG(shdatatogb[46]),
.OBH(shdatatogb[47]),
.OCA(),
.OCB(),
.OCC(),
.OCD(),
.OCE(),
.OCF(),
.OCG(),
.OCH(),
.ODA(vrtovaj[40]),
.ODB(vrtovaj[41]),
.ODC(vrtovaj[42]),
.ODD(vrtovaj[43]),
.ODE(vrtovaj[44]),
.ODF(vrtovaj[45]),
.ODG(vrtovaj[46]),
.ODH(vrtovaj[47]),
.OEA(vrtovak[40]),
.OEB(vrtovak[41]),
.OEC(vrtovak[42]),
.OED(vrtovak[43]),
.OEE(vrtovak[44]),
.OEF(vrtovak[45]),
.OEG(vrtovak[46]),
.OEH(vrtovak[47]),
.OFA(vrtovb[40]),
.OFB(vrtovb[41]),
.OFC(vrtovb[42]),
.OFD(vrtovb[43]),
.OFE(vrtovb[44]),
.OFF(vrtovb[45]),
.OFG(vrtovb[46]),
.OFH(vrtovb[47]),
.OGA(scaljtovl[40]),
.OGB(scaljtovl[41]),
.OGC(scaljtovl[42]),
.OGD(scaljtovl[43]),
.OGE(scaljtovl[44]),
.OGF(scaljtovl[45]),
.OGG(scaljtovl[46]),
.OGH(scaljtovl[47]),
.OHA(vrtovlk[40]),
.OHB(vrtovlk[41]),
.OHC(vrtovlk[42]),
.OHD(vrtovlk[43]),
.OHE(vrtovlk[44]),
.OHF(vrtovlk[45]),
.OHG(vrtovlk[46]),
.OHH(vrtovlk[47]),
.OIA(vrtofaj[40]),
.OIB(vrtofaj[41]),
.OIC(vrtofaj[42]),
.OID(vrtofaj[43]),
.OIE(vrtofaj[44]),
.OIF(vrtofaj[45]),
.OIG(vrtofaj[46]),
.OIH(vrtofaj[47]),
.OJA(vrtofak[40]),
.OJB(vrtofak[41]),
.OJC(vrtofak[42]),
.OJD(vrtofak[43]),
.OJE(vrtofak[44]),
.OJF(vrtofak[45]),
.OJG(vrtofak[46]),
.OJH(vrtofak[47]),
.OKA(vrtomulj[40]),
.OKB(vrtomulj[41]),
.OKC(vrtomulj[42]),
.OKD(vrtomulj[43]),
.OKE(vrtomulj[44]),
.OKF(vrtomulj[45]),
.OKG(vrtomulj[46]),
.OKH(vrtomulj[47]),
.OLA(vrtomulk[40]),
.OLB(vrtomulk[41]),
.OLC(vrtomulk[42]),
.OLD(vrtomulk[43]),
.OLE(vrtomulk[44]),
.OLF(vrtomulk[45]),
.OLG(vrtomulk[46]),
.OLH(vrtomulk[47]),
.OMA(vrtolm[40]),
.OMB(vrtolm[41]),
.OMC(vrtolm[42]),
.OMD(vrtolm[43]),
.OME(vrtolm[44]),
.OMF(vrtolm[45]),
.OMG(vrtolm[46]),
.OMH(vrtolm[47]),
.ONA(),
.ONB(),
.ONC(),
.OND(),
.ONE(),
.ONF(),
.ONG(),
.ONH(),
.OOA(vrtocm[40]),
.OOB(vrtocm[41]),
.OOC(vrtocm[42]),
.OOD(vrtocm[43]),
.OOE(vrtocm[44]),
.OOF(vrtocm[45]),
.OOG(vrtocm[46]),
.OOH(vrtocm[47]),
.OQA(sregbrdata[5]),
.OQB(),
.ORA(lmparityeafrvr[5]));



vr vr6 ( 
.IAA(v0addr7[0]),
.IAB(v0addr7[1]),
.IAC(v0addr7[2]),
.IAD(v0addr7[3]),
.IAE(v0addr7[4]),
.IAF(v0addr7[5]),
.IAG(v0vectmode[6]),
.IAH(v0vectstep[6]),
.IBA(v1addr7[0]),
.IBB(v1addr7[1]),
.IBC(v1addr7[2]),
.IBD(v1addr7[3]),
.IBE(v1addr7[4]),
.IBF(v1addr7[5]),
.IBG(v1vectmode[6]),
.IBH(v1vectstep[6]),
.ICA(v2addr7[0]),
.ICB(v2addr7[1]),
.ICC(v2addr7[2]),
.ICD(v2addr7[3]),
.ICE(v2addr7[4]),
.ICF(v2addr7[5]),
.ICG(v2vectmode[6]),
.ICH(v2vectstep[6]),
.IDA(v3addr7[0]),
.IDB(v3addr7[1]),
.IDC(v3addr7[2]),
.IDD(v3addr7[3]),
.IDE(v3addr7[4]),
.IDF(v3addr7[5]),
.IDG(v3vectmode[6]),
.IDH(v3vectstep[6]),
.IEA(v4addr7[0]),
.IEB(v4addr7[1]),
.IEC(v4addr7[2]),
.IED(v4addr7[3]),
.IEE(v4addr7[4]),
.IEF(v4addr7[5]),
.IEG(v4vectmode[6]),
.IEH(v4vectstep[6]),
.IFA(v5addr7[0]),
.IFB(v5addr7[1]),
.IFC(v5addr7[2]),
.IFD(v5addr7[3]),
.IFE(v5addr7[4]),
.IFFF(v5addr7[5]),
.IFG(v5vectmode[6]),
.IFH(v5vectstep[6]),
.IGA(v6addr7[0]),
.IGB(v6addr7[1]),
.IGC(v6addr7[2]),
.IGD(v6addr7[3]),
.IGE(v6addr7[4]),
.IGF(v6addr7[5]),
.IGG(v6vectmode[6]),
.IGH(v6vectstep[6]),
.IHA(v7addr7[0]),
.IHB(v7addr7[1]),
.IHC(v7addr7[2]),
.IHD(v7addr7[3]),
.IHE(v7addr7[4]),
.IHF(v7addr7[5]),
.IHG(v7vectmode[6]),
.IHH(v7vectstep[6]),
.IIA(gatovr[48]),
.IIB(gatovr[49]),
.IIC(gatovr[50]),
.IID(gatovr[51]),
.IIE(gatovr[52]),
.IIF(gatovr[53]),
.IIG(gatovr[54]),
.IIH(gatovr[55]),
.IJA(gbtovr[48]),
.IJB(gbtovr[49]),
.IJC(gbtovr[50]),
.IJD(gbtovr[51]),
.IJE(gbtovr[52]),
.IJF(gbtovr[53]),
.IJG(gbtovr[54]),
.IJH(gbtovr[55]),
.IKA(vbtovr[48]),
.IKB(vbtovr[49]),
.IKC(vbtovr[50]),
.IKD(vbtovr[51]),
.IKE(vbtovr[52]),
.IKF(vbtovr[53]),
.IKG(vbtovr[54]),
.IKH(vbtovr[55]),
.IMA(vltovr[48]),
.IMB(vltovr[49]),
.IMC(vltovr[50]),
.IMD(vltovr[51]),
.IME(vltovr[52]),
.IMF(vltovr[53]),
.IMG(vltovr[54]),
.IMH(vltovr[55]),
.INA(fctovr[48]),
.INB(fctovr[49]),
.INC(fctovr[50]),
.IND(fctovr[51]),
.INE(fctovr[52]),
.INF(fctovr[53]),
.ING(fctovr[54]),
.INH(fctovr[55]),
.IOA(metovr[48]),
.IOB(metovr[49]),
.IOC(metovr[50]),
.IOD(metovr[51]),
.IOE(metovr[52]),
.IOF(metovr[53]),
.IOG(metovr[54]),
.IOH(metovr[55]),
.IPA(watovr[48]),
.IPB(watovr[49]),
.IPC(watovr[50]),
.IPD(watovr[51]),
.IPE(watovr[52]),
.IPF(watovr[53]),
.IPG(watovr[54]),
.IPH(watovr[55]),
.IQA(commemtovr[48]),
.IQB(commemtovr[49]),
.IQC(commemtovr[50]),
.IQD(commemtovr[51]),
.IQE(commemtovr[52]),
.IQF(commemtovr[53]),
.IQG(commemtovr[54]),
.IQH(commemtovr[55]),
.IRA(jbtovr[48]),
.IRB(jbtovr[49]),
.IRC(jbtovr[50]),
.IRD(jbtovr[51]),
.IRE(jbtovr[52]),
.IRF(jbtovr[53]),
.IRG(jbtovr[54]),
.IRH(jbtovr[55]),
.ISA(vector7srccode[0]),
.ISB(vector7srccode[1]),
.ISC(vector7srccode[2]),
.ISD(vector7srccode[3]),
.ISE(vector7srccode[4]),
.ISF(vector7srccode[5]),
.ISG(vector7srccode[6]),
.ITA(scaldesttovr6[0]),
.ITB(scaldesttovr6[1]),
.ITC(scaldesttovr6[2]),
.ITD(scaldesttovr6[3]),
.ITE(scaldesttovr6[4]),
.ITF(scaldesttovr6[5]),
.IZZ (sysclock),
.IZH (ihold),
.OAA(scdatatoga[48]),
.OAB(scdatatoga[49]),
.OAC(scdatatoga[50]),
.OAD(scdatatoga[51]),
.OAE(scdatatoga[52]),
.OAF(scdatatoga[53]),
.OAG(scdatatoga[54]),
.OAH(scdatatoga[55]),
.OBA(shdatatogb[48]),
.OBB(shdatatogb[49]),
.OBC(shdatatogb[50]),
.OBD(shdatatogb[51]),
.OBE(shdatatogb[52]),
.OBF(shdatatogb[53]),
.OBG(shdatatogb[54]),
.OBH(shdatatogb[55]),
.OCA(),
.OCB(),
.OCC(),
.OCD(),
.OCE(),
.OCF(),
.OCG(),
.OCH(),
.ODA(vrtovaj[48]),
.ODB(vrtovaj[49]),
.ODC(vrtovaj[50]),
.ODD(vrtovaj[51]),
.ODE(vrtovaj[52]),
.ODF(vrtovaj[53]),
.ODG(vrtovaj[54]),
.ODH(vrtovaj[55]),
.OEA(vrtovak[48]),
.OEB(vrtovak[49]),
.OEC(vrtovak[50]),
.OED(vrtovak[51]),
.OEE(vrtovak[52]),
.OEF(vrtovak[53]),
.OEG(vrtovak[54]),
.OEH(vrtovak[55]),
.OFA(vrtovb[48]),
.OFB(vrtovb[49]),
.OFC(vrtovb[50]),
.OFD(vrtovb[51]),
.OFE(vrtovb[52]),
.OFF(vrtovb[53]),
.OFG(vrtovb[54]),
.OFH(vrtovb[55]),
.OGA(scaljtovl[48]),
.OGB(scaljtovl[49]),
.OGC(scaljtovl[50]),
.OGD(scaljtovl[51]),
.OGE(scaljtovl[52]),
.OGF(scaljtovl[53]),
.OGG(scaljtovl[54]),
.OGH(scaljtovl[55]),
.OHA(vrtovlk[48]),
.OHB(vrtovlk[49]),
.OHC(vrtovlk[50]),
.OHD(vrtovlk[51]),
.OHE(vrtovlk[52]),
.OHF(vrtovlk[53]),
.OHG(vrtovlk[54]),
.OHH(vrtovlk[55]),
.OIA(vrtofaj[48]),
.OIB(vrtofaj[49]),
.OIC(vrtofaj[50]),
.OID(vrtofaj[51]),
.OIE(vrtofaj[52]),
.OIF(vrtofaj[53]),
.OIG(vrtofaj[54]),
.OIH(vrtofaj[55]),
.OJA(vrtofak[48]),
.OJB(vrtofak[49]),
.OJC(vrtofak[50]),
.OJD(vrtofak[51]),
.OJE(vrtofak[52]),
.OJF(vrtofak[53]),
.OJG(vrtofak[54]),
.OJH(vrtofak[55]),
.OKA(vrtomulj[48]),
.OKB(vrtomulj[49]),
.OKC(vrtomulj[50]),
.OKD(vrtomulj[51]),
.OKE(vrtomulj[52]),
.OKF(vrtomulj[53]),
.OKG(vrtomulj[54]),
.OKH(vrtomulj[55]),
.OLA(vrtomulk[48]),
.OLB(vrtomulk[49]),
.OLC(vrtomulk[50]),
.OLD(vrtomulk[51]),
.OLE(vrtomulk[52]),
.OLF(vrtomulk[53]),
.OLG(vrtomulk[54]),
.OLH(vrtomulk[55]),
.OMA(vrtolm[48]),
.OMB(vrtolm[49]),
.OMC(vrtolm[50]),
.OMD(vrtolm[51]),
.OME(vrtolm[52]),
.OMF(vrtolm[53]),
.OMG(vrtolm[54]),
.OMH(vrtolm[55]),
.ONA(),
.ONB(),
.ONC(),
.OND(),
.ONE(),
.ONF(),
.ONG(),
.ONH(),
.OOA(vrtocm[48]),
.OOB(vrtocm[49]),
.OOC(vrtocm[50]),
.OOD(vrtocm[51]),
.OOE(vrtocm[52]),
.OOF(vrtocm[53]),
.OOG(vrtocm[54]),
.OOH(vrtocm[55]),
.OQA(sregbrdata[6]),
.OQB(),
.ORA(lmparityeafrvr[6]));



vr vr7 ( 
.IAA(v0addr8[0]),
.IAB(v0addr8[1]),
.IAC(v0addr8[2]),
.IAD(v0addr8[3]),
.IAE(v0addr8[4]),
.IAF(v0addr8[5]),
.IAG(v0vectmode[7]),
.IAH(v0vectstep[7]),
.IBA(v1addr8[0]),
.IBB(v1addr8[1]),
.IBC(v1addr8[2]),
.IBD(v1addr8[3]),
.IBE(v1addr8[4]),
.IBF(v1addr8[5]),
.IBG(v1vectmode[7]),
.IBH(v1vectstep[7]),
.ICA(v2addr8[0]),
.ICB(v2addr8[1]),
.ICC(v2addr8[2]),
.ICD(v2addr8[3]),
.ICE(v2addr8[4]),
.ICF(v2addr8[5]),
.ICG(v2vectmode[7]),
.ICH(v2vectstep[7]),
.IDA(v3addr8[0]),
.IDB(v3addr8[1]),
.IDC(v3addr8[2]),
.IDD(v3addr8[3]),
.IDE(v3addr8[4]),
.IDF(v3addr8[5]),
.IDG(v3vectmode[7]),
.IDH(v3vectstep[7]),
.IEA(v4addr8[0]),
.IEB(v4addr8[1]),
.IEC(v4addr8[2]),
.IED(v4addr8[3]),
.IEE(v4addr8[4]),
.IEF(v4addr8[5]),
.IEG(v4vectmode[7]),
.IEH(v4vectstep[7]),
.IFA(v5addr8[0]),
.IFB(v5addr8[1]),
.IFC(v5addr8[2]),
.IFD(v5addr8[3]),
.IFE(v5addr8[4]),
.IFFF(v5addr8[5]),
.IFG(v5vectmode[7]),
.IFH(v5vectstep[7]),
.IGA(v6addr8[0]),
.IGB(v6addr8[1]),
.IGC(v6addr8[2]),
.IGD(v6addr8[3]),
.IGE(v6addr8[4]),
.IGF(v6addr8[5]),
.IGG(v6vectmode[7]),
.IGH(v6vectstep[7]),
.IHA(v7addr8[0]),
.IHB(v7addr8[1]),
.IHC(v7addr8[2]),
.IHD(v7addr8[3]),
.IHE(v7addr8[4]),
.IHF(v7addr8[5]),
.IHG(v7vectmode[7]),
.IHH(v7vectstep[7]),
.IIA(gatovr[56]),
.IIB(gatovr[57]),
.IIC(gatovr[58]),
.IID(gatovr[59]),
.IIE(gatovr[60]),
.IIF(gatovr[61]),
.IIG(gatovr[62]),
.IIH(gatovr[63]),
.IJA(gbtovr[56]),
.IJB(gbtovr[57]),
.IJC(gbtovr[58]),
.IJD(gbtovr[59]),
.IJE(gbtovr[60]),
.IJF(gbtovr[61]),
.IJG(gbtovr[62]),
.IJH(gbtovr[63]),
.IKA(vbtovr[56]),
.IKB(vbtovr[57]),
.IKC(vbtovr[58]),
.IKD(vbtovr[59]),
.IKE(vbtovr[60]),
.IKF(vbtovr[61]),
.IKG(vbtovr[62]),
.IKH(vbtovr[63]),
.IMA(vltovr[56]),
.IMB(vltovr[57]),
.IMC(vltovr[58]),
.IMD(vltovr[59]),
.IME(vltovr[60]),
.IMF(vltovr[61]),
.IMG(vltovr[62]),
.IMH(vltovr[63]),
.INA(fctovr[56]),
.INB(fctovr[57]),
.INC(fctovr[58]),
.IND(fctovr[59]),
.INE(fctovr[60]),
.INF(fctovr[61]),
.ING(fctovr[62]),
.INH(fctovr[63]),
.IOA(metovr[56]),
.IOB(metovr[57]),
.IOC(metovr[58]),
.IOD(metovr[59]),
.IOE(metovr[60]),
.IOF(metovr[61]),
.IOG(metovr[62]),
.IOH(metovr[63]),
.IPA(watovr[56]),
.IPB(watovr[57]),
.IPC(watovr[58]),
.IPD(watovr[59]),
.IPE(watovr[60]),
.IPF(watovr[61]),
.IPG(watovr[62]),
.IPH(watovr[63]),
.IQA(commemtovr[56]),
.IQB(commemtovr[57]),
.IQC(commemtovr[58]),
.IQD(commemtovr[59]),
.IQE(commemtovr[60]),
.IQF(commemtovr[61]),
.IQG(commemtovr[62]),
.IQH(commemtovr[63]),
.IRA(jbtovr[56]),
.IRB(jbtovr[57]),
.IRC(jbtovr[58]),
.IRD(jbtovr[59]),
.IRE(jbtovr[60]),
.IRF(jbtovr[61]),
.IRG(jbtovr[62]),
.IRH(jbtovr[63]),
.ISA(vector8srccode[0]),
.ISB(vector8srccode[1]),
.ISC(vector8srccode[2]),
.ISD(vector8srccode[3]),
.ISE(vector8srccode[4]),
.ISF(vector8srccode[5]),
.ISG(vector8srccode[6]),
.ITA(scaldesttovr7[0]),
.ITB(scaldesttovr7[1]),
.ITC(scaldesttovr7[2]),
.ITD(scaldesttovr7[3]),
.ITE(scaldesttovr7[4]),
.ITF(scaldesttovr7[5]),
.IZZ (sysclock),
.IZH (ihold),
.OAA(scdatatoga[56]),
.OAB(scdatatoga[57]),
.OAC(scdatatoga[58]),
.OAD(scdatatoga[59]),
.OAE(scdatatoga[60]),
.OAF(scdatatoga[61]),
.OAG(scdatatoga[62]),
.OAH(scdatatoga[63]),
.OBA(shdatatogb[56]),
.OBB(shdatatogb[57]),
.OBC(shdatatogb[58]),
.OBD(shdatatogb[59]),
.OBE(shdatatogb[60]),
.OBF(shdatatogb[61]),
.OBG(shdatatogb[62]),
.OBH(shdatatogb[63]),
.OCA(),
.OCB(),
.OCC(),
.OCD(),
.OCE(),
.OCF(),
.OCG(),
.OCH(),
.ODA(vrtovaj[56]),
.ODB(vrtovaj[57]),
.ODC(vrtovaj[58]),
.ODD(vrtovaj[59]),
.ODE(vrtovaj[60]),
.ODF(vrtovaj[61]),
.ODG(vrtovaj[62]),
.ODH(vrtovaj[63]),
.OEA(vrtovak[56]),
.OEB(vrtovak[57]),
.OEC(vrtovak[58]),
.OED(vrtovak[59]),
.OEE(vrtovak[60]),
.OEF(vrtovak[61]),
.OEG(vrtovak[62]),
.OEH(vrtovak[63]),
.OFA(vrtovb[56]),
.OFB(vrtovb[57]),
.OFC(vrtovb[58]),
.OFD(vrtovb[59]),
.OFE(vrtovb[60]),
.OFF(vrtovb[61]),
.OFG(vrtovb[62]),
.OFH(vrtovb[63]),
.OGA(scaljtovl[56]),
.OGB(scaljtovl[57]),
.OGC(scaljtovl[58]),
.OGD(scaljtovl[59]),
.OGE(scaljtovl[60]),
.OGF(scaljtovl[61]),
.OGG(scaljtovl[62]),
.OGH(scaljtovl[63]),
.OHA(vrtovlk[56]),
.OHB(vrtovlk[57]),
.OHC(vrtovlk[58]),
.OHD(vrtovlk[59]),
.OHE(vrtovlk[60]),
.OHF(vrtovlk[61]),
.OHG(vrtovlk[62]),
.OHH(vrtovlk[63]),
.OIA(vrtofaj[56]),
.OIB(vrtofaj[57]),
.OIC(vrtofaj[58]),
.OID(vrtofaj[59]),
.OIE(vrtofaj[60]),
.OIF(vrtofaj[61]),
.OIG(vrtofaj[62]),
.OIH(vrtofaj[63]),
.OJA(vrtofak[56]),
.OJB(vrtofak[57]),
.OJC(vrtofak[58]),
.OJD(vrtofak[59]),
.OJE(vrtofak[60]),
.OJF(vrtofak[61]),
.OJG(vrtofak[62]),
.OJH(vrtofak[63]),
.OKA(vrtomulj[56]),
.OKB(vrtomulj[57]),
.OKC(vrtomulj[58]),
.OKD(vrtomulj[59]),
.OKE(vrtomulj[60]),
.OKF(vrtomulj[61]),
.OKG(vrtomulj[62]),
.OKH(vrtomulj[63]),
.OLA(vrtomulk[56]),
.OLB(vrtomulk[57]),
.OLC(vrtomulk[58]),
.OLD(vrtomulk[59]),
.OLE(vrtomulk[60]),
.OLF(vrtomulk[61]),
.OLG(vrtomulk[62]),
.OLH(vrtomulk[63]),
.OMA(vrtolm[56]),
.OMB(vrtolm[57]),
.OMC(vrtolm[58]),
.OMD(vrtolm[59]),
.OME(vrtolm[60]),
.OMF(vrtolm[61]),
.OMG(vrtolm[62]),
.OMH(vrtolm[63]),
.ONA(),
.ONB(),
.ONC(),
.OND(),
.ONE(),
.ONF(),
.ONG(),
.ONH(),
.OOA(vrtocm[56]),
.OOB(vrtocm[57]),
.OOC(vrtocm[58]),
.OOD(vrtocm[59]),
.OOE(vrtocm[60]),
.OOF(vrtocm[61]),
.OOG(vrtocm[62]),
.OOH(vrtocm[63]),
.OQA(sregbrdata[7]),
.OQB(vasregsign),
.ORA(lmparityeafrvr[7]));


wa wa0 ( 
.IAA(vrtolm[0]),
.IAB(vrtolm[1]),
.IAC(vrtolm[2]),
.IAD(vrtolm[3]),
.IAE(vrtolm[4]),
.IAF(vrtolm[5]),
.IAG(vrtolm[6]),
.IAH(vrtolm[7]),
.IAI(vrtolm[8]),
.IAJ(vrtolm[9]),
.IAK(vrtolm[10]),
.IAL(vrtolm[11]),
.IAM(vrtolm[12]),
.IAN(vrtolm[13]),
.IAO(vrtolm[14]),
.IAP(vrtolm[15]),
.IBA(vrtolm[16]),
.IBB(vrtolm[17]),
.IBC(vrtolm[18]),
.IBD(vrtolm[19]),
.IBE(vrtolm[20]),
.IBF(vrtolm[21]),
.IBG(vrtolm[22]),
.IBH(vrtolm[23]),
.IBI(vrtolm[24]),
.IBJ(vrtolm[25]),
.IBK(vrtolm[26]),
.IBL(vrtolm[27]),
.IBM(vrtolm[28]),
.IBN(vrtolm[29]),
.IBO(vrtolm[30]),
.IBP(vrtolm[31]),
.ICA(vrtolm[32]),
.ICB(vrtolm[33]),
.ICC(vrtolm[34]),
.ICD(vrtolm[35]),
.ICE(vrtolm[36]),
.ICF(vrtolm[37]),
.ICG(vrtolm[38]),
.ICH(vrtolm[39]),
.ICI(vrtolm[40]),
.ICJ(vrtolm[41]),
.ICK(vrtolm[42]),
.ICL(vrtolm[43]),
.ICM(vrtolm[44]),
.ICN(vrtolm[45]),
.ICO(vrtolm[46]),
.ICP(vrtolm[47]),
.IDA(vrtolm[48]),
.IDB(vrtolm[49]),
.IDC(vrtolm[50]),
.IDD(vrtolm[51]),
.IDE(vrtolm[52]),
.IDF(vrtolm[53]),
.IDG(vrtolm[54]),
.IDH(vrtolm[55]),
.IDI(vrtolm[56]),
.IDJ(vrtolm[57]),
.IDK(vrtolm[58]),
.IDL(vrtolm[59]),
.IDM(vrtolm[60]),
.IDN(vrtolm[61]),
.IDO(vrtolm[62]),
.IDP(vrtolm[63]),
.IEA(wadatalm[0]),
.IEB(wadatalm[1]),
.IEC(wadatalm[2]),
.IED(wadatalm[3]),
.IEE(wadatalm[4]),
.IEF(wadatalm[5]),
.IEG(wadatalm[6]),
.IEH(wadatalm[7]),
.IEI(wadatalm[8]),
.IEJ(wadatalm[9]),
.IEK(wadatalm[10]),
.IEL(wadatalm[11]),
.IEM(wadatalm[12]),
.IEN(wadatalm[13]),
.IEO(wadatalm[14]),
.IEP(wadatalm[15]),
.IFA(wadatalm[16]),
.IFB(wadatalm[17]),
.IFC(wadatalm[18]),
.IFD(wadatalm[19]),
.IFE(wadatalm[20]),
.IFFF(wadatalm[21]),
.IFG(wadatalm[22]),
.IFH(wadatalm[23]),
.IFI(wadatalm[24]),
.IFJ(wadatalm[25]),
.IFK(wadatalm[26]),
.IFL(wadatalm[27]),
.IFM(wadatalm[28]),
.IFN(wadatalm[29]),
.IFO(wadatalm[30]),
.IFP(wadatalm[31]),
.IGA(parceltowa[0]),
.IGB(parceltowa[1]),
.IGC(parceltowa[2]),
.IGD(parceltowa[3]),
.IGE(parceltowa[4]),
.IGF(parceltowa[5]),
.IGG(parceltowa[6]),
.IGH(parceltowa[7]),
.IGI(parceltowa[8]),
.IGJ(parceltowa[9]),
.IGK(parceltowa[10]),
.IGL(parceltowa[11]),
.IGM(parceltowa[12]),
.IGN(parceltowa[13]),
.IGO(parceltowa[14]),
.IGP(parceltowa[15]),
.IHA(goissuetowa[0]),
.IHB(goissuetowa[1]),
.IIA(constreadwa),
.IIB(constwritewa),
.IJA(enteradtowa),
.IJB(entervrtowa),
.IJC(enterardtowa),
.IJD(advlmadrtowa),
.IKA(jamecnt[0]),
.IKB(jamecnt[1]),
.IKC(jamecnt[2]),
.IKD(jamecnt[3]),
.IKE(jamecnt[4]),
.IKF(jamecnt[5]),
.IZZ (sysclock),
.OAA(watovr[0]),
.OAB(watovr[1]),
.OAC(watovr[2]),
.OAD(watovr[3]),
.OAE(watovr[4]),
.OAF(watovr[5]),
.OAG(watovr[6]),
.OAH(watovr[7]),
.OAI(watovr[8]),
.OAJ(watovr[9]),
.OAK(watovr[10]),
.OAL(watovr[11]),
.OAM(watovr[12]),
.OAN(watovr[13]),
.OAO(watovr[14]),
.OAP(watovr[15]),
.OBA(watovr[16]),
.OBB(watovr[17]),
.OBC(watovr[18]),
.OBD(watovr[19]),
.OBE(watovr[20]),
.OBF(watovr[21]),
.OBG(watovr[22]),
.OBH(watovr[23]),
.OBI(watovr[24]),
.OBJ(watovr[25]),
.OBK(watovr[26]),
.OBL(watovr[27]),
.OBM(watovr[28]),
.OBN(watovr[29]),
.OBO(watovr[30]),
.OBP(watovr[31]),
.OCA(watovr[32]),
.OCB(watovr[33]),
.OCC(watovr[34]),
.OCD(watovr[35]),
.OCE(watovr[36]),
.OCF(watovr[37]),
.OCG(watovr[38]),
.OCH(watovr[39]),
.OCI(watovr[40]),
.OCJ(watovr[41]),
.OCK(watovr[42]),
.OCL(watovr[43]),
.OCM(watovr[44]),
.OCN(watovr[45]),
.OCO(watovr[46]),
.OCP(watovr[47]),
.ODA(watovr[48]),
.ODB(watovr[49]),
.ODC(watovr[50]),
.ODD(watovr[51]),
.ODE(watovr[52]),
.ODF(watovr[53]),
.ODG(watovr[54]),
.ODH(watovr[55]),
.ODI(watovr[56]),
.ODJ(watovr[57]),
.ODK(watovr[58]),
.ODL(watovr[59]),
.ODM(watovr[60]),
.ODN(watovr[61]),
.ODO(watovr[62]),
.ODP(watovr[63]),
.OEA(watoar[0]),
.OEB(watoar[1]),
.OEC(watoar[2]),
.OED(watoar[3]),
.OEE(watoar[4]),
.OEF(watoar[5]),
.OEG(watoar[6]),
.OEH(watoar[7]),
.OEI(watoar[8]),
.OEJ(watoar[9]),
.OEK(watoar[10]),
.OEL(watoar[11]),
.OEM(watoar[12]),
.OEN(watoar[13]),
.OEO(watoar[14]),
.OEP(watoar[15]),
.OFA(watoar[16]),
.OFB(watoar[17]),
.OFC(watoar[18]),
.OFD(watoar[19]),
.OFE(watoar[20]),
.OFF(watoar[21]),
.OFG(watoar[22]),
.OFH(watoar[23]),
.OFI(watoar[24]),
.OFJ(watoar[25]),
.OFK(watoar[26]),
.OFL(watoar[27]),
.OFM(watoar[28]),
.OFN(watoar[29]),
.OFO(watoar[30]),
.OFP(watoar[31]),
.OGA(wajamecnt[0]),
.OGB(wajamecnt[1]),
.OGC(wajamecnt[2]),
.OGD(wajamecnt[3]),
.OGE(wajamecnt[4]),
.OGF(wajamecnt[5]));

   // fakeifs to replace cpu1-3 if modules for semaphore loop
   
fakeif fk1 (
.IZZ(sysclock),
.IAA(semaphorefl_0[0]),
.IAB(semaphorefl_0[0]),
.OAA(semaphorefl_1[0]),
.OAB(semaphorefl_1[0]) );
   

fakeif fk2 (
.IZZ(sysclock),
.IAA(semaphorefl_1[0]),
.IAB(semaphorefl_1[0]),
.OAA(semaphorefl_2[0]),
.OAB(semaphorefl_2[0]) );
   

fakeif fk3 (
.IZZ(sysclock),
.IAA(semaphorefl_2[0]),
.IAB(semaphorefl_2[0]),
.OAA(semaphorefl_3[0]),
.OAB(semaphorefl_3[1]) );
   
            
            
endmodule;
