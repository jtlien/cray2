module va( IZZ,
 IAA, 
 IAB, 
 IAC, 
 IAD, 
 IAE, 
 IAF, 
 IAG, 
 IAH, 
 IAI, 
 IAJ, 
 IAK, 
 IAL, 
 IAM, 
 IAN, 
 IAO, 
 IAP, 
 IBA, 
 IBB, 
 IBC, 
 IBD, 
 IBE, 
 IBF, 
 IBG, 
 IBH, 
 IBI, 
 IBJ, 
 IBK, 
 IBL, 
 IBM, 
 IBN, 
 IBO, 
 IBP, 
 ICA, 
 ICB, 
 ICC, 
 ICD, 
 ICE, 
 ICF, 
 ICG, 
 ICH, 
 ICI, 
 ICJ, 
 ICK, 
 ICL, 
 ICM, 
 ICN, 
 ICO, 
 ICP, 
 IDA, 
 IDB, 
 IDC, 
 IDD, 
 IDE, 
 IDF, 
 IDG, 
 IDH, 
 IDI, 
 IDJ, 
 IDK, 
 IDL, 
 IDM, 
 IDN, 
 IDO, 
 IDP, 
 IEA, 
 IEB, 
 IEC, 
 IED, 
 IEE, 
 IEF, 
 IEG, 
 IEH, 
 IEI, 
 IEJ, 
 IEK, 
 IEL, 
 IEM, 
 IEN, 
 IEO, 
 IEP, 
 IFA, 
 IFB, 
 IFC, 
 IFD, 
 IFE, 
 IFFF , 
 IFG, 
 IFH, 
 IFI, 
 IFJ, 
 IFK, 
 IFL, 
 IFM, 
 IFN, 
 IFO, 
 IFP, 
 IGA, 
 IGB, 
 IGC, 
 IGD, 
 IGE, 
 IGF, 
 IGG, 
 IGH, 
 IGI, 
 IGJ, 
 IGK, 
 IGL, 
 IGM, 
 IGN, 
 IGO, 
 IGP, 
 IHA, 
 IHB, 
 IHC, 
 IHD, 
 IHE, 
 IHF, 
 IHG, 
 IHH, 
 IHI, 
 IHJ, 
 IHK, 
 IHL, 
 IHM, 
 IHN, 
 IHO, 
 IHP, 
 IMA, 
 IRA, 
 IRB, 
 IRC, 
 IRD, 
 OAA, 
 OAB, 
 OAC, 
 OAD, 
 OAE, 
 OAF, 
 OAG, 
 OAH, 
 OAI, 
 OAJ, 
 OAK, 
 OAL, 
 OAM, 
 OAN, 
 OAO, 
 OAP, 
 OBA, 
 OBB, 
 OBC, 
 OBD, 
 OBE, 
 OBF, 
 OBG, 
 OBH, 
 OBI, 
 OBJ, 
 OBK, 
 OBL, 
 OBM, 
 OBN, 
 OBO, 
 OBP, 
 OCA, 
 OCB, 
 OCC, 
 OCD, 
 OCE, 
 OCF, 
 OCG, 
 OCH, 
 OCI, 
 OCJ, 
 OCK, 
 OCL, 
 OCM, 
 OCN, 
 OCO, 
 OCP, 
 ODA, 
 ODB, 
 ODC, 
 ODD, 
 ODE, 
 ODF, 
 ODG, 
 ODH, 
 ODI, 
 ODJ, 
 ODK, 
 ODL, 
 ODM, 
 ODN, 
 ODO, 
 ODP, 
 OEA, 
 OEB, 
 OEC, 
 OFA, 
 OFB, 
ONA ); 
    
 input IZZ; 
 input IAA; 
 input IAB; 
 input IAC; 
 input IAD; 
 input IAE; 
 input IAF; 
 input IAG; 
 input IAH; 
 input IAI; 
 input IAJ; 
 input IAK; 
 input IAL; 
 input IAM; 
 input IAN; 
 input IAO; 
 input IAP; 
 input IBA; 
 input IBB; 
 input IBC; 
 input IBD; 
 input IBE; 
 input IBF; 
 input IBG; 
 input IBH; 
 input IBI; 
 input IBJ; 
 input IBK; 
 input IBL; 
 input IBM; 
 input IBN; 
 input IBO; 
 input IBP; 
 input ICA; 
 input ICB; 
 input ICC; 
 input ICD; 
 input ICE; 
 input ICF; 
 input ICG; 
 input ICH; 
 input ICI; 
 input ICJ; 
 input ICK; 
 input ICL; 
 input ICM; 
 input ICN; 
 input ICO; 
 input ICP; 
 input IDA; 
 input IDB; 
 input IDC; 
 input IDD; 
 input IDE; 
 input IDF; 
 input IDG; 
 input IDH; 
 input IDI; 
 input IDJ; 
 input IDK; 
 input IDL; 
 input IDM; 
 input IDN; 
 input IDO; 
 input IDP; 
 input IEA; 
 input IEB; 
 input IEC; 
 input IED; 
 input IEE; 
 input IEF; 
 input IEG; 
 input IEH; 
 input IEI; 
 input IEJ; 
 input IEK; 
 input IEL; 
 input IEM; 
 input IEN; 
 input IEO; 
 input IEP; 
 input IFA; 
 input IFB; 
 input IFC; 
 input IFD; 
 input IFE; 
 input IFFF ; 
 input IFG; 
 input IFH; 
 input IFI; 
 input IFJ; 
 input IFK; 
 input IFL; 
 input IFM; 
 input IFN; 
 input IFO; 
 input IFP; 
 input IGA; 
 input IGB; 
 input IGC; 
 input IGD; 
 input IGE; 
 input IGF; 
 input IGG; 
 input IGH; 
 input IGI; 
 input IGJ; 
 input IGK; 
 input IGL; 
 input IGM; 
 input IGN; 
 input IGO; 
 input IGP; 
 input IHA; 
 input IHB; 
 input IHC; 
 input IHD; 
 input IHE; 
 input IHF; 
 input IHG; 
 input IHH; 
 input IHI; 
 input IHJ; 
 input IHK; 
 input IHL; 
 input IHM; 
 input IHN; 
 input IHO; 
 input IHP; 
 input IMA; 
 input IRA; 
 input IRB; 
 input IRC; 
 input IRD; 
 output OAA; 
 output OAB; 
 output OAC; 
 output OAD; 
 output OAE; 
 output OAF; 
 output OAG; 
 output OAH; 
 output OAI; 
 output OAJ; 
 output OAK; 
 output OAL; 
 output OAM; 
 output OAN; 
 output OAO; 
 output OAP; 
 output OBA; 
 output OBB; 
 output OBC; 
 output OBD; 
 output OBE; 
 output OBF; 
 output OBG; 
 output OBH; 
 output OBI; 
 output OBJ; 
 output OBK; 
 output OBL; 
 output OBM; 
 output OBN; 
 output OBO; 
 output OBP; 
 output OCA; 
 output OCB; 
 output OCC; 
 output OCD; 
 output OCE; 
 output OCF; 
 output OCG; 
 output OCH; 
 output OCI; 
 output OCJ; 
 output OCK; 
 output OCL; 
 output OCM; 
 output OCN; 
 output OCO; 
 output OCP; 
 output ODA; 
 output ODB; 
 output ODC; 
 output ODD; 
 output ODE; 
 output ODF; 
 output ODG; 
 output ODH; 
 output ODI; 
 output ODJ; 
 output ODK; 
 output ODL; 
 output ODM; 
 output ODN; 
 output ODO; 
 output ODP; 
 output OEA; 
 output OEB; 
 output OEC; 
 output OFA; 
 output OFB; 
 output ONA; 
  
  
reg  aaa ;
reg  aab ;
reg  aac ;
reg  aad ;
reg  aba ;
reg  abb ;
reg  abc ;
reg  abd ;
reg  aca ;
reg  acb ;
reg  acc ;
reg  acd ;
reg  ada ;
reg  adb ;
reg  adc ;
reg  add ;
reg  aea ;
reg  aeb ;
reg  aec ;
reg  aed ;
reg  afa ;
reg  afb ;
reg  afc ;
reg  afd ;
reg  aga ;
reg  agb ;
reg  agc ;
reg  agd ;
reg  aha ;
reg  ahb ;
reg  ahc ;
reg  ahd ;
reg  aia ;
reg  aib ;
reg  aic ;
reg  aid ;
reg  aja ;
reg  ajb ;
reg  ajc ;
reg  ajd ;
reg  aka ;
reg  akb ;
reg  akc ;
reg  akd ;
reg  ala ;
reg  alb ;
reg  alc ;
reg  ald ;
reg  ama ;
reg  amb ;
reg  amc ;
reg  amd ;
reg  ana ;
reg  anb ;
reg  anc ;
reg  andd  ;
reg  aoa ;
reg  aob ;
reg  aoc ;
reg  aod ;
reg  apa ;
reg  apb ;
reg  apc ;
reg  apd ;
reg  BAA ;
reg  BAB ;
reg  BAC ;
reg  BAD ;
reg  BBA ;
reg  BBB ;
reg  BBC ;
reg  BBD ;
reg  BBF ;
reg  BBG ;
reg  BCA ;
reg  BCB ;
reg  BCC ;
reg  BCD ;
reg  BCF ;
reg  BCG ;
reg  BDA ;
reg  BDB ;
reg  BDC ;
reg  BDD ;
reg  BDF ;
reg  BDG ;
reg  BEA ;
reg  BEB ;
reg  BEC ;
reg  BED ;
reg  BEF ;
reg  BEG ;
reg  BFA ;
reg  BFB ;
reg  BFC ;
reg  BFD ;
reg  BFF ;
reg  BFG ;
reg  BGA ;
reg  BGB ;
reg  BGC ;
reg  BGD ;
reg  BGF ;
reg  BGG ;
reg  BHA ;
reg  BHB ;
reg  BHC ;
reg  BHD ;
reg  BHF ;
reg  BHG ;
reg  BIA ;
reg  BIB ;
reg  BIC ;
reg  BID ;
reg  BIF ;
reg  BIG ;
reg  BJA ;
reg  BJB ;
reg  BJC ;
reg  BJD ;
reg  BJF ;
reg  BJG ;
reg  BKA ;
reg  BKB ;
reg  BKC ;
reg  BKD ;
reg  BKF ;
reg  BKG ;
reg  BLA ;
reg  BLB ;
reg  BLC ;
reg  BLD ;
reg  BLF ;
reg  BMA ;
reg  BMB ;
reg  BMC ;
reg  BMD ;
reg  BMF ;
reg  BMG ;
reg  BNA ;
reg  BNB ;
reg  BNC ;
reg  BND ;
reg  BNF ;
reg  BNG ;
reg  BOA ;
reg  BOB ;
reg  BOC ;
reg  BOD ;
reg  BOF ;
reg  BOG ;
reg  BPA ;
reg  BPB ;
reg  BPC ;
reg  BPD ;
reg  dfb ;
reg  gaa ;
reg  gab ;
reg  gac ;
reg  gad ;
reg  gba ;
reg  gbb ;
reg  gbc ;
reg  gbd ;
reg  gca ;
reg  gcb ;
reg  gcc ;
reg  gcd ;
reg  gda ;
reg  gdb ;
reg  gdc ;
reg  gdd ;
reg  gea ;
reg  geb ;
reg  gec ;
reg  ged ;
reg  gfa ;
reg  gfb ;
reg  gfc ;
reg  gfd ;
reg  gga ;
reg  ggb ;
reg  ggc ;
reg  ggd ;
reg  gha ;
reg  ghb ;
reg  ghc ;
reg  ghd ;
reg  gia ;
reg  gib ;
reg  gic ;
reg  gid ;
reg  gja ;
reg  gjb ;
reg  gjc ;
reg  gjd ;
reg  gka ;
reg  gkb ;
reg  gkc ;
reg  gkd ;
reg  gla ;
reg  glb ;
reg  glc ;
reg  gld ;
reg  gma ;
reg  gmb ;
reg  gmc ;
reg  gmd ;
reg  gna ;
reg  gnb ;
reg  gnc ;
reg  gnd ;
reg  goa ;
reg  gob ;
reg  goc ;
reg  god ;
reg  gpa ;
reg  gpb ;
reg  gpc ;
reg  gpd ;
reg  hba ;
reg  hbb ;
reg  hbc ;
reg  hbd ;
reg  hca ;
reg  hcb ;
reg  hcc ;
reg  hcd ;
reg  hda ;
reg  hdb ;
reg  hdc ;
reg  hdd ;
reg  hea ;
reg  heb ;
reg  hec ;
reg  hed ;
reg  hfa ;
reg  hfb ;
reg  hfc ;
reg  hfd ;
reg  hga ;
reg  hgb ;
reg  hgc ;
reg  hgd ;
reg  hha ;
reg  hhb ;
reg  hhc ;
reg  hhd ;
reg  hia ;
reg  hib ;
reg  hic ;
reg  hid ;
reg  hja ;
reg  hjb ;
reg  hjc ;
reg  hjd ;
reg  hka ;
reg  hkb ;
reg  hkc ;
reg  hkd ;
reg  hla ;
reg  hlb ;
reg  hlc ;
reg  hld ;
reg  hma ;
reg  hmb ;
reg  hmc ;
reg  hmd ;
reg  hna ;
reg  hnb ;
reg  hnc ;
reg  hnd ;
reg  hoa ;
reg  hob ;
reg  hoc ;
reg  hod ;
reg  hpa ;
reg  hpb ;
reg  hpc ;
reg  hpd ;
reg  KAB ;
reg  KAC ;
reg  KAD ;
reg  KBC ;
reg  KBD ;
reg  KCD ;
reg  lbc ;
reg  lbd ;
reg  lcd ;
reg  maa ;
reg  mab ;
reg  mac ;
reg  mba ;
reg  mbb ;
reg  mbc ;
reg  mca ;
reg  mcb ;
reg  mcc ;
reg  mda ;
reg  mdb ;
reg  mdc ;
reg  nba ;
reg  nbb ;
reg  nbc ;
reg  nca ;
reg  ncb ;
reg  ncc ;
reg  nda ;
reg  ndb ;
reg  ndc ;
reg  OAA ;
reg  OAB ;
reg  OAC ;
reg  OAD ;
reg  OAE ;
reg  OAF ;
reg  OAG ;
reg  OAH ;
reg  OAI ;
reg  OAJ ;
reg  OAK ;
reg  OAL ;
reg  OAM ;
reg  OAN ;
reg  OAO ;
reg  OAP ;
reg  OBA ;
reg  OBB ;
reg  OBC ;
reg  OBD ;
reg  OBE ;
reg  OBF ;
reg  OBG ;
reg  OBH ;
reg  OBI ;
reg  OBJ ;
reg  OBK ;
reg  OBL ;
reg  OBM ;
reg  OBN ;
reg  OBO ;
reg  OBP ;
reg  OCA ;
reg  OCB ;
reg  OCC ;
reg  OCD ;
reg  OCE ;
reg  OCF ;
reg  OCG ;
reg  OCH ;
reg  OCI ;
reg  OCJ ;
reg  OCK ;
reg  OCL ;
reg  OCM ;
reg  OCN ;
reg  OCO ;
reg  OCP ;
reg  ODA ;
reg  ODB ;
reg  ODC ;
reg  ODD ;
reg  ODE ;
reg  ODF ;
reg  ODG ;
reg  ODH ;
reg  ODI ;
reg  ODJ ;
reg  ODK ;
reg  ODL ;
reg  ODM ;
reg  ODN ;
reg  ODO ;
reg  ODP ;
reg  oea ;
reg  OEB ;
reg  OEC ;
reg  OFA ;
reg  OFB ;
reg  ONA ;
reg  qaa ;
reg  QAB ;
reg  QAC ;
reg  qad ;
reg  qba ;
reg  QBB ;
reg  qbc ;
reg  QBD ;
reg  QBE ;
reg  QBF ;
reg  QBI ;
reg  QCA ;
reg  QCB ;
reg  QCE ;
reg  QCF ;
reg  QCG ;
reg  QDA ;
reg  QDB ;
reg  QDC ;
reg  QDD ;
reg  QDE ;
reg  qea ;
reg  QEB ;
reg  QEC ;
reg  QED ;
reg  QEE ;
reg  QEF ;
reg  QFA ;
reg  QFB ;
reg  QFC ;
reg  QFD ;
reg  qga ;
reg  qgb ;
reg  QHA ;
reg  QIA ;
reg  QIB ;
reg  QJA ;
reg  QJB ;
reg  QJC ;
reg  QJD ;
reg  QJE ;
reg  QNA ;
reg  QNB ;
reg  QNC ;
reg  SAA ;
reg  SAB ;
reg  SAC ;
reg  SAD ;
reg  SBA ;
reg  SBB ;
reg  SBC ;
reg  SBD ;
reg  SCA ;
reg  SCB ;
reg  SCC ;
reg  SCD ;
reg  SDA ;
reg  SDB ;
reg  SDC ;
reg  SDD ;
reg  SEA ;
reg  SEB ;
reg  SEC ;
reg  SED ;
reg  SFA ;
reg  SFB ;
reg  SFC ;
reg  SFD ;
reg  SGA ;
reg  SGB ;
reg  SGC ;
reg  SGD ;
reg  SHA ;
reg  SHB ;
reg  SHC ;
reg  SHD ;
reg  SIA ;
reg  SIB ;
reg  SIC ;
reg  SID ;
reg  SJA ;
reg  SJB ;
reg  SJC ;
reg  SJD ;
reg  SKA ;
reg  SKB ;
reg  SKC ;
reg  SKD ;
reg  SLA ;
reg  SLB ;
reg  SLC ;
reg  SLD ;
reg  SMA ;
reg  SMB ;
reg  SMC ;
reg  SMD ;
reg  SNA ;
reg  SNB ;
reg  SNC ;
reg  SND ;
reg  SOA ;
reg  SOB ;
reg  SOC ;
reg  SOD ;
reg  SPA ;
reg  SPB ;
reg  SPC ;
reg  SPD ;
reg  TAA ;
reg  TAB ;
reg  TAC ;
reg  TAD ;
reg  TAE ;
reg  TAF ;
reg  TAG ;
reg  TAH ;
reg  TDA ;
reg  TDB ;
reg  TDC ;
reg  TDD ;
reg  TDE ;
reg  TDF ;
reg  TDG ;
reg  TDH ;
reg  TDI ;
reg  TDJ ;
reg  TDK ;
reg  TDL ;
reg  TDM ;
reg  TDN ;
reg  TDO ;
reg  TDP ;
reg  TEA ;
reg  TEB ;
reg  TEC ;
reg  TED ;
reg  TFA ;
reg  TFB ;
reg  TFC ;
reg  TFD ;
reg  TGA ;
reg  TGB ;
reg  TGC ;
reg  TGD ;
reg  tha ;
reg  thb ;
reg  thc ;
reg  thd ;
reg  TIA ;
reg  TIB ;
reg  TIC ;
reg  TID ;
reg  tja ;
reg  tjb ;
reg  tjc ;
reg  tjd ;
reg  tka ;
reg  tkb ;
reg  UAA ;
reg  UAB ;
reg  UAC ;
reg  UAD ;
reg  UBA ;
reg  UBB ;
reg  UBC ;
reg  UBD ;
reg  UCA ;
reg  UCB ;
reg  UCC ;
reg  UCD ;
reg  UDA ;
reg  UDB ;
reg  UDC ;
reg  UDD ;
reg  UEA ;
reg  UEB ;
reg  UEC ;
reg  UED ;
reg  UFA ;
reg  UFB ;
reg  UFC ;
reg  UFD ;
reg  UGA ;
reg  UGB ;
reg  UGC ;
reg  UGD ;
reg  UHA ;
reg  UHB ;
reg  UHC ;
reg  UHD ;
reg  UIA ;
reg  UIB ;
reg  UIC ;
reg  UID ;
reg  UJA ;
reg  UJB ;
reg  UJC ;
reg  UJD ;
reg  UKA ;
reg  UKB ;
reg  UKC ;
reg  UKD ;
reg  ULA ;
reg  ULB ;
reg  ULC ;
reg  ULD ;
reg  UMA ;
reg  UMB ;
reg  UMC ;
reg  UMD ;
reg  UNA ;
reg  UNB ;
reg  UNC ;
reg  UND ;
reg  UOA ;
reg  UOB ;
reg  UOC ;
reg  UOD ;
reg  UPA ;
reg  UPB ;
reg  UPC ;
reg  UPD ;
reg  UPE ;
reg  XAA ;
reg  XAB ;
reg  XAC ;
reg  XAD ;
reg  XBA ;
reg  XBB ;
reg  XBC ;
reg  XBD ;
reg  XCA ;
reg  XCB ;
reg  XCC ;
reg  XCD ;
reg  XDA ;
reg  XDB ;
reg  XDC ;
reg  XDD ;
reg  XEA ;
reg  XEB ;
reg  XEC ;
reg  XED ;
reg  XFA ;
reg  XFB ;
reg  XFC ;
reg  XFD ;
reg  XGA ;
reg  XGB ;
reg  XGC ;
reg  XGD ;
reg  XHA ;
reg  XHB ;
reg  XHC ;
reg  XHD ;
reg  XIB ;
reg  XIC ;
reg  XID ;
reg  XJA ;
reg  XJB ;
reg  XJC ;
reg  XJD ;
reg  XKA ;
reg  XKB ;
reg  XKC ;
reg  XKD ;
reg  XLA ;
reg  XLB ;
reg  XLC ;
reg  XLD ;
reg  XMA ;
reg  XMB ;
reg  XMC ;
reg  XMD ;
reg  XNA ;
reg  XNB ;
reg  XNC ;
reg  XND ;
reg  XOA ;
reg  XOB ;
reg  XOC ;
reg  XOD ;
reg  XPA ;
reg  XPB ;
reg  XPC ;
reg  XPD ;
wire  AAA ;
wire  AAB ;
wire  AAC ;
wire  AAD ;
wire  ABA ;
wire  ABB ;
wire  ABC ;
wire  ABD ;
wire  ACA ;
wire  ACB ;
wire  ACC ;
wire  ACD ;
wire  ADA ;
wire  ADB ;
wire  ADC ;
wire  ADD ;
wire  AEA ;
wire  AEB ;
wire  AEC ;
wire  AED ;
wire  AFA ;
wire  AFB ;
wire  AFC ;
wire  AFD ;
wire  AGA ;
wire  AGB ;
wire  AGC ;
wire  AGD ;
wire  AHA ;
wire  AHB ;
wire  AHC ;
wire  AHD ;
wire  AIA ;
wire  AIB ;
wire  AIC ;
wire  AID ;
wire  AJA ;
wire  AJB ;
wire  AJC ;
wire  AJD ;
wire  AKA ;
wire  AKB ;
wire  AKC ;
wire  AKD ;
wire  ALA ;
wire  ALB ;
wire  ALC ;
wire  ALD ;
wire  AMA ;
wire  AMB ;
wire  AMC ;
wire  AMD ;
wire  ANA ;
wire  ANB ;
wire  ANC ;
wire  ANDD  ;
wire  AOA ;
wire  AOB ;
wire  AOC ;
wire  AOD ;
wire  APA ;
wire  APB ;
wire  APC ;
wire  APD ;
wire  baa ;
wire  bab ;
wire  bac ;
wire  bad ;
wire  bba ;
wire  bbb ;
wire  bbc ;
wire  bbd ;
wire  bbf ;
wire  bbg ;
wire  bca ;
wire  bcb ;
wire  bcc ;
wire  bcd ;
wire  bcf ;
wire  bcg ;
wire  bda ;
wire  bdb ;
wire  bdc ;
wire  bdd ;
wire  bdf ;
wire  bdg ;
wire  bea ;
wire  beb ;
wire  bec ;
wire  bed ;
wire  bef ;
wire  beg ;
wire  bfa ;
wire  bfb ;
wire  bfc ;
wire  bfd ;
wire  bff ;
wire  bfg ;
wire  bga ;
wire  bgb ;
wire  bgc ;
wire  bgd ;
wire  bgf ;
wire  bgg ;
wire  bha ;
wire  bhb ;
wire  bhc ;
wire  bhd ;
wire  bhf ;
wire  bhg ;
wire  bia ;
wire  bib ;
wire  bic ;
wire  bid ;
wire  bif ;
wire  big ;
wire  bja ;
wire  bjb ;
wire  bjc ;
wire  bjd ;
wire  bjf ;
wire  bjg ;
wire  bka ;
wire  bkb ;
wire  bkc ;
wire  bkd ;
wire  bkf ;
wire  bkg ;
wire  bla ;
wire  blb ;
wire  blc ;
wire  bld ;
wire  blf ;
wire  blg ;
wire  BLG ;
wire  bma ;
wire  bmb ;
wire  bmc ;
wire  bmd ;
wire  bmf ;
wire  bmg ;
wire  bna ;
wire  bnb ;
wire  bnc ;
wire  bnd ;
wire  bnf ;
wire  bng ;
wire  boa ;
wire  bob ;
wire  boc ;
wire  bod ;
wire  bof ;
wire  bog ;
wire  bpa ;
wire  bpb ;
wire  bpc ;
wire  bpd ;
wire  caa ;
wire  CAA ;
wire  cab ;
wire  CAB ;
wire  cac ;
wire  CAC ;
wire  cad ;
wire  CAD ;
wire  cae ;
wire  CAE ;
wire  cbb ;
wire  CBB ;
wire  cbc ;
wire  CBC ;
wire  cbd ;
wire  CBD ;
wire  cbe ;
wire  CBE ;
wire  ccb ;
wire  CCB ;
wire  ccc ;
wire  CCC ;
wire  ccd ;
wire  CCD ;
wire  cce ;
wire  CCE ;
wire  cdb ;
wire  CDB ;
wire  cdc ;
wire  CDC ;
wire  cdd ;
wire  CDD ;
wire  cde ;
wire  CDE ;
wire  ceb ;
wire  CEB ;
wire  cec ;
wire  CEC ;
wire  ced ;
wire  CED ;
wire  cee ;
wire  CEE ;
wire  cfb ;
wire  CFB ;
wire  cfc ;
wire  CFC ;
wire  cfd ;
wire  CFD ;
wire  cfe ;
wire  CFE ;
wire  cgb ;
wire  CGB ;
wire  cgc ;
wire  CGC ;
wire  cgd ;
wire  CGD ;
wire  cge ;
wire  CGE ;
wire  chb ;
wire  CHB ;
wire  chc ;
wire  CHC ;
wire  chd ;
wire  CHD ;
wire  che ;
wire  CHE ;
wire  cib ;
wire  CIB ;
wire  cic ;
wire  CIC ;
wire  cid ;
wire  CID ;
wire  cie ;
wire  CIE ;
wire  cjb ;
wire  CJB ;
wire  cjc ;
wire  CJC ;
wire  cjd ;
wire  CJD ;
wire  cje ;
wire  CJE ;
wire  ckb ;
wire  CKB ;
wire  ckc ;
wire  CKC ;
wire  ckd ;
wire  CKD ;
wire  cke ;
wire  CKE ;
wire  clb ;
wire  CLB ;
wire  clc ;
wire  CLC ;
wire  cld ;
wire  CLD ;
wire  cle ;
wire  CLE ;
wire  cmb ;
wire  CMB ;
wire  cmc ;
wire  CMC ;
wire  cmd ;
wire  CMD ;
wire  cme ;
wire  CME ;
wire  cnb ;
wire  CNB ;
wire  cnc ;
wire  CNC ;
wire  cnd ;
wire  CND ;
wire  cne ;
wire  CNE ;
wire  cob ;
wire  COB ;
wire  coc ;
wire  COC ;
wire  cod ;
wire  COD ;
wire  coe ;
wire  COE ;
wire  cpb ;
wire  CPB ;
wire  cpc ;
wire  CPC ;
wire  cpd ;
wire  CPD ;
wire  dbb ;
wire  DBB ;
wire  dbc ;
wire  DBC ;
wire  dbd ;
wire  DBD ;
wire  dcb ;
wire  DCB ;
wire  dcc ;
wire  DCC ;
wire  dcd ;
wire  DCD ;
wire  ddb ;
wire  DDB ;
wire  ddc ;
wire  DDC ;
wire  ddd ;
wire  DDD ;
wire  deb ;
wire  DEB ;
wire  dec ;
wire  DEC ;
wire  ded ;
wire  DED ;
wire  DFB ;
wire  dfc ;
wire  DFC ;
wire  dfd ;
wire  DFD ;
wire  dgb ;
wire  DGB ;
wire  dgc ;
wire  DGC ;
wire  dgd ;
wire  DGD ;
wire  dhb ;
wire  DHB ;
wire  dhc ;
wire  DHC ;
wire  dhd ;
wire  DHD ;
wire  dib ;
wire  DIB ;
wire  dic ;
wire  DIC ;
wire  did ;
wire  DID ;
wire  djb ;
wire  DJB ;
wire  djc ;
wire  DJC ;
wire  djd ;
wire  DJD ;
wire  dkb ;
wire  DKB ;
wire  dkc ;
wire  DKC ;
wire  dkd ;
wire  DKD ;
wire  dlb ;
wire  DLB ;
wire  dlc ;
wire  DLC ;
wire  dld ;
wire  DLD ;
wire  dmb ;
wire  DMB ;
wire  dmc ;
wire  DMC ;
wire  dmd ;
wire  DMD ;
wire  dnb ;
wire  DNB ;
wire  dnc ;
wire  DNC ;
wire  dnd ;
wire  DND ;
wire  dob ;
wire  DOB ;
wire  doc ;
wire  DOC ;
wire  dod ;
wire  DOD ;
wire  dpb ;
wire  DPB ;
wire  dpc ;
wire  DPC ;
wire  dpd ;
wire  DPD ;
wire  eaa ;
wire  EAA ;
wire  eab ;
wire  EAB ;
wire  eac ;
wire  EAC ;
wire  ead ;
wire  EAD ;
wire  eba ;
wire  EBA ;
wire  ebb ;
wire  EBB ;
wire  ebc ;
wire  EBC ;
wire  ebd ;
wire  EBD ;
wire  eca ;
wire  ECA ;
wire  ecb ;
wire  ECB ;
wire  ecc ;
wire  ECC ;
wire  ecd ;
wire  ECD ;
wire  eda ;
wire  EDA ;
wire  edb ;
wire  EDB ;
wire  edc ;
wire  EDC ;
wire  edd ;
wire  EDD ;
wire  eea ;
wire  EEA ;
wire  eeb ;
wire  EEB ;
wire  eec ;
wire  EEC ;
wire  eed ;
wire  EED ;
wire  efa ;
wire  EFA ;
wire  efb ;
wire  EFB ;
wire  efc ;
wire  EFC ;
wire  efd ;
wire  EFD ;
wire  ega ;
wire  EGA ;
wire  egb ;
wire  EGB ;
wire  egc ;
wire  EGC ;
wire  egd ;
wire  EGD ;
wire  eha ;
wire  EHA ;
wire  ehb ;
wire  EHB ;
wire  ehc ;
wire  EHC ;
wire  ehd ;
wire  EHD ;
wire  eia ;
wire  EIA ;
wire  eib ;
wire  EIB ;
wire  eic ;
wire  EIC ;
wire  eid ;
wire  EID ;
wire  eja ;
wire  EJA ;
wire  ejb ;
wire  EJB ;
wire  ejc ;
wire  EJC ;
wire  ejd ;
wire  EJD ;
wire  eka ;
wire  EKA ;
wire  ekb ;
wire  EKB ;
wire  ekc ;
wire  EKC ;
wire  ekd ;
wire  EKD ;
wire  ela ;
wire  ELA ;
wire  elb ;
wire  ELB ;
wire  elc ;
wire  ELC ;
wire  eld ;
wire  ELD ;
wire  ema ;
wire  EMA ;
wire  emb ;
wire  EMB ;
wire  emc ;
wire  EMC ;
wire  emd ;
wire  EMD ;
wire  ena ;
wire  ENA ;
wire  enb ;
wire  ENB ;
wire  enc ;
wire  ENC ;
wire  endd ;
wire  ENDD  ;
wire  eoa ;
wire  EOA ;
wire  eob ;
wire  EOB ;
wire  eoc ;
wire  EOC ;
wire  eod ;
wire  EOD ;
wire  epa ;
wire  EPA ;
wire  epb ;
wire  EPB ;
wire  epc ;
wire  EPC ;
wire  epd ;
wire  EPD ;
wire  fab ;
wire  FAB ;
wire  fac ;
wire  FAC ;
wire  fad ;
wire  FAD ;
wire  fae ;
wire  FAE ;
wire  faf ;
wire  FAF ;
wire  fag ;
wire  FAG ;
wire  fah ;
wire  FAH ;
wire  fai ;
wire  FAI ;
wire  faj ;
wire  FAJ ;
wire  fak ;
wire  FAK ;
wire  fal ;
wire  FAL ;
wire  fam ;
wire  FAM ;
wire  fan ;
wire  FAN ;
wire  fao ;
wire  FAO ;
wire  fbf ;
wire  FBF ;
wire  fbg ;
wire  FBG ;
wire  fbj ;
wire  FBJ ;
wire  fbk ;
wire  FBK ;
wire  fbn ;
wire  FBN ;
wire  fbo ;
wire  FBO ;
wire  GAA ;
wire  GAB ;
wire  GAC ;
wire  GAD ;
wire  GBA ;
wire  GBB ;
wire  GBC ;
wire  GBD ;
wire  GCA ;
wire  GCB ;
wire  GCC ;
wire  GCD ;
wire  GDA ;
wire  GDB ;
wire  GDC ;
wire  GDD ;
wire  GEA ;
wire  GEB ;
wire  GEC ;
wire  GED ;
wire  GFA ;
wire  GFB ;
wire  GFC ;
wire  GFD ;
wire  GGA ;
wire  GGB ;
wire  GGC ;
wire  GGD ;
wire  GHA ;
wire  GHB ;
wire  GHC ;
wire  GHD ;
wire  GIA ;
wire  GIB ;
wire  GIC ;
wire  GID ;
wire  GJA ;
wire  GJB ;
wire  GJC ;
wire  GJD ;
wire  GKA ;
wire  GKB ;
wire  GKC ;
wire  GKD ;
wire  GLA ;
wire  GLB ;
wire  GLC ;
wire  GLD ;
wire  GMA ;
wire  GMB ;
wire  GMC ;
wire  GMD ;
wire  GNA ;
wire  GNB ;
wire  GNC ;
wire  GND ;
wire  GOA ;
wire  GOB ;
wire  GOC ;
wire  GOD ;
wire  GPA ;
wire  GPB ;
wire  GPC ;
wire  GPD ;
wire  HBA ;
wire  HBB ;
wire  HBC ;
wire  HBD ;
wire  HCA ;
wire  HCB ;
wire  HCC ;
wire  HCD ;
wire  HDA ;
wire  HDB ;
wire  HDC ;
wire  HDD ;
wire  HEA ;
wire  HEB ;
wire  HEC ;
wire  HED ;
wire  HFA ;
wire  HFB ;
wire  HFC ;
wire  HFD ;
wire  HGA ;
wire  HGB ;
wire  HGC ;
wire  HGD ;
wire  HHA ;
wire  HHB ;
wire  HHC ;
wire  HHD ;
wire  HIA ;
wire  HIB ;
wire  HIC ;
wire  HID ;
wire  HJA ;
wire  HJB ;
wire  HJC ;
wire  HJD ;
wire  HKA ;
wire  HKB ;
wire  HKC ;
wire  HKD ;
wire  HLA ;
wire  HLB ;
wire  HLC ;
wire  HLD ;
wire  HMA ;
wire  HMB ;
wire  HMC ;
wire  HMD ;
wire  HNA ;
wire  HNB ;
wire  HNC ;
wire  HND ;
wire  HOA ;
wire  HOB ;
wire  HOC ;
wire  HOD ;
wire  HPA ;
wire  HPB ;
wire  HPC ;
wire  HPD ;
wire  iaa ;
wire  iab ;
wire  iac ;
wire  iad ;
wire  iae ;
wire  iaf ;
wire  iag ;
wire  iah ;
wire  iai ;
wire  iaj ;
wire  iak ;
wire  ial ;
wire  iam ;
wire  ian ;
wire  iao ;
wire  iap ;
wire  iba ;
wire  ibb ;
wire  ibc ;
wire  ibd ;
wire  ibe ;
wire  ibf ;
wire  ibg ;
wire  ibh ;
wire  ibi ;
wire  ibj ;
wire  ibk ;
wire  ibl ;
wire  ibm ;
wire  ibn ;
wire  ibo ;
wire  ibp ;
wire  ica ;
wire  icb ;
wire  icc ;
wire  icd ;
wire  ice ;
wire  icf ;
wire  icg ;
wire  ich ;
wire  ici ;
wire  icj ;
wire  ick ;
wire  icl ;
wire  icm ;
wire  icn ;
wire  ico ;
wire  icp ;
wire  ida ;
wire  idb ;
wire  idc ;
wire  idd ;
wire  ide ;
wire  idf ;
wire  idg ;
wire  idh ;
wire  idi ;
wire  idj ;
wire  idk ;
wire  idl ;
wire  idm ;
wire  idn ;
wire  ido ;
wire  idp ;
wire  iea ;
wire  ieb ;
wire  iec ;
wire  ied ;
wire  iee ;
wire  ief ;
wire  ieg ;
wire  ieh ;
wire  iei ;
wire  iej ;
wire  iek ;
wire  iel ;
wire  iem ;
wire  ien ;
wire  ieo ;
wire  iep ;
wire  ifa ;
wire  ifb ;
wire  ifc ;
wire  ifd ;
wire  ife ;
wire  ifff  ;
wire  ifg ;
wire  ifh ;
wire  ifi ;
wire  ifj ;
wire  ifk ;
wire  ifl ;
wire  ifm ;
wire  ifn ;
wire  ifo ;
wire  ifp ;
wire  iga ;
wire  igb ;
wire  igc ;
wire  igd ;
wire  ige ;
wire  igf ;
wire  igg ;
wire  igh ;
wire  igi ;
wire  igj ;
wire  igk ;
wire  igl ;
wire  igm ;
wire  ign ;
wire  igo ;
wire  igp ;
wire  iha ;
wire  ihb ;
wire  ihc ;
wire  ihd ;
wire  ihe ;
wire  ihf ;
wire  ihg ;
wire  ihh ;
wire  ihi ;
wire  ihj ;
wire  ihk ;
wire  ihl ;
wire  ihm ;
wire  ihn ;
wire  iho ;
wire  ihp ;
wire  ima ;
wire  ira ;
wire  irb ;
wire  irc ;
wire  ird ;
wire  jaa ;
wire  JAA ;
wire  jab ;
wire  JAB ;
wire  jac ;
wire  JAC ;
wire  jad ;
wire  JAD ;
wire  jae ;
wire  JAE ;
wire  jaf ;
wire  JAF ;
wire  jag ;
wire  JAG ;
wire  jah ;
wire  JAH ;
wire  jai ;
wire  JAI ;
wire  jaj ;
wire  JAJ ;
wire  jak ;
wire  JAK ;
wire  jal ;
wire  JAL ;
wire  jam ;
wire  JAM ;
wire  jan ;
wire  JAN ;
wire  jao ;
wire  JAO ;
wire  jap ;
wire  JAP ;
wire  jba ;
wire  JBA ;
wire  jbb ;
wire  JBB ;
wire  jca ;
wire  JCA ;
wire  jda ;
wire  JDA ;
wire  jqa ;
wire  JQA ;
wire  kab ;
wire  kac ;
wire  kad ;
wire  kbc ;
wire  kbd ;
wire  kcd ;
wire  LBC ;
wire  LBD ;
wire  LCD ;
wire  MAA ;
wire  MAB ;
wire  MAC ;
wire  MBA ;
wire  MBB ;
wire  MBC ;
wire  MCA ;
wire  MCB ;
wire  MCC ;
wire  MDA ;
wire  MDB ;
wire  MDC ;
wire  NBA ;
wire  NBB ;
wire  NBC ;
wire  NCA ;
wire  NCB ;
wire  NCC ;
wire  NDA ;
wire  NDB ;
wire  NDC ;
wire  oaa ;
wire  oab ;
wire  oac ;
wire  oad ;
wire  oae ;
wire  oaf ;
wire  oag ;
wire  oah ;
wire  oai ;
wire  oaj ;
wire  oak ;
wire  oal ;
wire  oam ;
wire  oan ;
wire  oao ;
wire  oap ;
wire  oba ;
wire  obb ;
wire  obc ;
wire  obd ;
wire  obe ;
wire  obf ;
wire  obg ;
wire  obh ;
wire  obi ;
wire  obj ;
wire  obk ;
wire  obl ;
wire  obm ;
wire  obn ;
wire  obo ;
wire  obp ;
wire  oca ;
wire  ocb ;
wire  occ ;
wire  ocd ;
wire  oce ;
wire  ocf ;
wire  ocg ;
wire  och ;
wire  oci ;
wire  ocj ;
wire  ock ;
wire  ocl ;
wire  ocm ;
wire  ocn ;
wire  oco ;
wire  ocp ;
wire  oda ;
wire  odb ;
wire  odc ;
wire  odd ;
wire  ode ;
wire  odf ;
wire  odg ;
wire  odh ;
wire  odi ;
wire  odj ;
wire  odk ;
wire  odl ;
wire  odm ;
wire  odn ;
wire  odo ;
wire  odp ;
wire  OEA ;
wire  oeb ;
wire  oec ;
wire  ofa ;
wire  ofb ;
wire  ona ;
wire  pab ;
wire  PAB ;
wire  pac ;
wire  PAC ;
wire  pad ;
wire  PAD ;
wire  pba ;
wire  PBA ;
wire  pbb ;
wire  PBB ;
wire  pbc ;
wire  PBC ;
wire  pbd ;
wire  PBD ;
wire  pca ;
wire  PCA ;
wire  pcb ;
wire  PCB ;
wire  pcc ;
wire  PCC ;
wire  pcd ;
wire  PCD ;
wire  pda ;
wire  PDA ;
wire  pdb ;
wire  PDB ;
wire  pdc ;
wire  PDC ;
wire  pdd ;
wire  PDD ;
wire  QAA ;
wire  qab ;
wire  qac ;
wire  QAD ;
wire  QBA ;
wire  qbb ;
wire  QBC ;
wire  qbd ;
wire  qbe ;
wire  qbf ;
wire  qbi ;
wire  qca ;
wire  qcb ;
wire  qce ;
wire  qcf ;
wire  qcg ;
wire  qda ;
wire  qdb ;
wire  qdc ;
wire  qdd ;
wire  qde ;
wire  QEA ;
wire  qeb ;
wire  qec ;
wire  qed ;
wire  qee ;
wire  qef ;
wire  qfa ;
wire  qfb ;
wire  qfc ;
wire  qfd ;
wire  QGA ;
wire  QGB ;
wire  qha ;
wire  qia ;
wire  qib ;
wire  qja ;
wire  qjb ;
wire  qjc ;
wire  qjd ;
wire  qje ;
wire  qna ;
wire  qnb ;
wire  qnc ;
wire  saa ;
wire  sab ;
wire  sac ;
wire  sad ;
wire  sba ;
wire  sbb ;
wire  sbc ;
wire  sbd ;
wire  sca ;
wire  scb ;
wire  scc ;
wire  scd ;
wire  sda ;
wire  sdb ;
wire  sdc ;
wire  sdd ;
wire  sea ;
wire  seb ;
wire  sec ;
wire  sed ;
wire  sfa ;
wire  sfb ;
wire  sfc ;
wire  sfd ;
wire  sga ;
wire  sgb ;
wire  sgc ;
wire  sgd ;
wire  sha ;
wire  shb ;
wire  shc ;
wire  shd ;
wire  sia ;
wire  sib ;
wire  sic ;
wire  sid ;
wire  sja ;
wire  sjb ;
wire  sjc ;
wire  sjd ;
wire  ska ;
wire  skb ;
wire  skc ;
wire  skd ;
wire  sla ;
wire  slb ;
wire  slc ;
wire  sld ;
wire  sma ;
wire  smb ;
wire  smc ;
wire  smd ;
wire  sna ;
wire  snb ;
wire  snc ;
wire  snd ;
wire  soa ;
wire  sob ;
wire  soc ;
wire  sod ;
wire  spa ;
wire  spb ;
wire  spc ;
wire  spd ;
wire  taa ;
wire  tab ;
wire  tac ;
wire  tad ;
wire  tae ;
wire  taf ;
wire  tag ;
wire  tah ;
wire  tda ;
wire  tdb ;
wire  tdc ;
wire  tdd ;
wire  tde ;
wire  tdf ;
wire  tdg ;
wire  tdh ;
wire  tdi ;
wire  tdj ;
wire  tdk ;
wire  tdl ;
wire  tdm ;
wire  tdn ;
wire  tdo ;
wire  tdp ;
wire  tea ;
wire  teb ;
wire  tec ;
wire  ted ;
wire  tfa ;
wire  tfb ;
wire  tfc ;
wire  tfd ;
wire  tga ;
wire  tgb ;
wire  tgc ;
wire  tgd ;
wire  THA ;
wire  THB ;
wire  THC ;
wire  THD ;
wire  tia ;
wire  tib ;
wire  tic ;
wire  tid ;
wire  TJA ;
wire  TJB ;
wire  TJC ;
wire  TJD ;
wire  TKA ;
wire  TKB ;
wire  uaa ;
wire  uab ;
wire  uac ;
wire  uad ;
wire  uba ;
wire  ubb ;
wire  ubc ;
wire  ubd ;
wire  uca ;
wire  ucb ;
wire  ucc ;
wire  ucd ;
wire  uda ;
wire  udb ;
wire  udc ;
wire  udd ;
wire  uea ;
wire  ueb ;
wire  uec ;
wire  ued ;
wire  ufa ;
wire  ufb ;
wire  ufc ;
wire  ufd ;
wire  uga ;
wire  ugb ;
wire  ugc ;
wire  ugd ;
wire  uha ;
wire  uhb ;
wire  uhc ;
wire  uhd ;
wire  uia ;
wire  uib ;
wire  uic ;
wire  uid ;
wire  uja ;
wire  ujb ;
wire  ujc ;
wire  ujd ;
wire  uka ;
wire  ukb ;
wire  ukc ;
wire  ukd ;
wire  ula ;
wire  ulb ;
wire  ulc ;
wire  uld ;
wire  uma ;
wire  umb ;
wire  umc ;
wire  umd ;
wire  una ;
wire  unb ;
wire  unc ;
wire  und ;
wire  uoa ;
wire  uob ;
wire  uoc ;
wire  uod ;
wire  upa ;
wire  upb ;
wire  upc ;
wire  upd ;
wire  upe ;
wire  waa ;
wire  WAA ;
wire  wab ;
wire  WAB ;
wire  wac ;
wire  WAC ;
wire  wad ;
wire  WAD ;
wire  wba ;
wire  WBA ;
wire  wbb ;
wire  WBB ;
wire  wbc ;
wire  WBC ;
wire  wbd ;
wire  WBD ;
wire  wca ;
wire  WCA ;
wire  wcb ;
wire  WCB ;
wire  wcc ;
wire  WCC ;
wire  wcd ;
wire  WCD ;
wire  wda ;
wire  WDA ;
wire  wdb ;
wire  WDB ;
wire  wdc ;
wire  WDC ;
wire  wdd ;
wire  WDD ;
wire  wea ;
wire  WEA ;
wire  web ;
wire  WEB ;
wire  wec ;
wire  WEC ;
wire  wed ;
wire  WED ;
wire  wfa ;
wire  WFA ;
wire  wfb ;
wire  WFB ;
wire  wfc ;
wire  WFC ;
wire  wfd ;
wire  WFD ;
wire  wga ;
wire  WGA ;
wire  wgb ;
wire  WGB ;
wire  wgc ;
wire  WGC ;
wire  wgd ;
wire  WGD ;
wire  wha ;
wire  WHA ;
wire  whb ;
wire  WHB ;
wire  whc ;
wire  WHC ;
wire  whd ;
wire  WHD ;
wire  wib ;
wire  WIB ;
wire  wic ;
wire  WIC ;
wire  wid ;
wire  WID ;
wire  wja ;
wire  WJA ;
wire  wjb ;
wire  WJB ;
wire  wjc ;
wire  WJC ;
wire  wjd ;
wire  WJD ;
wire  wka ;
wire  WKA ;
wire  wkb ;
wire  WKB ;
wire  wkc ;
wire  WKC ;
wire  wkd ;
wire  WKD ;
wire  wla ;
wire  WLA ;
wire  wlb ;
wire  WLB ;
wire  wlc ;
wire  WLC ;
wire  wld ;
wire  WLD ;
wire  wma ;
wire  WMA ;
wire  wmb ;
wire  WMB ;
wire  wmc ;
wire  WMC ;
wire  wmd ;
wire  WMD ;
wire  wna ;
wire  WNA ;
wire  wnb ;
wire  WNB ;
wire  wnc ;
wire  WNC ;
wire  wnd ;
wire  WND ;
wire  woa ;
wire  WOA ;
wire  wob ;
wire  WOB ;
wire  woc ;
wire  WOC ;
wire  wod ;
wire  WOD ;
wire  wpa ;
wire  WPA ;
wire  wpb ;
wire  WPB ;
wire  wpc ;
wire  WPC ;
wire  wpd ;
wire  WPD ;
wire  xaa ;
wire  xab ;
wire  xac ;
wire  xad ;
wire  xba ;
wire  xbb ;
wire  xbc ;
wire  xbd ;
wire  xca ;
wire  xcb ;
wire  xcc ;
wire  xcd ;
wire  xda ;
wire  xdb ;
wire  xdc ;
wire  xdd ;
wire  xea ;
wire  xeb ;
wire  xec ;
wire  xed ;
wire  xfa ;
wire  xfb ;
wire  xfc ;
wire  xfd ;
wire  xga ;
wire  xgb ;
wire  xgc ;
wire  xgd ;
wire  xha ;
wire  xhb ;
wire  xhc ;
wire  xhd ;
wire  xib ;
wire  xic ;
wire  xid ;
wire  xja ;
wire  xjb ;
wire  xjc ;
wire  xjd ;
wire  xka ;
wire  xkb ;
wire  xkc ;
wire  xkd ;
wire  xla ;
wire  xlb ;
wire  xlc ;
wire  xld ;
wire  xma ;
wire  xmb ;
wire  xmc ;
wire  xmd ;
wire  xna ;
wire  xnb ;
wire  xnc ;
wire  xnd ;
wire  xoa ;
wire  xob ;
wire  xoc ;
wire  xod ;
wire  xpa ;
wire  xpb ;
wire  xpc ;
wire  xpd ;
wire  ZZI ;
wire  ZZO ;
assign ZZI = 1'b1;
assign ZZO = 1'b0;
assign GAA = ~gaa;  //complement 
assign GAB = ~gab;  //complement 
assign HIC = ~hic;  //complement 
assign GAC = ~gac;  //complement 
assign GAD = ~gad;  //complement 
assign GIA = ~gia;  //complement 
assign HIA = ~hia;  //complement 
assign HIB = ~hib;  //complement 
assign GIB = ~gib;  //complement 
assign dib =  bia  ; 
assign DIB = ~dib;  //complement 
assign dic =  aib & bia  |  bib  ; 
assign DIC = ~dic;  //complement 
assign GIC = ~gic;  //complement 
assign did =  bia & aib & aic  |  bib & aic  |  bic  ; 
assign DID = ~did; //complement 
assign GID = ~gid;  //complement 
assign HID = ~hid;  //complement 
assign tda = ~TDA;  //complement 
assign taa = ~TAA;  //complement 
assign TKA = ~tka;  //complement 
assign TKB = ~tkb;  //complement 
assign caa =  qfd  ; 
assign CAA = ~caa;  //complement 
assign cab =  aaa & qfd  |  baa  ; 
assign CAB = ~cab;  //complement 
assign EAA = ZZO & ~AAA & ~BAA  |  ZZO & ~AAA & BAA  |  ZZI & AAA & ~BAA  |  ZZO & AAA & BAA; 
assign eaa = ~EAA;  //complement 
assign EAB = ZZO & ~AAB & ~BAB  |         ZZO & ~AAB & BAB  |  ZZI & AAB & ~BAB  |  ZZO & AAB & BAB ; 
assign eab = ~EAB;  //complement 
assign CAC =  QFD & BAA & BAB  |  AAA & BAB  |  AAB  ; 
assign cac = ~CAC; //complement 
assign qfc = ~QFC;  //complement 
assign qfd = ~QFD;  //complement 
assign qia = ~QIA;  //complement 
assign qib = ~QIB;  //complement 
assign EAC = ZZO & ~AAC & ~BAC  |  ZZO & ~AAC & BAC  |  ZZI & AAC & ~BAC  |  ZZO & AAC & BAC; 
assign eac = ~EAC;  //complement 
assign EAD = ZZO & ~AAD & ~BAD  |         ZZO & ~AAD & BAD  |  ZZI & AAD & ~BAD  |  ZZO & AAD & BAD ; 
assign ead = ~EAD;  //complement 
assign CID =  AIA & BIB & BIC  |  AIB & BIC  |  AIC  ; 
assign cid = ~CID; //complement 
assign CAD =  QFD & BAA & BAB & BAC  |  AAA & BAB & BAC  |  AAB & BAC  |  AAC  ; 
assign cad = ~CAD;  //complement 
assign CIC =  BIB & AIA  |  AIB  ; 
assign cic = ~CIC;  //complement 
assign CAE =  QFD & BAA & BAB & BAC & BAD  |  AAA & BAB & BAC & BAD  |  AAB & BAC & BAD  |  AAC & BAD  |  AAD  ; 
assign cae = ~CAE;  //complement 
assign FAI =  BIA & BEF & BIG & BID  ; 
assign fai = ~FAI;  //complement  
assign kab = ~KAB;  //complement 
assign PCA =  KAC & LBC  |  KBC  ; 
assign pca = ~PCA; //complement 
assign EIA = ZZO & ~AIA & ~BIA  |  ZZO & ~AIA & BIA  |  ZZI & AIA & ~BIA  |  ZZO & AIA & BIA; 
assign eia = ~EIA;  //complement 
assign EIB = ZZO & ~AIB & ~BIB  |         ZZO & ~AIB & BIB  |  ZZI & AIB & ~BIB  |  ZZO & AIB & BIB ; 
assign eib = ~EIB;  //complement 
assign CIB =  AIA  ; 
assign cib = ~CIB;  //complement 
assign bib = ~BIB;  //complement 
assign bif = ~BIF;  //complement 
assign EIC = ZZO & ~AIC & ~BIC  |  ZZO & ~AIC & BIC  |  ZZI & AIC & ~BIC  |  ZZO & AIC & BIC; 
assign eic = ~EIC;  //complement 
assign EID = ZZO & ~AID & ~BID  |         ZZO & ~AID & BID  |  ZZI & AID & ~BID  |  ZZO & AID & BID ; 
assign eid = ~EID;  //complement 
assign bic = ~BIC;  //complement 
assign big = ~BIG;  //complement 
assign qde = ~QDE;  //complement 
assign tdi = ~TDI;  //complement 
assign CIE =  AEA & BIB & BIC & BID  |  AIB & BIC & BID  |  AIC & BID  |  AID  ; 
assign cie = ~CIE;  //complement 
assign AAA = ~aaa;  //complement 
assign baa = ~BAA;  //complement 
assign xaa = ~XAA;  //complement 
assign xab = ~XAB;  //complement 
assign xib = ~XIB;  //complement 
assign WAA =  SAA & xaa  |  saa & XAA  |  saa & xaa  |  SAA & XAA  ; 
assign waa = ~WAA; //complement 
assign wib =  SAA & xaa  |  saa & XAA  |  saa & xaa  |  saa & xaa  ; 
assign WIB = ~wib;  //complement 
assign saa = ~SAA;  //complement 
assign sab = ~SAB;  //complement 
assign AAB = ~aab;  //complement 
assign AAC = ~aac;  //complement 
assign oaa = ~OAA;  //complement 
assign oab = ~OAB;  //complement 
assign WAB =  SAB & xab & xib  |  sab & XAB & xib  |  sab & xab & XIB  |  SAB & XAB & XIB  ; 
assign wab = ~WAB; //complement 
assign wic =  SAB & xab & xib  |  sab & XAB & xib  |  sab & xab & XIB  |  sab & xab & xib  ; 
assign WIC = ~wic;  //complement 
assign uaa = ~UAA;  //complement 
assign uab = ~UAB;  //complement 
assign bac = ~BAC;  //complement 
assign xac = ~XAC;  //complement 
assign xad = ~XAD;  //complement 
assign xic = ~XIC;  //complement 
assign xid = ~XID;  //complement 
assign WAC =  SAC & xac & xic  |  sac & XAC & xic  |  sac & xac & XIC  |  SAC & XAC & XIC  ; 
assign wac = ~WAC; //complement 
assign wid =  SAC & xac & xic  |  sac & XAC & xic  |  sac & xac & XIC  |  sac & xac & xic  ; 
assign WID = ~wid;  //complement 
assign sac = ~SAC;  //complement 
assign sad = ~SAD;  //complement 
assign AAD = ~aad;  //complement 
assign bad = ~BAD;  //complement 
assign oac = ~OAC;  //complement 
assign oad = ~OAD;  //complement 
assign WAD =  SAD & xad & xid  |  sad & XAD & xid  |  sad & xad & XID  |  SAD & XAD & XID  ; 
assign wad = ~WAD; //complement 
assign wja =  SAD & xad & xid  |  sad & XAD & xid  |  sad & xad & XID  |  sad & xad & xid  ; 
assign WJA = ~wja;  //complement 
assign uac = ~UAC;  //complement 
assign uad = ~UAD;  //complement 
assign AIA = ~aia;  //complement 
assign bia = ~BIA;  //complement 
assign jaa =  uaa & uab & uac & uad  ; 
assign JAA = ~jaa;  //complement  
assign tea = ~TEA;  //complement 
assign teb = ~TEB;  //complement 
assign tec = ~TEC;  //complement 
assign ted = ~TED;  //complement 
assign sia = ~SIA;  //complement 
assign sib = ~SIB;  //complement 
assign AIB = ~aib;  //complement 
assign oca = ~OCA;  //complement 
assign ocb = ~OCB;  //complement 
assign qja = ~QJA;  //complement 
assign uib = ~UIB;  //complement 
assign uia = ~UIA;  //complement 
assign AIC = ~aic;  //complement 
assign jai =  uia & uib & uic & uid  ; 
assign JAI = ~jai;  //complement  
assign JCA =  QDA & qeb & qec  ; 
assign jca = ~JCA;  //complement 
assign bab = ~BAB;  //complement 
assign sic = ~SIC;  //complement 
assign sid = ~SID;  //complement 
assign AID = ~aid;  //complement 
assign bid = ~BID;  //complement 
assign occ = ~OCC;  //complement 
assign ocd = ~OCD;  //complement 
assign qda = ~QDA;  //complement 
assign qdb = ~QDB;  //complement 
assign qdc = ~QDC;  //complement 
assign qdd = ~QDD;  //complement 
assign uic = ~UIC;  //complement 
assign uid = ~UID;  //complement 
assign GBA = ~gba;  //complement 
assign HBA = ~hba;  //complement 
assign GBB = ~gbb;  //complement 
assign HBB = ~hbb;  //complement 
assign dbb =  bba  ; 
assign DBB = ~dbb;  //complement 
assign dbc =  abb & bba  |  bbb  ; 
assign DBC = ~dbc;  //complement 
assign HJC = ~hjc;  //complement 
assign GBC = ~gbc;  //complement 
assign HBC = ~hbc;  //complement 
assign dbd =  bba & abb & abc  |  bbb & abc  |  bbc  ; 
assign DBD = ~dbd; //complement 
assign GBD = ~gbd;  //complement 
assign HBD = ~hbd;  //complement 
assign GJA = ~gja;  //complement 
assign HJA = ~hja;  //complement 
assign HJB = ~hjb;  //complement 
assign GJB = ~gjb;  //complement 
assign djb =  bja  ; 
assign DJB = ~djb;  //complement 
assign djc =  ajb & bja  |  bjb  ; 
assign DJC = ~djc;  //complement 
assign GJC = ~gjc;  //complement 
assign djd =  bja & ajb & ajc  |  bjb & ajc  |  bjc  ; 
assign DJD = ~djd; //complement 
assign GJD = ~gjd;  //complement 
assign HJD = ~hjd;  //complement 
assign bca = ~BCA;  //complement 
assign tab = ~TAB;  //complement 
assign sca = ~SCA;  //complement 
assign EBA = ZZO & ~ABA & ~BBA  |  ZZO & ~ABA & BBA  |  ZZI & ABA & ~BBA  |  ZZO & ABA & BBA; 
assign eba = ~EBA;  //complement 
assign EBB = ZZO & ~ABB & ~BBB  |         ZZO & ~ABB & BBB  |  ZZI & ABB & ~BBB  |  ZZO & ABB & BBB ; 
assign ebb = ~EBB;  //complement 
assign CBB =  ABA  ; 
assign cbb = ~CBB;  //complement 
assign CBC =  BBB & ABA  |  ABB  ; 
assign cbc = ~CBC;  //complement 
assign bbb = ~BBB;  //complement 
assign bbf = ~BBF;  //complement 
assign EBC = ZZO & ~ABC & ~BBC  |  ZZO & ~ABC & BBC  |  ZZI & ABC & ~BBC  |  ZZO & ABC & BBC; 
assign ebc = ~EBC;  //complement 
assign EBD = ZZO & ~ABD & ~ABD  |         ZZO & ~ABD & ABD  |  ZZI & ABD & ~ABD  |  ZZO & ABD & ABD ; 
assign ebd = ~EBD;  //complement 
assign CJD =  AJA & BJB & BJC  |  AJB & BJC  |  AJC  ; 
assign cjd = ~CJD; //complement 
assign CBD =  ABA & BBB & BBC  |  ABB & BBC  |  ABC  ; 
assign cbd = ~CBD; //complement 
assign bbc = ~BBC;  //complement 
assign bbg = ~BBG;  //complement 
assign CJB =  AJA  ; 
assign cjb = ~CJB;  //complement 
assign FAB =  BBA & BBF & BBG & BBD  ; 
assign fab = ~FAB;  //complement  
assign CBE =  ABA & BBB & BBC & BBD  |  ABB & BBC & BBD  |  ABC & BBD  |  ABD  ; 
assign cbe = ~CBE;  //complement 
assign PAB =  MAA  ; 
assign pab = ~PAB;  //complement 
assign NCA = ~nca;  //complement 
assign FAJ =  BJA & BJF & BJG & BJD  ; 
assign faj = ~FAJ;  //complement  
assign FBJ =  BJA & BJF & BJG & BJD  ; 
assign fbj = ~FBJ;  //complement 
assign kac = ~KAC;  //complement 
assign PCB =  KAC & LBC & NCA  |  KBC & NCA  |  MCA  ; 
assign pcb = ~PCB; //complement 
assign EJA = ZZO & ~AJA & ~BJA  |  ZZO & ~AJA & BJA  |  ZZI & AJA & ~BJA  |  ZZO & AJA & BJA; 
assign eja = ~EJA;  //complement 
assign EJB = ZZO & ~AJB & ~BJB  |         ZZO & ~AJB & BJB  |  ZZI & AJB & ~BJB  |  ZZO & AJB & BJB ; 
assign ejb = ~EJB;  //complement 
assign CJC =  BJB & AJA  |  AJB  ; 
assign cjc = ~CJC;  //complement 
assign bjb = ~BJB;  //complement 
assign bjf = ~BJF;  //complement 
assign EJC = ZZO & ~AJC & ~BJC  |  ZZO & ~AJC & BJC  |  ZZI & AJC & ~BJC  |  ZZO & AJC & BJC; 
assign ejc = ~EJC;  //complement 
assign EJD = ZZO & ~AJD & ~BJD  |         ZZO & ~AJD & BJD  |  ZZI & AJD & ~BJD  |  ZZO & AJD & BJD ; 
assign ejd = ~EJD;  //complement 
assign MAA = ~maa;  //complement 
assign uka = ~UKA;  //complement 
assign bjc = ~BJC;  //complement 
assign bjg = ~BJG;  //complement 
assign tdj = ~TDJ;  //complement 
assign tdb = ~TDB;  //complement 
assign MDA = ~mda;  //complement 
assign CJE =  AJA & BJB & BJC & BJD  |  AJB & BJC & BJD  |  AJC & BJD  |  AJD  ; 
assign cje = ~CJE;  //complement 
assign MCA = ~mca;  //complement 
assign ABA = ~aba;  //complement 
assign bba = ~BBA;  //complement 
assign xja = ~XJA;  //complement 
assign xjb = ~XJB;  //complement 
assign xka = ~XKA;  //complement 
assign WBA =  SBA & xba & xja  |  sba & XBA & xja  |  sba & xba & XJA  |  SBA & XBA & XJA  ; 
assign wba = ~WBA; //complement 
assign wjb =  SBA & xba & xja  |  sba & XBA & xja  |  sba & xba & XJA  |  sba & xba & xja  ; 
assign WJB = ~wjb;  //complement 
assign sba = ~SBA;  //complement 
assign sbb = ~SBB;  //complement 
assign ABB = ~abb;  //complement 
assign oae = ~OAE;  //complement 
assign oaf = ~OAF;  //complement 
assign WBB =  SBB & xbb & xjb  |  sbb & XBB & xjb  |  sbb & xbb & XJB  |  SBB & XBB & XJB  ; 
assign wbb = ~WBB; //complement 
assign wjc =  SBB & xbb & xjb  |  sbb & XBB & xjb  |  sbb & xbb & XJB  |  sbb & xbb & xjb  ; 
assign WJC = ~wjc;  //complement 
assign uba = ~UBA;  //complement 
assign ubb = ~UBB;  //complement 
assign ABC = ~abc;  //complement 
assign xbc = ~XBC;  //complement 
assign xbd = ~XBD;  //complement 
assign xjc = ~XJC;  //complement 
assign xjd = ~XJD;  //complement 
assign WBC =  SBC & xbc & xjc  |  sbc & XBC & xjc  |  sbc & xbc & XJC  |  SBC & XBC & XJC  ; 
assign wbc = ~WBC; //complement 
assign wjd =  SBC & xbc & xjc  |  sbc & XBC & xjc  |  sbc & xbc & XJC  |  sbc & xbc & xjc  ; 
assign WJD = ~wjd;  //complement 
assign sbc = ~SBC;  //complement 
assign sbd = ~SBD;  //complement 
assign ABD = ~abd;  //complement 
assign bbd = ~BBD;  //complement 
assign oag = ~OAG;  //complement 
assign oah = ~OAH;  //complement 
assign WBD =  SBD & xbd & xjd  |  sbd & XBD & xjd  |  sbd & xbd & XJD  |  SBD & XBD & XJD  ; 
assign wbd = ~WBD; //complement 
assign wka =  SBD & xbd & xjd  |  sbd & XBD & xjd  |  sbd & xbd & XJD  |  sbd & xbd & xjd  ; 
assign WKA = ~wka;  //complement 
assign ubc = ~UBC;  //complement 
assign ubd = ~UBD;  //complement 
assign AJA = ~aja;  //complement 
assign bja = ~BJA;  //complement 
assign jab =  uba & ubb & ubc & ubd  ; 
assign JAB = ~jab;  //complement  
assign tfa = ~TFA;  //complement 
assign tfb = ~TFB;  //complement 
assign tfc = ~TFC;  //complement 
assign tfd = ~TFD;  //complement 
assign sja = ~SJA;  //complement 
assign sjb = ~SJB;  //complement 
assign AJB = ~ajb;  //complement 
assign oce = ~OCE;  //complement 
assign ocf = ~OCF;  //complement 
assign uja = ~UJA;  //complement 
assign ujb = ~UJB;  //complement 
assign AJC = ~ajc;  //complement 
assign jaj =  uja & ujb & ujc & ujd  ; 
assign JAJ = ~jaj;  //complement  
assign xba = ~XBA;  //complement 
assign xbb = ~XBB;  //complement 
assign sjc = ~SJC;  //complement 
assign sjd = ~SJD;  //complement 
assign AJD = ~ajd;  //complement 
assign bjd = ~BJD;  //complement 
assign ocg = ~OCG;  //complement 
assign och = ~OCH;  //complement 
assign qbi = ~QBI;  //complement 
assign ujc = ~UJC;  //complement 
assign ujd = ~UJD;  //complement 
assign GCA = ~gca;  //complement 
assign HCA = ~hca;  //complement 
assign GCB = ~gcb;  //complement 
assign HCB = ~hcb;  //complement 
assign dcb =  bca  ; 
assign DCB = ~dcb;  //complement 
assign dcc =  acb & bca  |  bcb  ; 
assign DCC = ~dcc;  //complement 
assign HKC = ~hkc;  //complement 
assign GCC = ~gcc;  //complement 
assign HCC = ~hcc;  //complement 
assign dcd =  bca & acb & acc  |  bcb & acc  |  bcc  ; 
assign DCD = ~dcd; //complement 
assign GCD = ~gcd;  //complement 
assign HCD = ~hcd;  //complement 
assign GKA = ~gka;  //complement 
assign GKB = ~gkb;  //complement 
assign HKB = ~hkb;  //complement 
assign dkb =  bka  ; 
assign DKB = ~dkb;  //complement 
assign dkc =  akb & bka  |  bkb  ; 
assign DKC = ~dkc;  //complement 
assign GKC = ~gkc;  //complement 
assign dkd =  bka & akb & akc  |  bkb & akc  |  bkc  ; 
assign DKD = ~dkd; //complement 
assign GKD = ~gkd;  //complement 
assign HKD = ~hkd;  //complement 
assign HKA = ~hka;  //complement 
assign tdc = ~TDC;  //complement 
assign tac = ~TAC;  //complement 
assign MAB = ~mab;  //complement 
assign ECA = ZZO & ~ACA & ~BCA  |  ZZO & ~ACA & BCA  |  ZZI & ACA & ~BCA  |  ZZO & ACA & BCA; 
assign eca = ~ECA;  //complement 
assign ECB = ZZO & ~ACB & ~BCB  |         ZZO & ~ACB & BCB  |  ZZI & ACB & ~BCB  |  ZZO & ACB & BCB ; 
assign ecb = ~ECB;  //complement 
assign CCB =  ACA  ; 
assign ccb = ~CCB;  //complement 
assign CCC =  BCB & ACA  |  ACB  ; 
assign ccc = ~CCC;  //complement 
assign bcb = ~BCB;  //complement 
assign bcf = ~BCF;  //complement 
assign ECC = ZZO & ~ACC & ~BCC  |  ZZO & ~ACC & BCC  |  ZZI & ACC & ~BCC  |  ZZO & ACC & BCC; 
assign ecc = ~ECC;  //complement 
assign ECD = ZZO & ~ACD & ~BCD  |         ZZO & ~ACD & BCD  |  ZZI & ACD & ~BCD  |  ZZO & ACD & BCD ; 
assign ecd = ~ECD;  //complement 
assign CKE =  AKA & BKB & BKC & BKD  |  AKB & BKC & BKD  |  AKC & BKD  |  AKD  ; 
assign cke = ~CKE;  //complement 
assign CCD =  ACA & BCB & BCC  |  ACB & BCC  |  ACC  ; 
assign ccd = ~CCD; //complement 
assign bcc = ~BCC;  //complement 
assign bcg = ~BCG;  //complement 
assign FAC =  BCA & BCF & BCG & BCD  ; 
assign fac = ~FAC;  //complement  
assign CCE =  ACA & BCB & BCC & BCD  |  ACB & BCC & BCD  |  ACC & BCD  |  ACD  ; 
assign cce = ~CCE;  //complement 
assign PAC =  MAB  ; 
assign pac = ~PAC;  //complement 
assign NCB = ~ncb;  //complement 
assign FAK =  BKA & BKF & BKG & BKD  ; 
assign fak = ~FAK;  //complement  
assign FBK =  BKA & BKF & BKG & BKD  ; 
assign fbk = ~FBK;  //complement 
assign kad = ~KAD;  //complement 
assign PCC =  KAC & LBC & NCB  |  KBC & NCB  |  MCB  ; 
assign pcc = ~PCC; //complement 
assign EKA = ZZO & ~AKA & ~BKA  |  ZZO & ~AKA & BKA  |  ZZI & AKA & ~BKA  |  ZZO & AKA & BKA; 
assign eka = ~EKA;  //complement 
assign EKB = ZZO & ~AKB & ~BKB  |         ZZO & ~AKB & BKB  |  ZZI & AKB & ~BKB  |  ZZO & AKB & BKB ; 
assign ekb = ~EKB;  //complement 
assign CKB =  AKA  ; 
assign ckb = ~CKB;  //complement 
assign CKC =  BKB & AKA  |  AKB  ; 
assign ckc = ~CKC;  //complement 
assign bkb = ~BKB;  //complement 
assign bkf = ~BKF;  //complement 
assign EKC = ZZO & ~AKC & ~BKC  |  ZZO & ~AKC & BKC  |  ZZI & AKC & ~BKC  |  ZZO & AKC & BKC; 
assign ekc = ~EKC;  //complement 
assign EKD = ZZO & ~AKD & ~BKD  |         ZZO & ~AKD & BKD  |  ZZI & AKD & ~BKD  |  ZZO & AKD & BKD ; 
assign ekd = ~EKD;  //complement 
assign CKD =  AKA & BKB & BKC  |  AKB & BKC  |  AKC  ; 
assign ckd = ~CKD; //complement 
assign bkc = ~BKC;  //complement 
assign bkg = ~BKG;  //complement 
assign tdk = ~TDK;  //complement 
assign MCB = ~mcb;  //complement 
assign ACA = ~aca;  //complement 
assign xca = ~XCA;  //complement 
assign xcb = ~XCB;  //complement 
assign xkb = ~XKB;  //complement 
assign WCA =  SCA & xca & xka  |  sca & XCA & xka  |  sca & xca & XKA  |  SCA & XCA & XKA  ; 
assign wca = ~WCA; //complement 
assign wkb =  SCA & xca & xka  |  sca & XCA & xka  |  sca & xca & XKA  |  sca & xca & xka  ; 
assign WKB = ~wkb;  //complement 
assign scb = ~SCB;  //complement 
assign ACB = ~acb;  //complement 
assign oai = ~OAI;  //complement 
assign oaj = ~OAJ;  //complement 
assign WCB =  SCB & xcb & xkb  |  scb & XCB & xkb  |  scb & xcb & XKB  |  SCB & XCB & XKB  ; 
assign wcb = ~WCB; //complement 
assign wkc =  SCB & xcb & xkb  |  scb & XCB & xkb  |  scb & xcb & XKB  |  scb & xcb & xkb  ; 
assign WKC = ~wkc;  //complement 
assign uca = ~UCA;  //complement 
assign ucb = ~UCB;  //complement 
assign ACC = ~acc;  //complement 
assign xcc = ~XCC;  //complement 
assign xcd = ~XCD;  //complement 
assign xkc = ~XKC;  //complement 
assign xkd = ~XKD;  //complement 
assign WCC =  SCC & xcc & xkc  |  scc & XCC & xkc  |  scc & xcc & XKC  |  SCC & XCC & XKC  ; 
assign wcc = ~WCC; //complement 
assign wkd =  SCC & xcc & xkc  |  scc & XCC & xkc  |  scc & xcc & XKC  |  scc & xcc & xkc  ; 
assign WKD = ~wkd;  //complement 
assign scc = ~SCC;  //complement 
assign scd = ~SCD;  //complement 
assign ACD = ~acd;  //complement 
assign bcd = ~BCD;  //complement 
assign oak = ~OAK;  //complement 
assign oal = ~OAL;  //complement 
assign WCD =  SCD & xcd & xkd  |  scd & XCD & xkd  |  scd & xcd & XKD  |  SCD & XCD & XKD  ; 
assign wcd = ~WCD; //complement 
assign wla =  SCD & xcd & xkd  |  scd & XCD & xkd  |  scd & xcd & XKD  |  scd & xcd & xkd  ; 
assign WLA = ~wla;  //complement 
assign ucc = ~UCC;  //complement 
assign ucd = ~UCD;  //complement 
assign bka = ~BKA;  //complement 
assign jac =  uca & ucb & ucc & ucd  ; 
assign JAC = ~jac;  //complement  
assign tga = ~TGA;  //complement 
assign tgb = ~TGB;  //complement 
assign tgc = ~TGC;  //complement 
assign tgd = ~TGD;  //complement 
assign ska = ~SKA;  //complement 
assign skb = ~SKB;  //complement 
assign AKB = ~akb;  //complement 
assign oci = ~OCI;  //complement 
assign ocj = ~OCJ;  //complement 
assign qjb = ~QJB;  //complement 
assign ukb = ~UKB;  //complement 
assign AKC = ~akc;  //complement 
assign jak =  uka & ukb & ukc & ukd  ; 
assign JAK = ~jak;  //complement  
assign qbd = ~QBD;  //complement 
assign skc = ~SKC;  //complement 
assign skd = ~SKD;  //complement 
assign AKD = ~akd;  //complement 
assign bkd = ~BKD;  //complement 
assign ock = ~OCK;  //complement 
assign ocl = ~OCL;  //complement 
assign qca = ~QCA;  //complement 
assign qcb = ~QCB;  //complement 
assign ukc = ~UKC;  //complement 
assign ukd = ~UKD;  //complement 
assign GDA = ~gda;  //complement 
assign HDA = ~hda;  //complement 
assign GDB = ~gdb;  //complement 
assign HDB = ~hdb;  //complement 
assign ddb =  bda  ; 
assign DDB = ~ddb;  //complement 
assign ddc =  adb & bda  |  bdb  ; 
assign DDC = ~ddc;  //complement 
assign HLC = ~hlc;  //complement 
assign GDC = ~gdc;  //complement 
assign HDC = ~hdc;  //complement 
assign ddd =  bda & adb & adc  |  bdb & adc  |  bdc  ; 
assign DDD = ~ddd; //complement 
assign HLB = ~hlb;  //complement 
assign GDD = ~gdd;  //complement 
assign HDD = ~hdd;  //complement 
assign GLA = ~gla;  //complement 
assign HLA = ~hla;  //complement 
assign GLB = ~glb;  //complement 
assign dlb =  bla  ; 
assign DLB = ~dlb;  //complement 
assign dlc =  alb & bla  |  blb  ; 
assign DLC = ~dlc;  //complement 
assign GLC = ~glc;  //complement 
assign dld =  bla & alb & alc  |  blb & alc  |  blc  ; 
assign DLD = ~dld; //complement 
assign GLD = ~gld;  //complement 
assign HLD = ~hld;  //complement 
assign tdd = ~TDD;  //complement 
assign tad = ~TAD;  //complement 
assign MAC = ~mac;  //complement 
assign EDA = ZZO & ~ADA & ~BDA  |  ZZO & ~ADA & BDA  |  ZZI & ADA & ~BDA  |  ZZO & ADA & BDA; 
assign eda = ~EDA;  //complement 
assign EDB = ZZO & ~ADB & ~BDB  |         ZZO & ~ADB & BDB  |  ZZI & ADB & ~BDB  |  ZZO & ADB & BDB ; 
assign edb = ~EDB;  //complement 
assign CDB =  ADA  ; 
assign cdb = ~CDB;  //complement 
assign CDC =  BDB & ADA  |  ADB  ; 
assign cdc = ~CDC;  //complement 
assign bdb = ~BDB;  //complement 
assign bdf = ~BDF;  //complement 
assign EDC = ZZO & ~ADC & ~BDC  |  ZZO & ~ADC & BDC  |  ZZI & ADC & ~BDC  |  ZZO & ADC & BDC; 
assign edc = ~EDC;  //complement 
assign EDD = ZZO & ~ADD & ~BDD  |         ZZO & ~ADD & BDD  |  ZZI & ADD & ~BDD  |  ZZO & ADD & BDD ; 
assign edd = ~EDD;  //complement 
assign CLD =  ALA & BLB & BLC  |  ALB & BLC  |  ALC  ; 
assign cld = ~CLD; //complement 
assign CDD =  ADA & BDB & BDC  |  ADB & BDC  |  ADC  ; 
assign cdd = ~CDD; //complement 
assign bdc = ~BDC;  //complement 
assign bdg = ~BDG;  //complement 
assign FAD =  BDA & BDF & BDG & BDD  ; 
assign fad = ~FAD;  //complement  
assign CDE =  ADA & BDB & BDC & BDD  |  ADB & BDC & BDD  |  ADC & BDD  |  ADD  ; 
assign cde = ~CDE;  //complement 
assign PAD =  MAC  ; 
assign pad = ~PAD;  //complement 
assign NCC = ~ncc;  //complement 
assign FAL =  BLA & BLF & BLG & BLD  ; 
assign fal = ~FAL;  //complement  
assign kbc = ~KBC;  //complement 
assign PCD =  KAC & LBC & NCC  |  KBC & NCC  |  MCC  ; 
assign pcd = ~PCD; //complement 
assign ELA = ZZO & ~ALA & ~BLA  |  ZZO & ~ALA & BLA  |  ZZI & ALA & ~BLA  |  ZZO & ALA & BLA; 
assign ela = ~ELA;  //complement 
assign ELB = ZZO & ~ALB & ~BLB  |         ZZO & ~ALB & BLB  |  ZZI & ALB & ~BLB  |  ZZO & ALB & BLB ; 
assign elb = ~ELB;  //complement 
assign BLG =  ULC  |  SLC  ; 
assign blg = ~BLG;  //complement 
assign CLB =  ALA  ; 
assign clb = ~CLB;  //complement 
assign CLC =  BLB & ALA  |  ALB  ; 
assign clc = ~CLC;  //complement 
assign blb = ~BLB;  //complement 
assign blf = ~BLF;  //complement 
assign ELC = ZZO & ~ALC & ~BLC  |  ZZO & ~ALC & BLC  |  ZZI & ALC & ~BLC  |  ZZO & ALC & BLC; 
assign elc = ~ELC;  //complement 
assign ELD = ZZO & ~ALD & ~BLD  |         ZZO & ~ALD & BLD  |  ZZI & ALD & ~BLD  |  ZZO & ALD & BLD ; 
assign eld = ~ELD;  //complement 
assign blc = ~BLC;  //complement 
assign tdl = ~TDL;  //complement 
assign CLE =  ALA & BLB & BLC & BLD  |  ALB & BLC & BLD  |  ALC & BLD  |  ALD  ; 
assign cle = ~CLE;  //complement 
assign MCC = ~mcc;  //complement 
assign ADA = ~ada;  //complement 
assign bda = ~BDA;  //complement 
assign xda = ~XDA;  //complement 
assign xdb = ~XDB;  //complement 
assign xla = ~XLA;  //complement 
assign xlb = ~XLB;  //complement 
assign WDA =  SDA & xda & xla  |  sda & XDA & xla  |  sda & xda & XLA  |  SDA & XDA & XLA  ; 
assign wda = ~WDA; //complement 
assign wlb =  SDA & xda & xla  |  sda & XDA & xla  |  sda & xda & XLA  |  sda & xda & xla  ; 
assign WLB = ~wlb;  //complement 
assign sda = ~SDA;  //complement 
assign sdb = ~SDB;  //complement 
assign ADB = ~adb;  //complement 
assign ADC = ~adc;  //complement 
assign oam = ~OAM;  //complement 
assign oan = ~OAN;  //complement 
assign WDB =  SDB & xdb & xlb  |  sdb & XDB & xlb  |  sdb & xdb & XLB  |  SDB & XDB & XLB  ; 
assign wdb = ~WDB; //complement 
assign wlc =  SDB & xdb & xlb  |  sdb & XDB & xlb  |  sdb & xdb & XLB  |  sdb & xdb & xlb  ; 
assign WLC = ~wlc;  //complement 
assign uda = ~UDA;  //complement 
assign udb = ~UDB;  //complement 
assign xdc = ~XDC;  //complement 
assign xdd = ~XDD;  //complement 
assign xlc = ~XLC;  //complement 
assign xld = ~XLD;  //complement 
assign WDC =  SDC & xdc & xlc  |  sdc & XDC & xlc  |  sdc & xdc & XLC  |  SDC & XDC & XLC  ; 
assign wdc = ~WDC; //complement 
assign wld =  SDC & xdc & xlc  |  sdc & XDC & xlc  |  sdc & xdc & XLC  |  sdc & xdc & xlc  ; 
assign WLD = ~wld;  //complement 
assign sdc = ~SDC;  //complement 
assign sdd = ~SDD;  //complement 
assign ADD = ~add;  //complement 
assign bdd = ~BDD;  //complement 
assign oao = ~OAO;  //complement 
assign oap = ~OAP;  //complement 
assign WDD =  SDD & xdd & xld  |  sdd & XDD & xld  |  sdd & xdd & XLD  |  SDD & XDD & XLD  ; 
assign wdd = ~WDD; //complement 
assign wma =  SDD & xdd & xld  |  sdd & XDD & xld  |  sdd & xdd & XLD  |  sdd & xdd & xld  ; 
assign WMA = ~wma;  //complement 
assign udc = ~UDC;  //complement 
assign udd = ~UDD;  //complement 
assign ALA = ~ala;  //complement 
assign bla = ~BLA;  //complement 
assign jad =  uda & udb & udc & udd  ; 
assign JAD = ~jad;  //complement  
assign jqa =  qaa & qad  ; 
assign JQA = ~jqa;  //complement 
assign QAA = ~qaa;  //complement 
assign qab = ~QAB;  //complement 
assign qac = ~QAC;  //complement 
assign QAD = ~qad;  //complement 
assign sla = ~SLA;  //complement 
assign slb = ~SLB;  //complement 
assign ALB = ~alb;  //complement 
assign ocm = ~OCM;  //complement 
assign ocn = ~OCN;  //complement 
assign qbe = ~QBE;  //complement 
assign qbf = ~QBF;  //complement 
assign ula = ~ULA;  //complement 
assign ulb = ~ULB;  //complement 
assign ALC = ~alc;  //complement 
assign jal =  ula & ulb & ulc & uld  ; 
assign JAL = ~jal;  //complement  
assign JDA =  QBE & qbf  ; 
assign jda = ~JDA;  //complement 
assign qbb = ~QBB;  //complement 
assign slc = ~SLC;  //complement 
assign sld = ~SLD;  //complement 
assign ALD = ~ald;  //complement 
assign bld = ~BLD;  //complement 
assign oco = ~OCO;  //complement 
assign ocp = ~OCP;  //complement 
assign QBA = ~qba;  //complement 
assign QBC = ~qbc;  //complement 
assign ulc = ~ULC;  //complement 
assign uld = ~ULD;  //complement 
assign GEA = ~gea;  //complement 
assign HEA = ~hea;  //complement 
assign GEB = ~geb;  //complement 
assign HEB = ~heb;  //complement 
assign deb =  bea  ; 
assign DEB = ~deb;  //complement 
assign dec =  aeb & bea  |  beb  ; 
assign DEC = ~dec;  //complement 
assign GMC = ~gmc;  //complement 
assign HMC = ~hmc;  //complement 
assign GEC = ~gec;  //complement 
assign HEC = ~hec;  //complement 
assign bec = ~BEC;  //complement 
assign GED = ~ged;  //complement 
assign HED = ~hed;  //complement 
assign GMA = ~gma;  //complement 
assign HMA = ~hma;  //complement 
assign GMB = ~gmb;  //complement 
assign HMB = ~hmb;  //complement 
assign dmb =  bma  ; 
assign DMB = ~dmb;  //complement 
assign dmc =  amb & bma  |  bmb  ; 
assign DMC = ~dmc;  //complement 
assign ded =  bea & aeb & aec  |  beb & aec  |  bec  ; 
assign DED = ~ded; //complement 
assign HMD = ~hmd;  //complement 
assign GMD = ~gmd;  //complement 
assign dmd =  bma & amb & amc  |  bmb & amc  |  bmc  ; 
assign DMD = ~dmd; //complement 
assign tde = ~TDE;  //complement 
assign tae = ~TAE;  //complement 
assign EEA = ZZO & ~AEA & ~BEA  |  ZZO & ~AEA & BEA  |  ZZI & AEA & ~BEA  |  ZZO & AEA & BEA; 
assign eea = ~EEA;  //complement 
assign EEB = ZZO & ~AEB & ~BEB  |         ZZO & ~AEB & BEB  |  ZZI & AEB & ~BEB  |  ZZO & AEB & BEB ; 
assign eeb = ~EEB;  //complement 
assign CEB =  AEA  ; 
assign ceb = ~CEB;  //complement 
assign CEC =  BEB & AEA  |  AEB  ; 
assign cec = ~CEC;  //complement 
assign beb = ~BEB;  //complement 
assign bef = ~BEF;  //complement 
assign EEC = ZZO & ~AEC & ~BEC  |  ZZO & ~AEC & BEC  |  ZZI & AEC & ~BEC  |  ZZO & AEC & BEC; 
assign eec = ~EEC;  //complement 
assign EED = ZZO & ~AED & ~BED  |         ZZO & ~AED & BED  |  ZZI & AED & ~BED  |  ZZO & AED & BED ; 
assign eed = ~EED;  //complement 
assign CMD =  AMA & BMB & BMC  |  AMB & BMC  |  AMC  ; 
assign cmd = ~CMD; //complement 
assign CED =  AEA & BEB & BEC  |  AEB & BEC  |  AEC  ; 
assign ced = ~CED; //complement 
assign beg = ~BEG;  //complement 
assign FAE =  BEA & BEF & BEG & BED  ; 
assign fae = ~FAE;  //complement  
assign CEE =  AEA & BEB & BEC & BED  |  AEB & BEC & BED  |  AEC & BED  |  AED  ; 
assign cee = ~CEE;  //complement 
assign pba =  kab  ; 
assign PBA = ~pba;  //complement 
assign FAM =  BMA & BMF & BMG & BMD  ; 
assign fam = ~FAM;  //complement  
assign kbd = ~KBD;  //complement 
assign PDA =  KAD & LBD & LCD  |  KBD & LCD  |  KCD  ; 
assign pda = ~PDA;  //complement 
assign EMA = ZZO & ~AMA & ~BMA  |  ZZO & ~AMA & BMA  |  ZZI & AMA & ~BMA  |  ZZO & AMA & BMA; 
assign ema = ~EMA;  //complement 
assign EMB = ZZO & ~AMB & ~BMB  |         ZZO & ~AMB & BMB  |  ZZI & AMB & ~BMB  |  ZZO & AMB & BMB ; 
assign emb = ~EMB;  //complement 
assign CMB =  AMA  ; 
assign cmb = ~CMB;  //complement 
assign CMC =  BMB & AMA  |  AMB  ; 
assign cmc = ~CMC;  //complement 
assign bmb = ~BMB;  //complement 
assign bmf = ~BMF;  //complement 
assign EMC = ZZO & ~AMC & ~BMC  |  ZZO & ~AMC & BMC  |  ZZI & AMC & ~BMC  |  ZZO & AMC & BMC; 
assign emc = ~EMC;  //complement 
assign EMD = ZZO & ~AMD & ~BMD  |         ZZO & ~AMD & BMD  |  ZZI & AMD & ~BMD  |  ZZO & AMD & BMD ; 
assign emd = ~EMD;  //complement 
assign bmc = ~BMC;  //complement 
assign bmg = ~BMG;  //complement 
assign tdm = ~TDM;  //complement 
assign CME =  AMA & BMB & BMC & BMD  |  AMB & BMC & BMD  |  AMC & BMD  |  AMD  ; 
assign cme = ~CME;  //complement 
assign AEA = ~aea;  //complement 
assign bea = ~BEA;  //complement 
assign xea = ~XEA;  //complement 
assign xeb = ~XEB;  //complement 
assign xma = ~XMA;  //complement 
assign xmb = ~XMB;  //complement 
assign WEA =  SEA & xea & xma  |  sea & XEA & xma  |  sea & xea & XMA  |  SEA & XEA & XMA  ; 
assign wea = ~WEA; //complement 
assign wmb =  SEA & xea & xma  |  sea & XEA & xma  |  sea & xea & XMA  |  sea & xea & xma  ; 
assign WMB = ~wmb;  //complement 
assign sea = ~SEA;  //complement 
assign seb = ~SEB;  //complement 
assign AEB = ~aeb;  //complement 
assign AEC = ~aec;  //complement 
assign oba = ~OBA;  //complement 
assign obb = ~OBB;  //complement 
assign WEB =  SEB & xeb & xmb  |  seb & XEB & xmb  |  seb & xeb & XMB  |  SEB & XEB & XMB  ; 
assign web = ~WEB; //complement 
assign wmc =  SEB & xeb & xmb  |  seb & XEB & xmb  |  seb & xeb & XMB  |  seb & xeb & xmb  ; 
assign WMC = ~wmc;  //complement 
assign uea = ~UEA;  //complement 
assign ueb = ~UEB;  //complement 
assign xec = ~XEC;  //complement 
assign xed = ~XED;  //complement 
assign xmc = ~XMC;  //complement 
assign xmd = ~XMD;  //complement 
assign WEC =  SEC & xec & xmc  |  sec & XEC & xmc  |  sec & xec & XMC  |  SEC & XEC & XMC  ; 
assign wec = ~WEC; //complement 
assign wmd =  SEC & xec & xmc  |  sec & XEC & xmc  |  sec & xec & XMC  |  sec & xec & xmc  ; 
assign WMD = ~wmd;  //complement 
assign sec = ~SEC;  //complement 
assign sed = ~SED;  //complement 
assign AED = ~aed;  //complement 
assign bed = ~BED;  //complement 
assign obc = ~OBC;  //complement 
assign obd = ~OBD;  //complement 
assign WED =  SED & xed & xmd  |  sed & XED & xmd  |  sed & xed & XMD  |  SED & XED & XMD  ; 
assign wed = ~WED; //complement 
assign wna =  SED & xed & xmd  |  sed & XED & xmd  |  sed & xed & XMD  |  sed & xed & xmd  ; 
assign WNA = ~wna;  //complement 
assign uec = ~UEC;  //complement 
assign ued = ~UED;  //complement 
assign AMA = ~ama;  //complement 
assign bma = ~BMA;  //complement 
assign jae =  uea & ueb & uec & ued  ; 
assign JAE = ~jae;  //complement  
assign ona = ~ONA;  //complement 
assign qna = ~QNA;  //complement 
assign qnb = ~QNB;  //complement 
assign qnc = ~QNC;  //complement 
assign sma = ~SMA;  //complement 
assign smb = ~SMB;  //complement 
assign AMB = ~amb;  //complement 
assign oda = ~ODA;  //complement 
assign odb = ~ODB;  //complement 
assign qjc = ~QJC;  //complement 
assign uma = ~UMA;  //complement 
assign umb = ~UMB;  //complement 
assign AMC = ~amc;  //complement 
assign jam =  uma & umb & umc & umd  ; 
assign JAM = ~jam;  //complement  
assign jbb =  qja & qjb & qjc & qjd & qje  ; 
assign JBB = ~jbb;  //complement  
assign jba =  qja & qjb & qjc & qjd  ; 
assign JBA = ~jba;  //complement 
assign smc = ~SMC;  //complement 
assign smd = ~SMD;  //complement 
assign AMD = ~amd;  //complement 
assign bmd = ~BMD;  //complement 
assign odc = ~ODC;  //complement 
assign odd = ~ODD;  //complement 
assign umc = ~UMC;  //complement 
assign umd = ~UMD;  //complement 
assign GFA = ~gfa;  //complement 
assign HFA = ~hfa;  //complement 
assign GFB = ~gfb;  //complement 
assign HFB = ~hfb;  //complement 
assign dfc =  afb & bfa  |  bfb  ; 
assign DFC = ~dfc;  //complement 
assign DFB = ~dfb;  //complement 
assign HNC = ~hnc;  //complement 
assign GFC = ~gfc;  //complement 
assign HFC = ~hfc;  //complement 
assign dfd =  bfa & afb & afc  |  bfb & afc  |  bfc  ; 
assign DFD = ~dfd; //complement 
assign GFD = ~gfd;  //complement 
assign HFD = ~hfd;  //complement 
assign GNA = ~gna;  //complement 
assign HNA = ~hna;  //complement 
assign GNB = ~gnb;  //complement 
assign HNB = ~hnb;  //complement 
assign dnb =  bna  ; 
assign DNB = ~dnb;  //complement 
assign dnc =  anb & bna  |  bnb  ; 
assign DNC = ~dnc;  //complement 
assign GNC = ~gnc;  //complement 
assign dnd =  bna & anb & anc  |  bnb & anc  |  bnc  ; 
assign DND = ~dnd; //complement 
assign GND = ~gnd;  //complement 
assign HND = ~hnd;  //complement 
assign tdf = ~TDF;  //complement 
assign qee = ~QEE;  //complement 
assign qef = ~QEF;  //complement 
assign taf = ~TAF;  //complement 
assign MBA = ~mba;  //complement 
assign EFA = ZZO & ~AFA & ~BFA  |  ZZO & ~AFA & BFA  |  ZZI & AFA & ~BFA  |  ZZO & AFA & BFA; 
assign efa = ~EFA;  //complement 
assign EFB = ZZO & ~AFB & ~BFB  |         ZZO & ~AFB & BFB  |  ZZI & AFB & ~BFB  |  ZZO & AFB & BFB ; 
assign efb = ~EFB;  //complement 
assign CFB =  AFA  ; 
assign cfb = ~CFB;  //complement 
assign CFC =  BFB & AFA  |  AFB  ; 
assign cfc = ~CFC;  //complement 
assign bfb = ~BFB;  //complement 
assign bff = ~BFF;  //complement 
assign EFC = ZZO & ~AFC & ~BFC  |  ZZO & ~AFC & BFC  |  ZZI & AFC & ~BFC  |  ZZO & AFC & BFC; 
assign efc = ~EFC;  //complement 
assign EFD = ZZO & ~AFD & ~BFD  |         ZZO & ~AFD & BFD  |  ZZI & AFD & ~BFD  |  ZZO & AFD & BFD ; 
assign efd = ~EFD;  //complement 
assign CND =  ANA & BNB & BNC  |  ANB & BNC  |  ANC  ; 
assign cnd = ~CND; //complement 
assign CFD =  AFA & BFB & BFC  |  AFB & BFC  |  AFC  ; 
assign cfd = ~CFD; //complement 
assign bfc = ~BFC;  //complement 
assign bfg = ~BFG;  //complement 
assign NBA = ~nba;  //complement 
assign FAF =  BFA & BFF & BFG & BFD  ; 
assign faf = ~FAF;  //complement  
assign FBF =  BFA & BFF & BFG & BFD  ; 
assign fbf = ~FBF;  //complement 
assign CFE =  AFA & BFB & BFC & BFD  |  AFB & BFC & BFD  |  AFC & BFD  |  AFD  ; 
assign cfe = ~CFE;  //complement 
assign PBB =  KAB & NBA  |  MBA  ; 
assign pbb = ~PBB; //complement 
assign NDA = ~nda;  //complement 
assign FAN =  BNA & BNF & BNG & BND  ; 
assign fan = ~FAN;  //complement  
assign FBN =  BNA & BNF & BNG & BND  ; 
assign fbn = ~FBN;  //complement 
assign kcd = ~KCD;  //complement 
assign PDB =  KAD & LBD & LCD & NDA  |  KBD & LCD & NDA  |  KCD & NDA  |  MDA  ; 
assign pdb = ~PDB;  //complement 
assign ENA = ZZO & ~ANA & ~BNA  |  ZZO & ~ANA & BNA  |  ZZI & ANA & ~BNA  |  ZZO & ANA & BNA; 
assign ena = ~ENA;  //complement 
assign ENB = ZZO & ~ANB & ~BNB  |         ZZO & ~ANB & BNB  |  ZZI & ANB & ~BNB  |  ZZO & ANB & BNB ; 
assign enb = ~ENB;  //complement 
assign CNB =  ANA  ; 
assign cnb = ~CNB;  //complement 
assign CNC =  BNB & ANA  |  ANB  ; 
assign cnc = ~CNC;  //complement 
assign bnf = ~BNF;  //complement 
assign bnb = ~BNB;  //complement 
assign ENC = ZZO & ~ANC & ~BNC  |  ZZO & ~ANC & BNC  |  ZZI & ANC & ~BNC  |  ZZO & ANC & BNC; 
assign enc = ~ENC;  //complement 
assign ENDD  = ZZO & ~ANDD  & ~BND  |         ZZO & ~ANDD  & BND  |  ZZI & ANDD  & ~BND  |  ZZO & ANDD  & BND ; 
assign endd = ~ENDD ;  //complement 
assign bnc = ~BNC;  //complement 
assign bng = ~BNG;  //complement 
assign tdn = ~TDN;  //complement 
assign CNE =  ANA & BNB & BNC & BND  |  ANB & BNC & BND  |  ANC & BND  |  ANDD   ; 
assign cne = ~CNE;  //complement 
assign AFA = ~afa;  //complement 
assign bfa = ~BFA;  //complement 
assign xfa = ~XFA;  //complement 
assign xfb = ~XFB;  //complement 
assign xna = ~XNA;  //complement 
assign xnb = ~XNB;  //complement 
assign WFA =  SFA & xfa & xna  |  sfa & XFA & xna  |  sfa & xfa & XNA  |  SFA & XFA & XNA  ; 
assign wfa = ~WFA; //complement 
assign wnb =  SFA & xfa & xna  |  sfa & XFA & xna  |  sfa & xfa & XNA  |  sfa & xfa & xna  ; 
assign WNB = ~wnb;  //complement 
assign sfa = ~SFA;  //complement 
assign sfb = ~SFB;  //complement 
assign AFB = ~afb;  //complement 
assign obe = ~OBE;  //complement 
assign obf = ~OBF;  //complement 
assign WFB =  SFB & xfb & xnb  |  sfb & XFB & xnb  |  sfb & xfb & XNB  |  SFB & XFB & XNB  ; 
assign wfb = ~WFB; //complement 
assign wnc =  SFB & xfb & xnb  |  sfb & XFB & xnb  |  sfb & xfb & XNB  |  sfb & xfb & xnb  ; 
assign WNC = ~wnc;  //complement 
assign ufa = ~UFA;  //complement 
assign ufb = ~UFB;  //complement 
assign AFC = ~afc;  //complement 
assign xfc = ~XFC;  //complement 
assign xfd = ~XFD;  //complement 
assign xnc = ~XNC;  //complement 
assign xnd = ~XND;  //complement 
assign WFC =  SFC & xfc & xnc  |  sfc & XFC & xnc  |  sfc & xfc & XNC  |  SFC & XFC & XNC  ; 
assign wfc = ~WFC; //complement 
assign wnd =  SFC & xfc & xnc  |  sfc & XFC & xnc  |  sfc & xfc & XNC  |  sfc & xfc & xnc  ; 
assign WND = ~wnd;  //complement 
assign sfc = ~SFC;  //complement 
assign sfd = ~SFD;  //complement 
assign AFD = ~afd;  //complement 
assign bfd = ~BFD;  //complement 
assign obg = ~OBG;  //complement 
assign obh = ~OBH;  //complement 
assign WFD =  SFD & xfd & xnd  |  sfd & XFD & xnd  |  sfd & xfd & XND  |  SFD & XFD & XND  ; 
assign wfd = ~WFD; //complement 
assign woa =  SFD & xfd & xnd  |  sfd & XFD & xnd  |  sfd & xfd & XND  |  sfd & xfd & xnd  ; 
assign WOA = ~woa;  //complement 
assign ufc = ~UFC;  //complement 
assign ufd = ~UFD;  //complement 
assign ANA = ~ana;  //complement 
assign bna = ~BNA;  //complement 
assign jaf =  ufa & ufb & ufc & ufd  ; 
assign JAF = ~jaf;  //complement  
assign THA = ~tha;  //complement 
assign THB = ~thb;  //complement 
assign THC = ~thc;  //complement 
assign THD = ~thd;  //complement 
assign sna = ~SNA;  //complement 
assign snb = ~SNB;  //complement 
assign ANB = ~anb;  //complement 
assign ode = ~ODE;  //complement 
assign odf = ~ODF;  //complement 
assign OEA = ~oea;  //complement 
assign una = ~UNA;  //complement 
assign unb = ~UNB;  //complement 
assign ANC = ~anc;  //complement 
assign jan =  una & unb & unc & und  ; 
assign JAN = ~jan;  //complement  
assign QGA = ~qga;  //complement 
assign QGB = ~qgb;  //complement 
assign snc = ~SNC;  //complement 
assign snd = ~SND;  //complement 
assign ANDD  = ~andd ;  //complement 
assign bnd = ~BND;  //complement 
assign odg = ~ODG;  //complement 
assign odh = ~ODH;  //complement 
assign QEA = ~qea;  //complement 
assign qeb = ~QEB;  //complement 
assign qec = ~QEC;  //complement 
assign qed = ~QED;  //complement 
assign unc = ~UNC;  //complement 
assign und = ~UND;  //complement 
assign GGA = ~gga;  //complement 
assign HGA = ~hga;  //complement 
assign GGB = ~ggb;  //complement 
assign HGB = ~hgb;  //complement 
assign dgb =  bga  ; 
assign DGB = ~dgb;  //complement 
assign dgc =  agb & bga  |  bgb  ; 
assign DGC = ~dgc;  //complement 
assign HOC = ~hoc;  //complement 
assign GGC = ~ggc;  //complement 
assign HGC = ~hgc;  //complement 
assign dgd =  bga & agb & agc  |  bgb & agc  |  bgc  ; 
assign DGD = ~dgd; //complement 
assign HOB = ~hob;  //complement 
assign GGD = ~ggd;  //complement 
assign HGD = ~hgd;  //complement 
assign GOA = ~goa;  //complement 
assign HOA = ~hoa;  //complement 
assign GOB = ~gob;  //complement 
assign dob =  boa  ; 
assign DOB = ~dob;  //complement 
assign doc =  aob & boa  |  bob  ; 
assign DOC = ~doc;  //complement 
assign GOC = ~goc;  //complement 
assign dod =  boa & aob & aoc  |  bob & aoc  |  boc  ; 
assign DOD = ~dod; //complement 
assign GOD = ~god;  //complement 
assign HOD = ~hod;  //complement 
assign tdg = ~TDG;  //complement 
assign qcf = ~QCF;  //complement 
assign tag = ~TAG;  //complement 
assign MBB = ~mbb;  //complement 
assign EGA = ZZO & ~AGA & ~BGA  |  ZZO & ~AGA & BGA  |  ZZI & AGA & ~BGA  |  ZZO & AGA & BGA; 
assign ega = ~EGA;  //complement 
assign EGB = ZZO & ~AGB & ~BGB  |         ZZO & ~AGB & BGB  |  ZZI & AGB & ~BGB  |  ZZO & AGB & BGB ; 
assign egb = ~EGB;  //complement 
assign CGB =  AGA  ; 
assign cgb = ~CGB;  //complement 
assign CGC =  BGB & AGA  |  AGB  ; 
assign cgc = ~CGC;  //complement 
assign bgb = ~BGB;  //complement 
assign bgf = ~BGF;  //complement 
assign EGC = ZZO & ~AGC & ~BGC  |  ZZO & ~AGC & BGC  |  ZZI & AGC & ~BGC  |  ZZO & AGC & BGC; 
assign egc = ~EGC;  //complement 
assign EGD = ZZO & ~AGD & ~BGD  |         ZZO & ~AGD & BGD  |  ZZI & AGD & ~BGD  |  ZZO & AGD & BGD ; 
assign egd = ~EGD;  //complement 
assign COD =  AOA & BOB & BOC  |  AOB & BOC  |  AOC  ; 
assign cod = ~COD; //complement 
assign CGD =  AGA & BGB & BGC  |  AGB & BGC  |  AGC  ; 
assign cgd = ~CGD; //complement 
assign bgc = ~BGC;  //complement 
assign bgg = ~BGG;  //complement 
assign NBB = ~nbb;  //complement 
assign FAG =  BGA & BGF & BGG & BGD  ; 
assign fag = ~FAG;  //complement  
assign FBG =  BGA & BGF & BGG & BGD  ; 
assign fbg = ~FBG;  //complement 
assign CGE =  AGA & BGB & BGC & BGD  |  AGB & BGC & BGD  |  AGC & BGD  |  AGD  ; 
assign cge = ~CGE;  //complement 
assign PBC =  KAB & NBB  |  MBB  ; 
assign pbc = ~PBC; //complement 
assign NDB = ~ndb;  //complement 
assign FAO =  BOA & BOF & BOG & BOD  ; 
assign fao = ~FAO;  //complement  
assign FBO =  BOA & BOF & BOG & BOD  ; 
assign fbo = ~FBO;  //complement 
assign LCD = ~lcd;  //complement 
assign PDC =  KAD & LBD & LCD & NDB  |  KBD & LCD & NDB  |  KCD & NDB  |  MDB  ; 
assign pdc = ~PDC;  //complement 
assign EOA = ZZO & ~AOA & ~BOA  |  ZZO & ~AOA & BOA  |  ZZI & AOA & ~BOA  |  ZZO & AOA & BOA; 
assign eoa = ~EOA;  //complement 
assign EOB = ZZO & ~AOB & ~BOB  |         ZZO & ~AOB & BOB  |  ZZI & AOB & ~BOB  |  ZZO & AOB & BOB ; 
assign eob = ~EOB;  //complement 
assign COB =  AOA  ; 
assign cob = ~COB;  //complement 
assign COC =  BOB & AOA  |  AOB  ; 
assign coc = ~COC;  //complement 
assign bob = ~BOB;  //complement 
assign bof = ~BOF;  //complement 
assign EOC = ZZO & ~AOC & ~BOC  |  ZZO & ~AOC & BOC  |  ZZI & AOC & ~BOC  |  ZZO & AOC & BOC; 
assign eoc = ~EOC;  //complement 
assign EOD = ZZO & ~AOD & ~BOD  |         ZZO & ~AOD & BOD  |  ZZI & AOD & ~BOD  |  ZZO & AOD & BOD ; 
assign eod = ~EOD;  //complement 
assign boc = ~BOC;  //complement 
assign bog = ~BOG;  //complement 
assign tdo = ~TDO;  //complement 
assign AKA = ~aka;  //complement 
assign COE =  AOA & BOB & BOC & BOD  |  AOB & BOC & BOD  |  AOC & BOD  |  AOD  ; 
assign coe = ~COE;  //complement 
assign MDB = ~mdb;  //complement 
assign AGA = ~aga;  //complement 
assign bga = ~BGA;  //complement 
assign xga = ~XGA;  //complement 
assign xgb = ~XGB;  //complement 
assign xoa = ~XOA;  //complement 
assign xob = ~XOB;  //complement 
assign WGA =  SGA & xga & xoa  |  sga & XGA & xoa  |  sga & xga & XOA  |  SGA & XGA & XOA  ; 
assign wga = ~WGA; //complement 
assign wob =  SGA & xga & xoa  |  sga & XGA & xoa  |  sga & xga & XOA  |  sga & xga & xoa  ; 
assign WOB = ~wob;  //complement 
assign sga = ~SGA;  //complement 
assign sgb = ~SGB;  //complement 
assign AGB = ~agb;  //complement 
assign obi = ~OBI;  //complement 
assign obj = ~OBJ;  //complement 
assign WGB =  SGB & xgb & xob  |  sgb & XGB & xob  |  sgb & xgb & XOB  |  SGB & XGB & XOB  ; 
assign wgb = ~WGB; //complement 
assign woc =  SGB & xgb & xob  |  sgb & XGB & xob  |  sgb & xgb & XOB  |  sgb & xgb & xob  ; 
assign WOC = ~woc;  //complement 
assign uga = ~UGA;  //complement 
assign ugb = ~UGB;  //complement 
assign AGC = ~agc;  //complement 
assign xgc = ~XGC;  //complement 
assign xgd = ~XGD;  //complement 
assign xoc = ~XOC;  //complement 
assign xod = ~XOD;  //complement 
assign WGC =  SGC & xgc & xoc  |  sgc & XGC & xoc  |  sgc & xgc & XOC  |  SGC & XGC & XOC  ; 
assign wgc = ~WGC; //complement 
assign wod =  SGC & xgc & xoc  |  sgc & XGC & xoc  |  sgc & xgc & XOC  |  sgc & xgc & xoc  ; 
assign WOD = ~wod;  //complement 
assign sgc = ~SGC;  //complement 
assign sgd = ~SGD;  //complement 
assign AGD = ~agd;  //complement 
assign bgd = ~BGD;  //complement 
assign obk = ~OBK;  //complement 
assign obl = ~OBL;  //complement 
assign WGD =  SGD & xgd & xod  |  sgd & XGD & xod  |  sgd & xgd & XOD  |  SGD & XGD & XOD  ; 
assign wgd = ~WGD; //complement 
assign wpa =  SGD & xgd & xod  |  sgd & XGD & xod  |  sgd & xgd & XOD  |  sgd & xgd & xod  ; 
assign WPA = ~wpa;  //complement 
assign ugc = ~UGC;  //complement 
assign ugd = ~UGD;  //complement 
assign AOA = ~aoa;  //complement 
assign boa = ~BOA;  //complement 
assign jag =  uga & ugb & ugc & ugd  ; 
assign JAG = ~jag;  //complement  
assign tia = ~TIA;  //complement 
assign tib = ~TIB;  //complement 
assign tic = ~TIC;  //complement 
assign tid = ~TID;  //complement 
assign soa = ~SOA;  //complement 
assign sob = ~SOB;  //complement 
assign AOB = ~aob;  //complement 
assign odi = ~ODI;  //complement 
assign odj = ~ODJ;  //complement 
assign qjd = ~QJD;  //complement 
assign uoa = ~UOA;  //complement 
assign uob = ~UOB;  //complement 
assign AOC = ~aoc;  //complement 
assign qcg = ~QCG;  //complement 
assign jao =  uoa & uob & uoc & uod  ; 
assign JAO = ~jao;  //complement  
assign qce = ~QCE;  //complement 
assign qfa = ~QFA;  //complement 
assign qfb = ~QFB;  //complement 
assign soc = ~SOC;  //complement 
assign sod = ~SOD;  //complement 
assign AOD = ~aod;  //complement 
assign bod = ~BOD;  //complement 
assign odk = ~ODK;  //complement 
assign odl = ~ODL;  //complement 
assign qje = ~QJE;  //complement 
assign uoc = ~UOC;  //complement 
assign uod = ~UOD;  //complement 
assign GHA = ~gha;  //complement 
assign HHA = ~hha;  //complement 
assign GHB = ~ghb;  //complement 
assign HHB = ~hhb;  //complement 
assign dhb =  bha  ; 
assign DHB = ~dhb;  //complement 
assign dhc =  ahb & bha  |  bhb  ; 
assign DHC = ~dhc;  //complement 
assign HPC = ~hpc;  //complement 
assign GHC = ~ghc;  //complement 
assign HHC = ~hhc;  //complement 
assign dhd =  bha & ahb & ahc  |  bhb & ahc  |  bhc  ; 
assign DHD = ~dhd; //complement 
assign HPB = ~hpb;  //complement 
assign GHD = ~ghd;  //complement 
assign HHD = ~hhd;  //complement 
assign GPA = ~gpa;  //complement 
assign HPA = ~hpa;  //complement 
assign CPB =  APA  ; 
assign cpb = ~CPB;  //complement 
assign GPB = ~gpb;  //complement 
assign dpb =  bpa  ; 
assign DPB = ~dpb;  //complement 
assign dpc =  apb & bpa  |  bpb  ; 
assign DPC = ~dpc;  //complement 
assign GPC = ~gpc;  //complement 
assign dpd =  bpa & apb & apc  |  bpb & apc  |  bpc  ; 
assign DPD = ~dpd; //complement 
assign GPD = ~gpd;  //complement 
assign HPD = ~hpd;  //complement 
assign tdh = ~TDH;  //complement 
assign tah = ~TAH;  //complement 
assign MBC = ~mbc;  //complement 
assign EHA = ZZO & ~AHA & ~BHA  |  ZZO & ~AHA & BHA  |  ZZI & AHA & ~BHA  |  ZZO & AHA & BHA; 
assign eha = ~EHA;  //complement 
assign EHB = ZZO & ~AHB & ~BHB  |         ZZO & ~AHB & BHB  |  ZZI & AHB & ~BHB  |  ZZO & AHB & BHB ; 
assign ehb = ~EHB;  //complement 
assign CHB =  AHA  ; 
assign chb = ~CHB;  //complement 
assign CHC =  BHB & AHA  |  AHB  ; 
assign chc = ~CHC;  //complement 
assign bhb = ~BHB;  //complement 
assign bhf = ~BHF;  //complement 
assign EHC = ZZO & ~AHC & ~BHC  |  ZZO & ~AHC & BHC  |  ZZI & AHC & ~BHC  |  ZZO & AHC & BHC; 
assign ehc = ~EHC;  //complement 
assign EHD = ZZO & ~AHD & ~BHD  |         ZZO & ~AHD & BHD  |  ZZI & AHD & ~BHD  |  ZZO & AHD & BHD ; 
assign ehd = ~EHD;  //complement 
assign CPD =  APA & BPB & BPC  |  APB & BPC  |  APC  ; 
assign cpd = ~CPD; //complement 
assign CHD =  AHA & BHB & BHC  |  AHB & BHC  |  AHC  ; 
assign chd = ~CHD; //complement 
assign bhc = ~BHC;  //complement 
assign bhg = ~BHG;  //complement 
assign NBC = ~nbc;  //complement 
assign FAH =  BHA & BHF & BHG & BHD  ; 
assign fah = ~FAH;  //complement  
assign CHE =  AHA & BHB & BHC & BHD  |  AHB & BHC & BHD  |  AHC & BHD  |  AHD  ; 
assign che = ~CHE;  //complement 
assign PBD =  KAB & NBC  |  MBC  ; 
assign pbd = ~PBD; //complement 
assign NDC = ~ndc;  //complement 
assign LBC = ~lbc;  //complement 
assign LBD = ~lbd;  //complement 
assign PDD =  KAD & LBD & LCD & NDC  |  KBD & LCD & NDC  |  KCD & NDC  |  MDC  ; 
assign pdd = ~PDD;  //complement 
assign EPA = ZZO & ~APA & ~BPA  |  ZZO & ~APA & BPA  |  ZZI & APA & ~BPA  |  ZZO & APA & BPA; 
assign epa = ~EPA;  //complement 
assign EPB = ZZO & ~APB & ~BPB  |         ZZO & ~APB & BPB  |  ZZI & APB & ~BPB  |  ZZO & APB & BPB ; 
assign epb = ~EPB;  //complement 
assign CPC =  BPB & APA  |  APB  ; 
assign cpc = ~CPC;  //complement 
assign EPC = ZZO & ~APC & ~BPC  |  ZZO & ~APC & BPC  |  ZZI & APC & ~BPC  |  ZZO & APC & BPC; 
assign epc = ~EPC;  //complement 
assign EPD = ZZO & ~APD & ~BPD  |         ZZO & ~APD & BPD  |  ZZI & APD & ~BPD  |  ZZO & APD & BPD ; 
assign epd = ~EPD;  //complement 
assign tdp = ~TDP;  //complement 
assign MDC = ~mdc;  //complement 
assign AHA = ~aha;  //complement 
assign bha = ~BHA;  //complement 
assign xha = ~XHA;  //complement 
assign xhb = ~XHB;  //complement 
assign xpa = ~XPA;  //complement 
assign xpb = ~XPB;  //complement 
assign WHA =  SHA & xha & xpa  |  sha & XHA & xpa  |  sha & xha & XPA  |  SHA & XHA & XPA  ; 
assign wha = ~WHA; //complement 
assign wpb =  SHA & xha & xpa  |  sha & XHA & xpa  |  sha & xha & XPA  |  sha & xha & xpa  ; 
assign WPB = ~wpb;  //complement 
assign sha = ~SHA;  //complement 
assign shb = ~SHB;  //complement 
assign AHB = ~ahb;  //complement 
assign obm = ~OBM;  //complement 
assign obn = ~OBN;  //complement 
assign WHB =  SHB & xhb & xpb  |  shb & XHB & xpb  |  shb & xhb & XPB  |  SHB & XHB & XPB  ; 
assign whb = ~WHB; //complement 
assign wpc =  SHB & xhb & xpb  |  shb & XHB & xpb  |  shb & xhb & XPB  |  shb & xhb & xpb  ; 
assign WPC = ~wpc;  //complement 
assign uha = ~UHA;  //complement 
assign uhb = ~UHB;  //complement 
assign AHC = ~ahc;  //complement 
assign xhc = ~XHC;  //complement 
assign xhd = ~XHD;  //complement 
assign xpc = ~XPC;  //complement 
assign xpd = ~XPD;  //complement 
assign WHC =  SHC & xhc & xpc  |  shc & XHC & xpc  |  shc & xhc & XPC  |  SHC & XHC & XPC  ; 
assign whc = ~WHC; //complement 
assign wpd =  SHC & xhc & xpc  |  shc & XHC & xpc  |  shc & xhc & XPC  |  shc & xhc & xpc  ; 
assign WPD = ~wpd;  //complement 
assign shc = ~SHC;  //complement 
assign shd = ~SHD;  //complement 
assign AHD = ~ahd;  //complement 
assign bhd = ~BHD;  //complement 
assign obo = ~OBO;  //complement 
assign obp = ~OBP;  //complement 
assign WHD =  SHD & xhd & xpd  |  shd & XHD & xpd  |  shd & xhd & XPD  |  SHD & XHD & XPD  ; 
assign whd = ~WHD; //complement 
assign uhc = ~UHC;  //complement 
assign uhd = ~UHD;  //complement 
assign APA = ~apa;  //complement 
assign bpa = ~BPA;  //complement 
assign jah =  uha & uhb & uhc & uhd  ; 
assign JAH = ~jah;  //complement  
assign TJA = ~tja;  //complement 
assign TJB = ~tjb;  //complement 
assign TJC = ~tjc;  //complement 
assign TJD = ~tjd;  //complement 
assign spa = ~SPA;  //complement 
assign spb = ~SPB;  //complement 
assign APB = ~apb;  //complement 
assign bpb = ~BPB;  //complement 
assign odm = ~ODM;  //complement 
assign odn = ~ODN;  //complement 
assign oeb = ~OEB;  //complement 
assign oec = ~OEC;  //complement 
assign upa = ~UPA;  //complement 
assign upb = ~UPB;  //complement 
assign APC = ~apc;  //complement 
assign bpc = ~BPC;  //complement 
assign jap =  upa & upb & upc  ; 
assign JAP = ~jap;  //complement  
assign ofa = ~OFA;  //complement 
assign ofb = ~OFB;  //complement 
assign spc = ~SPC;  //complement 
assign spd = ~SPD;  //complement 
assign APD = ~apd;  //complement 
assign bpd = ~BPD;  //complement 
assign odo = ~ODO;  //complement 
assign odp = ~ODP;  //complement 
assign qha = ~QHA;  //complement 
assign upe = ~UPE;  //complement 
assign upc = ~UPC;  //complement 
assign upd = ~UPD;  //complement 
assign iaa = ~IAA; //complement 
assign iab = ~IAB; //complement 
assign iac = ~IAC; //complement 
assign iad = ~IAD; //complement 
assign iae = ~IAE; //complement 
assign iaf = ~IAF; //complement 
assign iag = ~IAG; //complement 
assign iah = ~IAH; //complement 
assign iai = ~IAI; //complement 
assign iaj = ~IAJ; //complement 
assign iak = ~IAK; //complement 
assign ial = ~IAL; //complement 
assign iam = ~IAM; //complement 
assign ian = ~IAN; //complement 
assign iao = ~IAO; //complement 
assign iap = ~IAP; //complement 
assign iba = ~IBA; //complement 
assign ibb = ~IBB; //complement 
assign ibc = ~IBC; //complement 
assign ibd = ~IBD; //complement 
assign ibe = ~IBE; //complement 
assign ibf = ~IBF; //complement 
assign ibg = ~IBG; //complement 
assign ibh = ~IBH; //complement 
assign ibi = ~IBI; //complement 
assign ibj = ~IBJ; //complement 
assign ibk = ~IBK; //complement 
assign ibl = ~IBL; //complement 
assign ibm = ~IBM; //complement 
assign ibn = ~IBN; //complement 
assign ibo = ~IBO; //complement 
assign ibp = ~IBP; //complement 
assign ica = ~ICA; //complement 
assign icb = ~ICB; //complement 
assign icc = ~ICC; //complement 
assign icd = ~ICD; //complement 
assign ice = ~ICE; //complement 
assign icf = ~ICF; //complement 
assign icg = ~ICG; //complement 
assign ich = ~ICH; //complement 
assign ici = ~ICI; //complement 
assign icj = ~ICJ; //complement 
assign ick = ~ICK; //complement 
assign icl = ~ICL; //complement 
assign icm = ~ICM; //complement 
assign icn = ~ICN; //complement 
assign ico = ~ICO; //complement 
assign icp = ~ICP; //complement 
assign ida = ~IDA; //complement 
assign idb = ~IDB; //complement 
assign idc = ~IDC; //complement 
assign idd = ~IDD; //complement 
assign ide = ~IDE; //complement 
assign idf = ~IDF; //complement 
assign idg = ~IDG; //complement 
assign idh = ~IDH; //complement 
assign idi = ~IDI; //complement 
assign idj = ~IDJ; //complement 
assign idk = ~IDK; //complement 
assign idl = ~IDL; //complement 
assign idm = ~IDM; //complement 
assign idn = ~IDN; //complement 
assign ido = ~IDO; //complement 
assign idp = ~IDP; //complement 
assign iea = ~IEA; //complement 
assign ieb = ~IEB; //complement 
assign iec = ~IEC; //complement 
assign ied = ~IED; //complement 
assign iee = ~IEE; //complement 
assign ief = ~IEF; //complement 
assign ieg = ~IEG; //complement 
assign ieh = ~IEH; //complement 
assign iei = ~IEI; //complement 
assign iej = ~IEJ; //complement 
assign iek = ~IEK; //complement 
assign iel = ~IEL; //complement 
assign iem = ~IEM; //complement 
assign ien = ~IEN; //complement 
assign ieo = ~IEO; //complement 
assign iep = ~IEP; //complement 
assign ifa = ~IFA; //complement 
assign ifb = ~IFB; //complement 
assign ifc = ~IFC; //complement 
assign ifd = ~IFD; //complement 
assign ife = ~IFE; //complement 
assign ifff  = ~IFFF ; //complement 
assign ifg = ~IFG; //complement 
assign ifh = ~IFH; //complement 
assign ifi = ~IFI; //complement 
assign ifj = ~IFJ; //complement 
assign ifk = ~IFK; //complement 
assign ifl = ~IFL; //complement 
assign ifm = ~IFM; //complement 
assign ifn = ~IFN; //complement 
assign ifo = ~IFO; //complement 
assign ifp = ~IFP; //complement 
assign iga = ~IGA; //complement 
assign igb = ~IGB; //complement 
assign igc = ~IGC; //complement 
assign igd = ~IGD; //complement 
assign ige = ~IGE; //complement 
assign igf = ~IGF; //complement 
assign igg = ~IGG; //complement 
assign igh = ~IGH; //complement 
assign igi = ~IGI; //complement 
assign igj = ~IGJ; //complement 
assign igk = ~IGK; //complement 
assign igl = ~IGL; //complement 
assign igm = ~IGM; //complement 
assign ign = ~IGN; //complement 
assign igo = ~IGO; //complement 
assign igp = ~IGP; //complement 
assign iha = ~IHA; //complement 
assign ihb = ~IHB; //complement 
assign ihc = ~IHC; //complement 
assign ihd = ~IHD; //complement 
assign ihe = ~IHE; //complement 
assign ihf = ~IHF; //complement 
assign ihg = ~IHG; //complement 
assign ihh = ~IHH; //complement 
assign ihi = ~IHI; //complement 
assign ihj = ~IHJ; //complement 
assign ihk = ~IHK; //complement 
assign ihl = ~IHL; //complement 
assign ihm = ~IHM; //complement 
assign ihn = ~IHN; //complement 
assign iho = ~IHO; //complement 
assign ihp = ~IHP; //complement 
assign ima = ~IMA; //complement 
assign ira = ~IRA; //complement 
assign irb = ~IRB; //complement 
assign irc = ~IRC; //complement 
assign ird = ~IRD; //complement 
always@(posedge IZZ )
   begin 
 gaa <=  caa & eaa  |  CAA & EAA  |  tda  ; 
 gab <=  cab & eab  |  CAB & EAB  |  tda  ; 
 hic <=  dic & eic  |  DIC & EEC  |  tdi  ; 
 gac <=  cac & eac  |  CAC & EAC  |  tda  ; 
 gad <=  cad & ead  |  CAD & EAD  |  tda  ; 
 gia <=  eia  |  tdi  ; 
 hia <=  EIA  |  tdi  ; 
 hib <=  dib & eib  |  DIB & EIB  |  tdi  ; 
 gib <=  cib & eib  |  CIB & EIB  |  tdi  ; 
 gic <=  cic & eic  |  CIC & EIC  |  tdi  ; 
 gid <=  cid & eid  |  CID & EID  |  tdi  ; 
 hid <=  did & eid  |  DID & EID  |  tdi  ; 
 TDA <= qef ; 
 TAA <= QCF ; 
 tka <= qib ; 
 tkb <= qib ; 
 QFC <= QFB ; 
 QFD <= QFC ; 
 QIA <= JCA ; 
 QIB <= QIA ; 
 KAB <=  CAE & FAB & FAC & FAD  |  CBE & FAC & FAD  |  CCE & FAD  |  CDE  ; 
 BIB <=  UIB  |  SIB  ; 
 BIF <=  UIB  |  SIB  ; 
 BIC <=  UIC  |  SIC  ; 
 BIG <=  UIC  |  SIC  ; 
 QDE <= QDD ; 
 TDI <= qde ; 
 aaa <=  uaa & TAA  |  waa  |  taa  ; 
 BAA <=  UAA & TAA  |  WAA  ; 
 XAA <= TKA & WAA ; 
 XAB <= TKA & WAB ; 
 XIB <= TKA & WIB ; 
 SAA <=  SAA & TEA  |  IAA & TFA  |  IEA & TGA  ; 
 SAB <=  SAB & TEA  |  IAB & TFA  |  IEB & TGA  ; 
 aab <=  uab & TAA  |  wab  |  wib & taa  ; 
 aac <=  uac & TAA  |  wac  |  wic & taa  ; 
 OAA <=  GAA  ; 
 OAB <=  GAB  ; 
 UAA <=  iea & THA  |  ZZI & TIA  |  IEA & TJA  ; 
 UAB <=  ieb & THA  |  UAA & TIA  |  IEB & TJA  ; 
 BAC <=  UAC & TAA  |  WAC  |  WIC & taa  ; 
 XAC <= TKB & WAC ; 
 XAD <= TKB & WAD ; 
 XIC <= TKB & WIC ; 
 XID <= TKB & WID ; 
 SAC <=  SAC & TEB  |  IAC & TFB  |  IEC & TGB  ; 
 SAD <=  SAD & TEB  |  IAD & TFB  |  IED & TGB  ; 
 aad <=  uad & TAA  |  wad  |  wid & taa  ; 
 BAD <=  UAD & TAA  |  WAD  |  WID & taa  ; 
 OAC <=  GAC  ; 
 OAD <=  GAD  ; 
 UAC <=  iec & THB  |  UAB & TIB  |  IEC & TJB  ; 
 UAD <=  ied & THB  |  UAC & TIB  |  IED & TJB  ; 
 aia <=  uia  |  sia  ; 
 BIA <=  UIA  |  SIA  ; 
 TEA <= qcb & qca ; 
 TEB <= qcb & qca ; 
 TEC <= qcb & qca ; 
 TED <= qcb & qca ; 
 SIA <=  SIA & TEC  |  ICA & TFC  |  IGA & TGC  ; 
 SIB <=  SIB & TEC  |  ICB & TFC  |  IGB & TGC  ; 
 aib <=  uib  |  sib  ; 
 OCA <=  GIA & pca  |  HEA & PCA  ; 
 OCB <=  GEB & pca  |  HIB & PCA  ; 
 QJA <=  JAA  |  JAB  |  JAE  |  JAJ  ; 
 UIB <=  igb & THC  |  UIA & TIC  |  IGB & TJC  ; 
 UIA <=  iga & THC  |  UHD & TIC  |  IGA & TJC  ; 
 aic <=  uic  |  sic  ; 
 BAB <=  UAB & TAA  |  WAB  |  WIB & taa  ; 
 SIC <=  SIC & TED  |  ICC & TFD  |  IGC & TGD  ; 
 SID <=  SID & TED  |  ICD & TFD  |  IGD & TGD  ; 
 aid <=  uid  |  sid  ; 
 BID <=  UID  |  SID  ; 
 OCC <=  GEC & pca  |  HIC & PCA  ; 
 OCD <=  GID & pca  |  HID & PCA  ; 
 QDA <= QBI ; 
 QDB <= QDA ; 
 QDC <= QDB ; 
 QDD <= QDC ; 
 UIC <=  igc & THD  |  UIB & TID  |  IGC & TJD  ; 
 UID <=  igd & THD  |  UIC & TID  |  IGD & TJD  ; 
 gba <=  eba  |  tdb  ; 
 hba <=  EBA  |  tdb  ; 
 gbb <=  cbb & ebb  |  CBB & EBB  |  tdb  ; 
 hbb <=  dbb & ebb  |  DBB & EBB  |  tdb  ; 
 hjc <=  djc & ejc  |  DJC & EJC  |  tdj  ; 
 gbc <=  cbc & ebc  |  CBC & EBC  |  tdb  ; 
 hbc <=  dbc & ebc  |  DBC & EBC  |  tdb  ; 
 gbd <=  cbd & ebd  |  CBD & EBD  |  tdb  ; 
 hbd <=  dbd & ebd  |  DBD & EBD  |  tdb  ; 
 gja <=  eja  |  tdj  ; 
 hja <=  EJA  |  tdj  ; 
 hjb <=  djb & ejb  |  DJB & EJB  |  tdj  ; 
 gjb <=  cjb & ejb  |  CJB & EJB  |  tdj  ; 
 gjc <=  cjc & ejc  |  CJC & EJC  |  tdj  ; 
 gjd <=  cjd & ejd  |  CJD & EJD  |  tdj  ; 
 hjd <=  djd & ejd  |  DJD & EJD  |  tdj  ; 
 BCA <=  UCA & TAC  |  WCA  |  WKA & tac  ; 
 TAB <= QCF ; 
 SCA <=  SCA & TEA  |  IAI & TFA  |  IEI & TGA  ; 
 BBB <=  UBB & TAB  |  WBB  |  WJB & tab  ; 
 BBF <=  UBB & TAB  |  WBB  |  WJB & tab  ; 
 BBC <=  UBC & TAB  |  WBC  |  WJC & tab  ; 
 BBG <=  UBC & TAB  |  WBC  |  WJC & tab  ; 
 nca <=  fai  ; 
 KAC <=  CAE & FAB & FAC & FAD  |  CBE & FAC & FAD  |  CCE & FAD  |  CDE  ; 
 BJB <=  UJB  |  SJB  ; 
 BJF <=  UJB  |  SJB  ; 
 maa <=  cae  ; 
 UKA <=  igi & THC  |  UJD & TIC  |  IGI & TJC  ; 
 BJC <=  UJC  |  SJC  ; 
 BJG <=  UJC  |  SJC  ; 
 TDJ <= qde ; 
 TDB <= qef ; 
 mda <=  cme  ; 
 mca <=  cie  ; 
 aba <=  uba & TAB  |  wba  |  wja & tab  ; 
 BBA <=  UBA & TAB  |  WBA  |  WJA & tab  ; 
 XJA <= TKA & WJA ; 
 XJB <= TKA & WJB ; 
 XKA <= TKA & WKA ; 
 SBA <=  SBA & TEA  |  IAE & TFA  |  IEE & TGA  ; 
 SBB <=  SBB & TEA  |  IAF & TFA  |  IEF & TGA  ; 
 abb <=  ubb & TAB  |  wbb  |  wjb & tab  ; 
 OAE <=  GBA & pab  |  HBA & PAB  ; 
 OAF <=  GBB & pab  |  HBB & PAB  ; 
 UBA <=  iee & THA  |  UAD & TIA  |  IEE & TJA  ; 
 UBB <=  ief & THA  |  UBA & TIA  |  IEF & TJA  ; 
 abc <=  ubc & TAB  |  wbc  |  wjc & tab  ; 
 XBC <= TKB & WBC ; 
 XBD <= TKB & WBD ; 
 XJC <= TKB & WJC ; 
 XJD <= TKB & WJD ; 
 SBC <=  SBC & TEB  |  IAG & TFB  |  IEG & TGB  ; 
 SBD <=  SBD & TEB  |  IAH & TFB  |  IEH & TGB  ; 
 abd <=  ubd & TAB  |  wbd  |  wjd & tab  ; 
 BBD <=  UBD & TAB  |  WBD  |  WJD & tab  ; 
 OAG <=  GBC & pab  |  HBC & PAB  ; 
 OAH <=  GBD & pab  |  HBD & PAB  ; 
 UBC <=  ieg & THB  |  UBB & TIB  |  IEG & TJB  ; 
 UBD <=  ieh & THB  |  UBC & TIB  |  IEH & TJB  ; 
 aja <=  uja  |  sja  ; 
 BJA <=  UJA  |  SJA  ; 
 TFA <= QCA ; 
 TFB <= QCA ; 
 TFC <= QCA ; 
 TFD <= QCA ; 
 SJA <=  SJA & TEC  |  ICE & TFC  |  IGE & TGC  ; 
 SJB <=  SJB & TEC  |  ICF & TFC  |  IGF & TGC  ; 
 ajb <=  ujb  |  sjb  ; 
 OCE <=  GJA & pcb  |  HJA & PCB  ; 
 OCF <=  GJB & pcb  |  HJB & PCB  ; 
 UJA <=  ige & THC  |  UID & TIC  |  IGE & TJC  ; 
 UJB <=  igf & THC  |  UJA & TIC  |  IGF & TJC  ; 
 ajc <=  ujc  |  sjc  ; 
 XBA <= TKA & WBA ; 
 XBB <= TKA & WBB ; 
 SJC <=  SJC & TED  |  ICG & TFD  |  IGG & TGD  ; 
 SJD <=  SJD & TED  |  ICH & TFD  |  IGH & TGD  ; 
 ajd <=  ujd  |  sjd  ; 
 BJD <=  UJD  |  SJD  ; 
 OCG <=  GJC & pcb  |  HJC & PCB  ; 
 OCH <=  GJD & pcb  |  HJD & PCB  ; 
 QBI <=  QBI & jqa  |  QAD  ; 
 UJC <=  igg & THD  |  UJB & TID  |  IGG & TJD  ; 
 UJD <=  igh & THD  |  UJC & TID  |  IGH & TJD  ; 
 gca <=  eca  |  tdc  ; 
 hca <=  ECA  |  tdc  ; 
 gcb <=  ccb & ecb  |  CCB & ECB  |  tdc  ; 
 hcb <=  dcb & ecb  |  DCB & ECB  |  tdc  ; 
 hkc <=  dkc & ekc  |  DKC & EKC  |  tdk  ; 
 gcc <=  ccc & ecc  |  CCC & ECC  |  tdc  ; 
 hcc <=  dcc & ecc  |  DCC & ECC  |  tdc  ; 
 gcd <=  ccd & ecd  |  CCD & ECD  |  tdc  ; 
 hcd <=  dcd & ecd  |  DCD & ECD  |  tdc  ; 
 gka <=  eka & ekb  |  tdk & EKB  ; 
 gkb <=  ckb & ekb  |  CKB & EKB  |  tdk  ; 
 hkb <=  dkb & ekb  |  DKB & EKB  |  tdk  ; 
 gkc <=  ckc & ekc  |  CKC & EKC  |  tdk  ; 
 gkd <=  ckd & ekd  |  CKD & EKD  |  tdk  ; 
 hkd <=  dkd & ekd  |  DKD & EKD  |  tdk  ; 
 hka <=  EKA  |  tdk  ; 
 TDC <= qef ; 
 TAC <= QCF ; 
 mab <=  cae & cbe & cbe  |  fab & cbe  ; 
 BCB <=  UCB & TAC  |  WCB  |  WKB & tac  ; 
 BCF <=  UCB & TAC  |  WCB  |  WKB & tac  ; 
 BCC <=  UCC & TAC  |  WCC  |  WKC & tac  ; 
 BCG <=  UCC & TAC  |  WCC  |  WKC & tac  ; 
 ncb <=  fai  |  faj  ; 
 KAD <=  CAE & FAB & FAC & FAD  |  CBE & FAC & FAD  |  CCE & FAD  |  CDE  ; 
 BKB <=  UKB  |  SKB  ; 
 BKF <=  UKB  |  SKB  ; 
 BKC <=  UKC  |  SKC  ; 
 BKG <=  UKC  |  SKC  ; 
 TDK <= qde ; 
 mcb <=  cie & cje & cje  |  fbj & cje  ; 
 aca <=  uca & TAC  |  wca  |  wka & tac  ; 
 XCA <= TKA & WCA ; 
 XCB <= TKA & WCB ; 
 XKB <= TKA & WKB ; 
 SCB <=  SCB & TEA  |  IAJ & TFA  |  IEJ & TGA  ; 
 acb <=  ucb & TAC  |  wcb  |  wkb & tac  ; 
 OAI <=  GCA & pac  |  HCA & PAC  ; 
 OAJ <=  GCB & pac  |  HCB & PAC  ; 
 UCA <=  iei & THA  |  UBD & TIA  |  IEI & TJA  ; 
 UCB <=  iej & THA  |  UCA & TIA  |  IEJ & TJA  ; 
 acc <=  ucc & TAC  |  wcc  |  wkc & tac  ; 
 XCC <= TKB & WCC ; 
 XCD <= TKB & WCD ; 
 XKC <= TKB & WKC ; 
 XKD <= TKB & WKD ; 
 SCC <=  SCC & TEB  |  IAK & TFB  |  IEK & TGB  ; 
 SCD <=  SCD & TEB  |  IAL & TFB  |  IEL & TGB  ; 
 acd <=  ucd & TAC  |  wcd  |  wkd & tac  ; 
 BCD <=  UCD & TAC  |  WCD  |  WKD & tac  ; 
 OAK <=  GCC & pac  |  HCC & PAC  ; 
 OAL <=  GCD & pac  |  HCD & PAC  ; 
 UCC <=  iek & THB  |  UCB & TIB  |  IEK & TJB  ; 
 UCD <=  iel & THB  |  UCC & TIB  |  IEL & TJB  ; 
 BKA <=  UKA  |  SKA  ; 
 TGA <= QCB ; 
 TGB <= QCB ; 
 TGC <= QCB ; 
 TGD <= QCB ; 
 SKA <=  SKA & TEC  |  ICI & TFC  |  IGI & TGC  ; 
 SKB <=  SKB & TEC  |  ICJ & TFC  |  IGJ & TGC  ; 
 akb <=  ukb  |  skb  ; 
 OCI <=  GKA & pcc  |  HKA & PCC  ; 
 OCJ <=  GKB & pcc  |  HKB & PCC  ; 
 QJB <=  JAC  |  JAD  |  JAK  |  JAL  ; 
 UKB <=  igj & THC  |  UKA & TIC  |  IGJ & TJC  ; 
 akc <=  ukc  |  skc  ; 
 QBD <=  QAC & QAB & QAA  |  QBD & jqa  ; 
 SKC <=  SKC & TED  |  ICK & TFD  |  IGK & TGD  ; 
 SKD <=  SKD & TED  |  ICL & TFD  |  IGL & TGD  ; 
 akd <=  ukd  |  skd  ; 
 BKD <=  UKD  |  SKD  ; 
 OCK <=  GKC & pcc  |  HKC & PCC  ; 
 OCL <=  GKD & pcc  |  HKD & PCC  ; 
 QCA <=  QBB  |  QBD  ; 
 QCB <=  QBA  |  QBC  |  QEB  ; 
 UKC <=  igk & THD  |  UKB & TID  |  IGK & TJD  ; 
 UKD <=  igl & THD  |  UKC & TID  |  IGL & TJD  ; 
 gda <=  eda  |  tdd  ; 
 hda <=  EDA  |  tdd  ; 
 gdb <=  cdb & edb  |  CDB & EDB  |  tdd  ; 
 hdb <=  ddb & edb  |  DDB & EDB  |  tdd  ; 
 hlc <=  dlc & elc  |  DLC & ELC  |  tdl  ; 
 gdc <=  cdc & edc  |  CDC & EDC  |  tdd  ; 
 hdc <=  ddc & edc  |  DDC & EDC  |  tdd  ; 
 hlb <=  dlb & elb  |  DLB & ELB  |  tdl  ; 
 gdd <=  cdd & edd  |  CDD & EDD  |  tdd  ; 
 hdd <=  ddd & edd  |  DDD & EDD  |  tdd  ; 
 gla <=  ela  |  tdl  ; 
 hla <=  ELA  |  tdl  ; 
 glb <=  clb & elb  |  CLB & ELB  |  tdl  ; 
 glc <=  clc & elc  |  CLC & ELC  |  tdl  ; 
 gld <=  cld & eld  |  CLD & ELD  |  tdl  ; 
 hld <=  dld & eld  |  DLD & ELD  |  tdl  ; 
 TDD <= qef ; 
 TAD <= QCF ; 
 mac <=  ZZI & cae & cbe & cce  |  ZZI & cae & cbe & cce  |  fab & cbe & cce  |  ZZI & fac & cce  ; 
 BDB <=  UDB & TAD  |  WDB  |  WLB & tad  ; 
 BDF <=  UDB & TAD  |  WDB  |  WLB & tad  ; 
 BDC <=  UDC & TAD  |  WDC  |  WLC & tad  ; 
 BDG <=  UDC & TAD  |  WDC  |  WLC & tad  ; 
 ncc <=  fai  |  faj  |  fak  ; 
 KBC <=  CEE & FAF & FAG & FAH  |  CFE & FAG & FAH  |  CGE & FAH  |  CHE  ; 
 BLB <=  ULB  |  SLB  ; 
 BLF <=  ULB  |  SLB  ; 
 BLC <=  ULC  |  SLC  ; 
 TDL <= qde ; 
 mcc <=  ZZI & cie & cje & cke  |  ZZI & cie & cje & cke  |  fbj & cje & cke  |  ZZI & fbk & cke  ; 
 ada <=  uda & TAD  |  wda  |  wla & tad  ; 
 BDA <=  UDA & TAD  |  WDA  |  WLA & tad  ; 
 XDA <= TKA & WDA ; 
 XDB <= TKA & WDB ; 
 XLA <= TKA & WLA ; 
 XLB <= TKA & WLB ; 
 SDA <=  SDA & TEA  |  IAM & TFA  |  IEM & TGA  ; 
 SDB <=  SDB & TEA  |  IAN & TFA  |  IEN & TGA  ; 
 adb <=  udb & TAD  |  wdb  |  wlb & tad  ; 
 adc <=  udc & TAD  |  wdc  |  wlc & tad  ; 
 OAM <=  GDA & pad  |  HDA & PAD  ; 
 OAN <=  GDB & pad  |  HDB & PAD  ; 
 UDA <=  iem & THA  |  UCD & TIA  |  IEM & TJA  ; 
 UDB <=  ien & THA  |  UDA & TIA  |  IEN & TJA  ; 
 XDC <= TKB & WDC ; 
 XDD <= TKB & WDD ; 
 XLC <= TKB & WLC ; 
 XLD <= TKB & WLD ; 
 SDC <=  SDC & TEB  |  IAO & TFB  |  IEO & TGB  ; 
 SDD <=  SDD & TEB  |  IAP & TFB  |  IEP & TGB  ; 
 add <=  udd & TAD  |  wdd  |  wld & tad  ; 
 BDD <=  UDD & TAD  |  WDD  |  WLD & tad  ; 
 OAO <=  GDC & pad  |  HDC & PAD  ; 
 OAP <=  GDD & pad  |  HDD & PAD  ; 
 UDC <=  ieo & THB  |  UDB & TIB  |  IEO & TJB  ; 
 UDD <=  iep & THB  |  UDC & TIB  |  IEP & TJB  ; 
 ala <=  ula  |  sla  ; 
 BLA <=  ULA  |  SLA  ; 
 qaa <= ira ; 
 QAB <= IRB ; 
 QAC <= IRC ; 
 qad <= ird ; 
 SLA <=  SLA & TEC  |  ICM & TFC  |  IGM & TGC  ; 
 SLB <=  SLB & TEC  |  ICN & TFC  |  IGN & TGC  ; 
 alb <=  ulb  |  slb  ; 
 OCM <=  GLA & pcd  |  HLA & PCD  ; 
 OCN <=  GLB & pcd  |  HLB & PCD  ; 
 QBE <=  QBE & jqa  |  QAA & QAA  ; 
 QBF <=  QBF & jqa  |  QAC & QAA  ; 
 ULA <=  igm & THC  |  UKD & TIC  |  IGM & TJC  ; 
 ULB <=  ign & THC  |  ULA & TIC  |  IGN & TJC  ; 
 alc <=  ulc  |  slc  ; 
 QBB <=  qac & QAB & QAA  |  QBB & jqa  ; 
 SLC <=  SLC & TED  |  ICO & TFD  |  IGO & TGD  ; 
 SLD <=  SLD & TED  |  ICP & TFD  |  IGP & TGD  ; 
 ald <=  uld  |  sld  ; 
 BLD <=  ULD  |  SLD  ; 
 OCO <=  GLC & pcd  |  HLC & PCD  ; 
 OCP <=  GLD & pcd  |  HLD & PCD  ; 
 qba <=  QAC  |  QAB  |  qaa  ; 
 qbc <=  qac  |  QAB  |  qaa  ; 
 ULC <=  igo & THD  |  ULB & TID  |  IGO & TJD  ; 
 ULD <=  igp & THD  |  ULC & TID  |  IGP & TJD  ; 
 gea <=  eea  |  tde  ; 
 hea <=  EEA  |  tde  ; 
 geb <=  ceb & eeb  |  CEB & EEB  |  tde  ; 
 heb <=  deb & eeb  |  DEB & EEB  |  tde  ; 
 gmc <=  cmc & emc  |  CMC & EMC  |  tdm  ; 
 hmc <=  dmc & emc  |  DMC & EMC  |  tdm  ; 
 gec <=  cec & eec  |  CEC & EEC  |  tde  ; 
 hec <=  dec & eec  |  DEC & EEC  |  tde  ; 
 BEC <=  UEC & TAE  |  WEC  |  WMC & tae  ; 
 ged <=  ced & eed  |  CED & EED  |  tde  ; 
 hed <=  ded & eed  |  DED & EED  |  tde  ; 
 gma <=  ema  |  tdm  ; 
 hma <=  EMA  |  tdm  ; 
 gmb <=  cmb & emb  |  CMB & EMB  |  tdm  ; 
 hmb <=  dmb & emb  |  DMB & EMB  |  tdm  ; 
 hmd <=  dmd & emd  |  DMD & EMD  |  tdm  ; 
 gmd <=  cmd & emd  |  CMD & EMD  |  tdm  ; 
 TDE <= qef ; 
 TAE <= QCF ; 
 BEB <=  UEB & TAE  |  WEB  |  WMB & tae  ; 
 BEF <=  UEB & TAE  |  WEB  |  WMB & tae  ; 
 BEG <=  UEC & TAE  |  WEC  |  WMC & tae  ; 
 KBD <=  CEE & FAF & FAG & FAH  |  CFE & FAG & FAH  |  CGE & FAH  |  CHE  ; 
 BMB <=  UMB  |  SMB  ; 
 BMF <=  UMB  |  SMB  ; 
 BMC <=  UMC  |  SMC  ; 
 BMG <=  UMC  |  SMC  ; 
 TDM <= qde ; 
 aea <=  uea & TAE  |  wea  |  wma & tae  ; 
 BEA <=  UEA & TAE  |  WEA  |  WMA & tae  ; 
 XEA <= TKA & WEA ; 
 XEB <= TKA & WEB ; 
 XMA <= TKA & WMA ; 
 XMB <= TKA & WMB ; 
 SEA <=  SEA & TEA  |  IBA & TFA  |  IFA & TGA  ; 
 SEB <=  SEB & TEA  |  IBB & TFA  |  IFB & TGA  ; 
 aeb <=  ueb & TAE  |  web  |  wmb & tae  ; 
 aec <=  uec & TAE  |  wec  |  wmc & tae  ; 
 OBA <=  GEA & pba  |  HEA & PBA  ; 
 OBB <=  GEB & pba  |  HEB & PBA  ; 
 UEA <=  ifa & THA  |  UDD & TIA  |  IFA & TJA  ; 
 UEB <=  ifb & THA  |  UEA & TIA  |  IFB & TJA  ; 
 XEC <= TKB & WEC ; 
 XED <= TKB & WED ; 
 XMC <= TKB & WMC ; 
 XMD <= TKB & WMD ; 
 SEC <=  SEC & TEB  |  IBC & TFB  |  IFC & TGB  ; 
 SED <=  SED & TEB  |  IBD & TFB  |  IFD & TGB  ; 
 aed <=  ued & TAE  |  wed  |  wmd & tae  ; 
 BED <=  UED & TAE  |  WED  |  WMD & tae  ; 
 OBC <=  GEC & pba  |  HEC & PBA  ; 
 OBD <=  GED & pba  |  HED & PBA  ; 
 UEC <=  ifc & THB  |  UEB & TIB  |  IFC & TJB  ; 
 UED <=  ifd & THB  |  UEC & TIB  |  IFD & TJB  ; 
 ama <=  uma  |  sma  ; 
 BMA <=  UMA  |  SMA  ; 
 ONA <= QNC ; 
 QNA <= JQA ; 
 QNB <= QNA ; 
 QNC <= QNB ; 
 SMA <=  SMA & TEC  |  IDA & TFC  |  IHA & TGC  ; 
 SMB <=  SMB & TEC  |  IDB & TFC  |  IHB & TGC  ; 
 amb <=  umb  |  smb  ; 
 ODA <=  GMA & pda  |  HMA & PDA  ; 
 ODB <=  GMB & pda  |  HMB & PDA  ; 
 QJC <=  JAE  |  JAF  |  JAM  |  JAN  ; 
 UMA <=  iha & THC  |  ULD & TIC  |  IHA & TJC  ; 
 UMB <=  ihb & THC  |  UMA & TIC  |  IHB & TJC  ; 
 amc <=  umc  |  smc  ; 
 SMC <=  SMC & TED  |  IDC & TFD  |  IHC & TGD  ; 
 SMD <=  SMD & TED  |  IDD & TFD  |  IHD & TGD  ; 
 amd <=  umd  |  smd  ; 
 BMD <=  UMD  |  SMD  ; 
 ODC <=  GMC & pda  |  HMC & PDA  ; 
 ODD <=  GMD & pda  |  HMD & PDA  ; 
 UMC <=  ihc & THD  |  UMB & TID  |  IHC & TJD  ; 
 UMD <=  ihd & THD  |  UMC & TID  |  IHD & TJD  ; 
 gfa <=  efa  |  tdf  ; 
 hfa <=  EFA  |  tdf  ; 
 gfb <=  cfb & efb  |  CFB & EFB  |  tdf  ; 
 hfb <=  dfb & efb  |  DFB & EFB  |  tdf  ; 
 dfb <=  bfa  ; 
 hnc <=  dnc & enc  |  DNC & ENC  |  tdn  ; 
 gfc <=  cfc & efc  |  CFC & EFC  |  tdf  ; 
 hfc <=  dfc & efc  |  DFC & EFC  |  tdf  ; 
 gfd <=  cfd & efd  |  CFD & EFD  |  tdf  ; 
 hfd <=  dfd & efd  |  DFD & EFD  |  tdf  ; 
 gna <=  ena  |  tdn  ; 
 hna <=  ENA  |  tdn  ; 
 gnb <=  cnb & enb  |  CNB & ENB  |  tdn  ; 
 hnb <=  dnb & enb  |  DNB & ENB  |  tdn  ; 
 gnc <=  cnc & enc  |  CNC & ENC  |  tdn  ; 
 gnd <=  cnd & endd  |  CND & ENDD   |  tdn  ; 
 hnd <=  dnd & endd  |  DND & ENDD   |  tdn  ; 
 TDF <= qef ; 
 QEE <= QED ; 
 QEF <= QEE ; 
 TAF <= QCF ; 
 mba <=  cee  ; 
 BFB <=  UFB & TAF  |  WFB  |  WNB & taf  ; 
 BFF <=  UFB & TAF  |  WFB  |  WNB & taf  ; 
 BFC <=  UFC & TAF  |  WFC  |  WNC & taf  ; 
 BFG <=  UFC & TAF  |  WFC  |  WNC & taf  ; 
 nba <=  fae  ; 
 nda <=  fam  ; 
 KCD <=  CIE & FAJ & FAK & FAL  |  CJE & FAK & FAL  |  CKE & FAL  |  CLE  ; 
 BNF <=  UNB  |  SNB  ; 
 BNB <=  UNB  |  SNB  ; 
 BNC <=  UNC  |  SNC  ; 
 BNG <=  UNC  |  SNC  ; 
 TDN <= qde ; 
 afa <=  ufa & TAF  |  wfa  |  wna & taf  ; 
 BFA <=  UFA & TAF  |  WFA  |  WNA & taf  ; 
 XFA <= TKA & WFA ; 
 XFB <= TKA & WFB ; 
 XNA <= TKA & WNA ; 
 XNB <= TKA & WNB ; 
 SFA <=  SFA & TEA  |  IBE & TFA  |  IFE & TGA  ; 
 SFB <=  SFB & TEA  |  IBF & TFA  |  IFFF  & TGA  ; 
 afb <=  ufb & TAF  |  wfb  |  wnb & taf  ; 
 OBE <=  GFA & pbb  |  HFA & PBB  ; 
 OBF <=  GFB & pbb  |  HFB & PBB  ; 
 UFA <=  ife & THA  |  UED & TIA  |  IFE & TJA  ; 
 UFB <=  ifff  & THA  |  UFA & TIA  |  IFFF  & TJA  ; 
 afc <=  ufc & TAF  |  wfc  |  wnc & taf  ; 
 XFC <= TKB & WFC ; 
 XFD <= TKB & WFD ; 
 XNC <= TKB & WNC ; 
 XND <= TKB & WND ; 
 SFC <=  SFC & TEB  |  IBG & TFB  |  IFG & TGB  ; 
 SFD <=  SFD & TEB  |  IBH & TFB  |  IFH & TGB  ; 
 afd <=  ufd & TAF  |  wfd  |  wnd & taf  ; 
 BFD <=  UFD & TAF  |  WFD  |  WND & taf  ; 
 OBG <=  GFC & pbb  |  HFC & PBB  ; 
 OBH <=  GFD & pbb  |  HFD & PBB  ; 
 UFC <=  ifg & THB  |  UFB & TIB  |  IFG & TJB  ; 
 UFD <=  ifh & THB  |  UFC & TIB  |  IFH & TJB  ; 
 ana <=  una  |  sna  ; 
 BNA <=  UNA  |  SNA  ; 
 tha <= qfa ; 
 thb <= qfa ; 
 thc <= qfa ; 
 thd <= qfa ; 
 SNA <=  SNA & TEC  |  IDE & TFC  |  IHE & TGC  ; 
 SNB <=  SNB & TEC  |  IDF & TFC  |  IHF & TGC  ; 
 anb <=  unb  |  snb  ; 
 ODE <=  GNA & pdb  |  HNA & PDB  ; 
 ODF <=  GNB & pdb  |  HNB & PDB  ; 
 oea <=  JBA  |  qga  ; 
 UNA <=  ihe & THC  |  UMD & TIC  |  IHE & TJC  ; 
 UNB <=  ihf & THC  |  UNA & TIC  |  IHF & TJC  ; 
 anc <=  unc  |  snc  ; 
 qga <=  jba & qed  |  qga & qed  ; 
 qgb <=  jbb & qed  |  qgb & qed  ; 
 SNC <=  SNC & TED  |  IDG & TFD  |  IHG & TGD  ; 
 SND <=  SND & TED  |  IDH & TFD  |  IHH & TGD  ; 
 andd  <=  und  |  snd  ; 
 BND <=  UND  |  SND  ; 
 ODG <=  GNC & pdb  |  HNC & PDB  ; 
 ODH <=  GND & pdb  |  HND & PDB  ; 
 qea <= qad ; 
 QEB <= QEA ; 
 QEC <= QEB ; 
 QED <= QEC ; 
 UNC <=  ihg & THD  |  UNB & TID  |  IHG & TJD  ; 
 UND <=  ihh & THD  |  UNC & TID  |  IHH & TJD  ; 
 gga <=  ega  |  tdg  ; 
 hga <=  EGA  |  tdg  ; 
 ggb <=  cgb & egb  |  CGB & EGB  |  tdg  ; 
 hgb <=  dgb & egb  |  DGB & EGB  |  tdg  ; 
 hoc <=  doc & eoc  |  DOC & EOC  |  tdo  ; 
 ggc <=  cgc & egc  |  CGC & EGC  |  tdg  ; 
 hgc <=  dgc & egc  |  DGC & EGC  |  tdg  ; 
 hob <=  dob & eob  |  DOB & EOB  |  tdo  ; 
 ggd <=  cgd & egd  |  CGD & EGD  |  tdg  ; 
 hgd <=  dgd & egd  |  DGD & EGD  |  tdg  ; 
 goa <=  eoa  |  tdo  ; 
 hoa <=  EOA  |  tdo  ; 
 gob <=  cob & eob  |  COB & EOB  |  tdo  ; 
 goc <=  coc & eoc  |  COC & EOC  |  tdo  ; 
 god <=  cod & eod  |  COD & EOD  |  tdo  ; 
 hod <=  dod & eod  |  DOD & EOD  |  tdo  ; 
 TDG <= qef ; 
 QCF <= QCE ; 
 TAG <= QCF ; 
 mbb <=  cee & cfe & cfe  |  fbf & cfe  ; 
 BGB <=  UGB & TAG  |  WGB  |  WOB & tag  ; 
 BGF <=  UGB & TAG  |  WGB  |  WOB & tag  ; 
 BGC <=  UGC & TAG  |  WGC  |  WOC & tag  ; 
 BGG <=  UGC & TAG  |  WGC  |  WOC & tag  ; 
 nbb <=  fae  |  faf  ; 
 ndb <=  fam  |  fan  ; 
 lcd <=  fai  |  faj  |  fak  |  fal  ; 
 BOB <=  UOB  |  SOB  ; 
 BOF <=  UOB  |  SOB  ; 
 BOC <=  UOC  |  SOC  ; 
 BOG <=  UOC  |  SOC  ; 
 TDO <= qde ; 
 aka <=  uka  |  ska  ; 
 mdb <=  cme & cne & cne  |  fbn & cne  ; 
 aga <=  uga & TAG  |  wga  |  woa & tag  ; 
 BGA <=  UGA & TAG  |  WGA  |  WOA & tag  ; 
 XGA <= TKA & WGA ; 
 XGB <= TKA & WGB ; 
 XOA <= TKA & WOA ; 
 XOB <= TKA & WOB ; 
 SGA <=  SGA & TEA  |  IBI & TFA  |  IFI & TGA  ; 
 SGB <=  SGB & TEA  |  IBJ & TFA  |  IFJ & TGA  ; 
 agb <=  ugb & TAG  |  wgb  |  wob & tag  ; 
 OBI <=  GGA & pbc  |  HGA & PBC  ; 
 OBJ <=  GGB & pbc  |  HGB & PBC  ; 
 UGA <=  ifi & THA  |  UFD & TIA  |  IFI & TJA  ; 
 UGB <=  ifj & THA  |  UGA & TIA  |  IFJ & TJA  ; 
 agc <=  ugc & TAG  |  wgc  |  woc & tag  ; 
 XGC <= TKB & WGC ; 
 XGD <= TKB & WGD ; 
 XOC <= TKB & WOC ; 
 XOD <= TKB & WOD ; 
 SGC <=  SGC & TEB  |  IBK & TFB  |  IFK & TGB  ; 
 SGD <=  SGD & TEB  |  IBL & TFB  |  IFL & TGB  ; 
 agd <=  ugd & TAG  |  wgd  |  wod & tag  ; 
 BGD <=  UGD & TAG  |  WGD  |  WOD & tag  ; 
 OBK <=  GGC & pbc  |  HGC & PBC  ; 
 OBL <=  GGD & pbc  |  HGD & PBC  ; 
 UGC <=  ifk & THB  |  UGB & TIB  |  IFK & TJB  ; 
 UGD <=  ifl & THB  |  UGC & TIB  |  IFL & TJB  ; 
 aoa <=  uoa  |  soa  ; 
 BOA <=  UOA  |  SOA  ; 
 TIA <= qcg & qfa ; 
 TIB <= qcg & qfa ; 
 TIC <= qcg & qfa ; 
 TID <= qcg & qfa ; 
 SOA <=  SOA & TEC  |  IDI & TFC  |  IHI & TGC  ; 
 SOB <=  SOB & TEC  |  IDJ & TFC  |  IHJ & TGC  ; 
 aob <=  uob  |  sob  ; 
 ODI <=  GOA & pdc  |  HOA & PDC  ; 
 ODJ <=  GOB & pdc  |  HOB & PDC  ; 
 QJD <=  JAG  |  JAH  ; 
 UOA <=  ihi & THC  |  UND & TIC  |  IHI & TJC  ; 
 UOB <=  ihj & THC  |  UOA & TIC  |  IHJ & TJC  ; 
 aoc <=  uoc  |  soc  ; 
 QCG <=  JDA  |  QEA  ; 
 QCE <= QBE ; 
 QFA <= QBF ; 
 QFB <= QFA ; 
 SOC <=  SOC & TED  |  IDK & TFD  |  IHK & TGD  ; 
 SOD <=  SOD & TED  |  IDL & TFD  |  IHL & TGD  ; 
 aod <=  uod  |  sod  ; 
 BOD <=  UOD  |  SOD  ; 
 ODK <=  GOC & pdc  |  HOC & PDC  ; 
 ODL <=  GOD & pdc  |  HOD & PDC  ; 
 QJE <=  JAO  |  JAP  ; 
 UOC <=  ihk & THD  |  UOB & TID  |  IHK & TJD  ; 
 UOD <=  ihl & THD  |  UOC & TID  |  IHL & TJD  ; 
 gha <=  eha  |  tdh  ; 
 hha <=  EHA  |  tdh  ; 
 ghb <=  chb & ehb  |  CHB & EHB  |  tdh  ; 
 hhb <=  dhb & ehb  |  DHB & EHB  |  tdh  ; 
 hpc <=  dpc & epc  |  DPC & EPC  |  tdp  ; 
 ghc <=  chc & ehc  |  CHC & EHC  |  tdh  ; 
 hhc <=  dhc & ehc  |  DHC & EHC  |  tdh  ; 
 hpb <=  dpb & epb  |  DPB & EPB  |  tdp  ; 
 ghd <=  chd & ehd  |  CHD & EHD  |  tdh  ; 
 hhd <=  dhd & ehd  |  DHD & EHD  |  tdh  ; 
 gpa <=  epa  |  tdp  ; 
 hpa <=  EPA  |  tdp  ; 
 gpb <=  cpb & epb  |  CPB & EPB  |  tdp  ; 
 gpc <=  cpc & epc  |  CPC & EPC  |  tdp  ; 
 gpd <=  cpd & epd  |  CPD & EPD  |  tdp  ; 
 hpd <=  dpd & epd  |  DPD & EPD  |  tdp  ; 
 TDH <= qef ; 
 TAH <= QCF ; 
 mbc <=  ZZI & cee & cfe & cge  |  ZZI & cee & cfe & cge  |  fbf & cfe & cge  |  ZZI & fbg & cge  ; 
 BHB <=  UHB & TAH  |  WHB  |  WPB & tah  ; 
 BHF <=  UHB & TAH  |  WHB  |  WPB & tah  ; 
 BHC <=  UHC & TAH  |  WHC  |  WPC & tah  ; 
 BHG <=  UHC & TAH  |  WHC  |  WPC & tah  ; 
 nbc <=  fae  |  faf  |  fag  ; 
 ndc <=  fam  |  fan  |  fao  ; 
 lbc <=  fae  |  faf  |  fag  |  fah  ; 
 lbd <=  fae  |  faf  |  fag  |  fah  ; 
 TDP <= qde ; 
 mdc <=  ZZI & cme & cne & coe  |  ZZI & cme & cne & coe  |  fbn & cne & coe  |  ZZI & fbo & coe  ; 
 aha <=  uha & TAH  |  wha  |  wpa & tah  ; 
 BHA <=  UHA & TAH  |  WHA  |  WPA & tah  ; 
 XHA <= TKA & WHA ; 
 XHB <= TKA & WHB ; 
 XPA <= TKA & WPA ; 
 XPB <= TKA & WPB ; 
 SHA <=  SHA & TEA  |  IBM & TFA  |  IFM & TGA  ; 
 SHB <=  SHB & TEA  |  IBN & TFA  |  IFN & TGA  ; 
 ahb <=  uhb & TAH  |  whb  |  wpb & tah  ; 
 OBM <=  GHA & pbd  |  HHA & PBD  ; 
 OBN <=  GHB & pbd  |  HHB & PBD  ; 
 UHA <=  ifm & THA  |  UGD & TIA  |  IFM & TJA  ; 
 UHB <=  ifn & THA  |  UHA & TIA  |  IFN & TJA  ; 
 ahc <=  uhc & TAH  |  whc  |  wpc & tah  ; 
 XHC <= TKB & WHC ; 
 XHD <= TKB & WHD ; 
 XPC <= TKB & WPC ; 
 XPD <= TKB & WPD ; 
 SHC <=  SHC & TEB  |  IBO & TFB  |  IFO & TGB  ; 
 SHD <=  SHD & TEB  |  IBP & TFB  |  IFP & TGB  ; 
 ahd <=  uhd & TAH  |  whd  |  wpd & tah  ; 
 BHD <=  UHD & TAH  |  WHD  |  WPD & tah  ; 
 OBO <=  GHC & pbd  |  HHC & PBD  ; 
 OBP <=  GHD & pbd  |  HHD & PBD  ; 
 UHC <=  ifo & THB  |  UHB & TIB  |  IFO & TJB  ; 
 UHD <=  ifp & THB  |  UHC & TIB  |  IFP & TJB  ; 
 apa <=  upa  |  spa  ; 
 BPA <=  UPA  |  SPA  ; 
 tja <= qcg ; 
 tjb <= qcg ; 
 tjc <= qcg ; 
 tjd <= qcg ; 
 SPA <=  SPA & TEC  |  IDM & TFC  |  IHM & TGC  ; 
 SPB <=  SPB & TEC  |  IDN & TFC  |  IHN & TGC  ; 
 apb <=  upb  |  spb  ; 
 BPB <=  UPB  |  SPB  ; 
 ODM <=  GPA & pdd  |  HPA & PDD  ; 
 ODN <=  GPB & pdd  |  HPB & PDD  ; 
 OEB <= QHA ; 
 OEC <= QHA ; 
 UPA <=  ihm & THC  |  UOD & TIC  |  IHM & TJC  ; 
 UPB <=  ihn & THC  |  UPA & TIC  |  IHN & TJC  ; 
 apc <=  upc  |  spc  ; 
 BPC <=  UPC  |  SPC  ; 
 OFA <= QGB & UPE ; 
 OFB <= QGB & UPE ; 
 SPC <=  SPC & TED  |  IDO & TFD  |  IHO & TGD  ; 
 SPD <=  SPD & TED  |  IDP & TFD  |  IHP & TGD  ; 
 apd <=  upd  |  spd  ; 
 BPD <=  UPD  |  SPD  ; 
 ODO <=  GPC & pdd  |  HPC & PDD  ; 
 ODP <=  GPD & pdd  |  HPD & PDD  ; 
 QHA <= QGB & jbb ; 
 UPE <= QGB & UPD ; 
 UPC <=  iho & THD  |  UPB & TID  |  IHO & TJD  ; 
 UPD <=  ihp & THD  |  UPC & TID  |  IHP & TJD  ; 
end 
endmodule;
