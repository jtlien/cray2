module mif( IZZ,
 IAA, 
 IAB, 
 IAC, 
 IAD, 
 IAE, 
 IAF, 
 IAG, 
 IAH, 
 IAI, 
 IAJ, 
 IAK, 
 IAL, 
 IAM, 
 IAN, 
 IAO, 
 IAP, 
 IBA, 
 IBB, 
 IBC, 
 IBD, 
 IBE, 
 IBF, 
 IBG, 
 IBH, 
 IBI, 
 IBJ, 
 IBK, 
 IBL, 
 IBM, 
 IBN, 
 IBO, 
 IBP, 
 ICA, 
 ICB, 
 ICC, 
 ICD, 
 ICE, 
 ICF, 
 ICG, 
 ICH, 
 ICI, 
 ICJ, 
 ICK, 
 ICL, 
 ICM, 
 ICN, 
 ICO, 
 ICP, 
 IDA, 
 IDB, 
 IDC, 
 IDD, 
 IDE, 
 IDF, 
 IDG, 
 IDH, 
 IDI, 
 IDJ, 
 IDK, 
 IDL, 
 IDM, 
 IDN, 
 IDO, 
 IDP, 
 IEA, 
 IEB, 
 IEC, 
 IED, 
 IEE, 
 IEF, 
 IEG, 
 IEH, 
 IEI, 
 IEJ, 
 IEK, 
 IEL, 
 IEM, 
 IEN, 
 IEO, 
 IEP, 
 IFA, 
 IFB, 
 IFC, 
 IFD, 
 IFE, 
 IFFF , 
 IFG, 
 IFH, 
 IFI, 
 IGA, 
 IGB, 
 IGC, 
 IHB, 
 IHC, 
 IJA, 
 IJB, 
 IJC, 
 IJD, 
 IKA, 
 IKB, 
 ILA, 
 ILB, 
 ILC, 
 IMA, 
 IMB, 
 IMC, 
 IMD, 
 IME, 
 IMF, 
 IMG, 
 INA, 
 IOA, 
 IOB, 
 IOC, 
 IOD, 
 IPA, 
 IPB, 
 IPC, 
 IPD, 
 IPE, 
 IPF, 
 IQA, 
 IQB, 
 IQC, 
 IQD, 
 IQE, 
 IQF, 
 IQG, 
 IQH, 
 IQI, 
 OAA, 
 OAB, 
 OAC, 
 OAD, 
 OAE, 
 OAF, 
 OAG, 
 OAH, 
 OAI, 
 OAJ, 
 OAK, 
 OAL, 
 OAM, 
 OAN, 
 OAO, 
 OAP, 
 OBA, 
 OBB, 
 OBC, 
 OBD, 
 OBE, 
 OBF, 
 OBG, 
 OBH, 
 OBI, 
 OBJ, 
 OBK, 
 OBL, 
 OBM, 
 OBN, 
 OBO, 
 OBP, 
 OCA, 
 OCB, 
 OCC, 
 OCD, 
 OCE, 
 OCF, 
 OCG, 
 OCH, 
 OCI, 
 OCJ, 
 OCK, 
 OCL, 
 OCM, 
 OCN, 
 OCO, 
 OCP, 
 ODA, 
 ODB, 
 ODC, 
 ODD, 
 ODE, 
 ODF, 
 ODG, 
 ODH, 
 ODI, 
 ODJ, 
 ODK, 
 ODL, 
 ODM, 
 ODN, 
 ODO, 
 ODP, 
 OEA, 
 OEB, 
 OEC, 
 OED, 
 OEE, 
 OEF, 
 OEG, 
 OEH, 
 OEI, 
 OEJ, 
 OEK, 
 OEL, 
 OEM, 
 OEN, 
 OEO, 
 OEP, 
 OEQ, 
 OER, 
 OES, 
 OET, 
 OEU, 
 OEV, 
 OEW, 
 OEX, 
 OEY, 
 OFA, 
 OFB, 
 OFC, 
 OGA, 
 OGB, 
 OGC, 
 OGD, 
 OGE, 
 OGF, 
 OGG, 
 OGH, 
 OGI, 
 OGJ, 
 OHA, 
 OHB, 
 OHC, 
 OHD, 
 OHE, 
 OIA, 
 OIB, 
 OIC, 
 OID, 
 OIE, 
 OIG, 
 OJA, 
 OJB, 
 OJC, 
 OJD, 
 OJE, 
 OKA, 
 OKB, 
 OLA, 
 OLB, 
 OLC, 
 OLD, 
 OLF, 
 OMA, 
 OMB, 
 OQA, 
 OQB, 
 ORA, 
 ORB, 
 ORC, 
 ORD, 
 ORE, 
 ORF, 
 OTA, 
 OTB, 
 OTC, 
 OTD, 
 OTE, 
OTF ); 
    
 input IZZ; 
 input IAA; 
 input IAB; 
 input IAC; 
 input IAD; 
 input IAE; 
 input IAF; 
 input IAG; 
 input IAH; 
 input IAI; 
 input IAJ; 
 input IAK; 
 input IAL; 
 input IAM; 
 input IAN; 
 input IAO; 
 input IAP; 
 input IBA; 
 input IBB; 
 input IBC; 
 input IBD; 
 input IBE; 
 input IBF; 
 input IBG; 
 input IBH; 
 input IBI; 
 input IBJ; 
 input IBK; 
 input IBL; 
 input IBM; 
 input IBN; 
 input IBO; 
 input IBP; 
 input ICA; 
 input ICB; 
 input ICC; 
 input ICD; 
 input ICE; 
 input ICF; 
 input ICG; 
 input ICH; 
 input ICI; 
 input ICJ; 
 input ICK; 
 input ICL; 
 input ICM; 
 input ICN; 
 input ICO; 
 input ICP; 
 input IDA; 
 input IDB; 
 input IDC; 
 input IDD; 
 input IDE; 
 input IDF; 
 input IDG; 
 input IDH; 
 input IDI; 
 input IDJ; 
 input IDK; 
 input IDL; 
 input IDM; 
 input IDN; 
 input IDO; 
 input IDP; 
 input IEA; 
 input IEB; 
 input IEC; 
 input IED; 
 input IEE; 
 input IEF; 
 input IEG; 
 input IEH; 
 input IEI; 
 input IEJ; 
 input IEK; 
 input IEL; 
 input IEM; 
 input IEN; 
 input IEO; 
 input IEP; 
 input IFA; 
 input IFB; 
 input IFC; 
 input IFD; 
 input IFE; 
 input IFFF ; 
 input IFG; 
 input IFH; 
 input IFI; 
 input IGA; 
 input IGB; 
 input IGC; 
 input IHB; 
 input IHC; 
 input IJA; 
 input IJB; 
 input IJC; 
 input IJD; 
 input IKA; 
 input IKB; 
 input ILA; 
 input ILB; 
 input ILC; 
 input IMA; 
 input IMB; 
 input IMC; 
 input IMD; 
 input IME; 
 input IMF; 
 input IMG; 
 input INA; 
 input IOA; 
 input IOB; 
 input IOC; 
 input IOD; 
 input IPA; 
 input IPB; 
 input IPC; 
 input IPD; 
 input IPE; 
 input IPF; 
 input IQA; 
 input IQB; 
 input IQC; 
 input IQD; 
 input IQE; 
 input IQF; 
 input IQG; 
 input IQH; 
 input IQI; 

 output OAA; 
 output OAB; 
 output OAC; 
 output OAD; 
 output OAE; 
 output OAF; 
 output OAG; 
 output OAH; 
 output OAI; 
 output OAJ; 
 output OAK; 
 output OAL; 
 output OAM; 
 output OAN; 
 output OAO; 
 output OAP; 
 output OBA; 
 output OBB; 
 output OBC; 
 output OBD; 
 output OBE; 
 output OBF; 
 output OBG; 
 output OBH; 
 output OBI; 
 output OBJ; 
 output OBK; 
 output OBL; 
 output OBM; 
 output OBN; 
 output OBO; 
 output OBP; 
 output OCA; 
 output OCB; 
 output OCC; 
 output OCD; 
 output OCE; 
 output OCF; 
 output OCG; 
 output OCH; 
 output OCI; 
 output OCJ; 
 output OCK; 
 output OCL; 
 output OCM; 
 output OCN; 
 output OCO; 
 output OCP; 
 output ODA; 
 output ODB; 
 output ODC; 
 output ODD; 
 output ODE; 
 output ODF; 
 output ODG; 
 output ODH; 
 output ODI; 
 output ODJ; 
 output ODK; 
 output ODL; 
 output ODM; 
 output ODN; 
 output ODO; 
 output ODP; 
 output OEA; 
 output OEB; 
 output OEC; 
 output OED; 
 output OEE; 
 output OEF; 
 output OEG; 
 output OEH; 
 output OEI; 
 output OEJ; 
 output OEK; 
 output OEL; 
 output OEM; 
 output OEN; 
 output OEO; 
 output OEP; 
 output OEQ; 
 output OER; 
 output OES; 
 output OET; 
 output OEU; 
 output OEV; 
 output OEW; 
 output OEX; 
 output OEY; 
 output OFA; 
 output OFB; 
 output OFC; 
 output OGA; 
 output OGB; 
 output OGC; 
 output OGD; 
 output OGE; 
 output OGF; 
 output OGG; 
 output OGH; 
 output OGI; 
 output OGJ; 
 output OHA; 
 output OHB; 
 output OHC; 
 output OHD; 
 output OHE; 
 output OIA; 
 output OIB; 
 output OIC; 
 output OID; 
 output OIE; 
 output OIG; 
 output OJA; 
 output OJB; 
 output OJC; 
 output OJD; 
 output OJE; 
 output OKA; 
 output OKB; 
 output OLA; 
 output OLB; 
 output OLC; 
 output OLD; 
 output OLF; 
 output OMA; 
 output OMB; 
 output OQA; 
 output OQB; 
 output ORA; 
 output ORB; 
 output ORC; 
 output ORD; 
 output ORE; 
 output ORF; 
 output OTA; 
 output OTB; 
 output OTC; 
 output OTD; 
 output OTE; 
 output OTF; 
  
  
reg  AAA ;
reg  AAB ;
reg  AAC ;
reg  AAD ;
reg  AAE ;
reg  AAF ;
reg  AAG ;
reg  AAH ;
reg  AAI ;
reg  AAJ ;
reg  AAK ;
reg  AAL ;
reg  AAM ;
reg  AAN ;
reg  AAO ;
reg  AAP ;
reg  ABA ;
reg  ABB ;
reg  ABC ;
reg  ABD ;
reg  ABE ;
reg  ABF ;
reg  ABG ;
reg  ABH ;
reg  ABI ;
reg  ABJ ;
reg  ABK ;
reg  ABL ;
reg  ABM ;
reg  ABN ;
reg  ABO ;
reg  ABP ;
reg  ach ;
reg  aci ;
reg  acj ;
reg  ack ;
reg  acl ;
reg  acm ;
reg  acn ;
reg  aco ;
reg  acp ;
reg  ada ;
reg  adb ;
reg  adc ;
reg  add ;
reg  ade ;
reg  adf ;
reg  adg ;
reg  adh ;
reg  adi ;
reg  adj ;
reg  adk ;
reg  adl ;
reg  adm ;
reg  adn ;
reg  ado ;
reg  AEH ;
reg  AEI ;
reg  AEJ ;
reg  AEK ;
reg  AEL ;
reg  AEM ;
reg  AEN ;
reg  AEO ;
reg  AEP ;
reg  AFA ;
reg  AFB ;
reg  AFC ;
reg  AFD ;
reg  AFE ;
reg  AFF ;
reg  AFG ;
reg  AFH ;
reg  AFI ;
reg  AFJ ;
reg  AFK ;
reg  AFL ;
reg  AFM ;
reg  AFN ;
reg  AFO ;
reg  AGH ;
reg  AGI ;
reg  AGJ ;
reg  AGK ;
reg  AGL ;
reg  AGM ;
reg  AGN ;
reg  AGO ;
reg  AGP ;
reg  AHA ;
reg  AHB ;
reg  AHC ;
reg  AHD ;
reg  AHE ;
reg  AHF ;
reg  AHG ;
reg  AHH ;
reg  AHI ;
reg  AHJ ;
reg  AHK ;
reg  AHL ;
reg  AHM ;
reg  AHN ;
reg  AHO ;
reg  AIH ;
reg  AII ;
reg  AIJ ;
reg  AIK ;
reg  AIL ;
reg  AIM ;
reg  AIN ;
reg  AIO ;
reg  AIP ;
reg  AJA ;
reg  AJB ;
reg  AJC ;
reg  AJD ;
reg  AJE ;
reg  AJF ;
reg  AJG ;
reg  AJH ;
reg  AJI ;
reg  AJJ ;
reg  AJK ;
reg  AJL ;
reg  AJM ;
reg  AJN ;
reg  AJO ;
reg  AKH ;
reg  AKI ;
reg  AKJ ;
reg  AKK ;
reg  AKL ;
reg  AKM ;
reg  AKN ;
reg  AKO ;
reg  AKP ;
reg  ALA ;
reg  ALB ;
reg  ALC ;
reg  ALD ;
reg  ALE ;
reg  ALF ;
reg  ALG ;
reg  ALH ;
reg  ALI ;
reg  ALJ ;
reg  ALK ;
reg  ALL ;
reg  ALM ;
reg  ALN ;
reg  ALO ;
reg  AMH ;
reg  AMI ;
reg  AMJ ;
reg  AMK ;
reg  AML ;
reg  AMM ;
reg  AMN ;
reg  AMO ;
reg  AMP ;
reg  ANA ;
reg  ANB ;
reg  ANC ;
reg  ANDD  ;
reg  ANE ;
reg  ANF ;
reg  ANG ;
reg  ANH ;
reg  ANI ;
reg  ANJ ;
reg  ANK ;
reg  ANL ;
reg  ANM ;
reg  ANN ;
reg  ANO ;
reg  AOH ;
reg  AOI ;
reg  AOJ ;
reg  AOK ;
reg  AOL ;
reg  AOM ;
reg  AON ;
reg  AOO ;
reg  AOP ;
reg  APA ;
reg  APB ;
reg  APC ;
reg  APD ;
reg  APE ;
reg  APF ;
reg  APG ;
reg  APH ;
reg  API ;
reg  APJ ;
reg  APK ;
reg  APL ;
reg  APM ;
reg  APN ;
reg  APO ;
reg  AQH ;
reg  AQI ;
reg  AQJ ;
reg  AQK ;
reg  AQL ;
reg  AQM ;
reg  AQN ;
reg  AQO ;
reg  AQP ;
reg  ARA ;
reg  ARB ;
reg  ARC ;
reg  ARD ;
reg  ARE ;
reg  ARF ;
reg  ARG ;
reg  ARH ;
reg  ARI ;
reg  ARJ ;
reg  ARK ;
reg  ARL ;
reg  ARM ;
reg  ARN ;
reg  ARO ;
reg  ASH ;
reg  ASI ;
reg  ASJ ;
reg  ASK ;
reg  ASL ;
reg  ASM ;
reg  ASN ;
reg  ASO ;
reg  ASP ;
reg  ATA ;
reg  ATB ;
reg  ATC ;
reg  ATD ;
reg  ATE ;
reg  ATF ;
reg  ATG ;
reg  ATH ;
reg  ATI ;
reg  ATJ ;
reg  ATK ;
reg  ATL ;
reg  ATM ;
reg  ATN ;
reg  ATO ;
reg  ATP ;
reg  BAH ;
reg  BAI ;
reg  BAJ ;
reg  BAK ;
reg  BAL ;
reg  BAM ;
reg  BAN ;
reg  BAO ;
reg  BAP ;
reg  BBA ;
reg  BBB ;
reg  BBC ;
reg  BBD ;
reg  BBE ;
reg  BBF ;
reg  BBG ;
reg  BBH ;
reg  BBI ;
reg  BBJ ;
reg  BBK ;
reg  BBL ;
reg  BBM ;
reg  BBN ;
reg  BBO ;
reg  BBP ;
reg  BCI ;
reg  BCJ ;
reg  BCK ;
reg  BCM ;
reg  BCN ;
reg  BCO ;
reg  BDA ;
reg  BDB ;
reg  BDC ;
reg  BDE ;
reg  BDF ;
reg  BDG ;
reg  BDI ;
reg  BDJ ;
reg  BDK ;
reg  BDM ;
reg  BDN ;
reg  BDO ;
reg  BEH ;
reg  BEI ;
reg  BEJ ;
reg  BEK ;
reg  BEL ;
reg  BEM ;
reg  BEN ;
reg  BEO ;
reg  BEP ;
reg  BFA ;
reg  BFB ;
reg  BFC ;
reg  BFD ;
reg  BFE ;
reg  BFF ;
reg  BFG ;
reg  BFH ;
reg  BFI ;
reg  BFJ ;
reg  BFK ;
reg  BFL ;
reg  CAA ;
reg  CAB ;
reg  CAC ;
reg  CCA ;
reg  CCB ;
reg  CDA ;
reg  CDB ;
reg  CEA ;
reg  CEB ;
reg  CFA ;
reg  CFB ;
reg  CGA ;
reg  CGB ;
reg  CHA ;
reg  CHB ;
reg  CIA ;
reg  CIB ;
reg  CJA ;
reg  CJB ;
reg  DAA ;
reg  DAB ;
reg  DAC ;
reg  DAD ;
reg  DAE ;
reg  DAF ;
reg  DAG ;
reg  DAH ;
reg  DAI ;
reg  DAJ ;
reg  DAK ;
reg  DAL ;
reg  DAM ;
reg  DAN ;
reg  DAO ;
reg  DAP ;
reg  DBA ;
reg  DBB ;
reg  DBC ;
reg  DBD ;
reg  DBE ;
reg  DBF ;
reg  DBG ;
reg  DBH ;
reg  DBI ;
reg  DBJ ;
reg  DBK ;
reg  DBL ;
reg  DBM ;
reg  DBN ;
reg  DBO ;
reg  DBP ;
reg  eaa ;
reg  eab ;
reg  eac ;
reg  ead ;
reg  eae ;
reg  eaf ;
reg  eag ;
reg  eah ;
reg  eai ;
reg  eaj ;
reg  eak ;
reg  eal ;
reg  eam ;
reg  ean ;
reg  eao ;
reg  eap ;
reg  ebj ;
reg  ebk ;
reg  ebl ;
reg  ebp ;
reg  eci ;
reg  ecj ;
reg  eck ;
reg  ecl ;
reg  ecm ;
reg  ecn ;
reg  eco ;
reg  EDA ;
reg  EDB ;
reg  EDC ;
reg  EDD ;
reg  EDE ;
reg  EDF ;
reg  EDG ;
reg  EDH ;
reg  EDI ;
reg  EDJ ;
reg  EDK ;
reg  EDL ;
reg  EDM ;
reg  EDN ;
reg  EDO ;
reg  EDP ;
reg  gaa ;
reg  gab ;
reg  gac ;
reg  GAE ;
reg  gaf ;
reg  gag ;
reg  gah ;
reg  gai ;
reg  gal ;
reg  gam ;
reg  gan ;
reg  gao ;
reg  gap ;
reg  gba ;
reg  gbc ;
reg  gbd ;
reg  gbe ;
reg  gbf ;
reg  gbg ;
reg  gbh ;
reg  gbi ;
reg  gbj ;
reg  gbk ;
reg  gbm ;
reg  gbn ;
reg  gbo ;
reg  gbp ;
reg  gca ;
reg  gcb ;
reg  gcc ;
reg  gcd ;
reg  gch ;
reg  gci ;
reg  gcj ;
reg  gck ;
reg  gcl ;
reg  gcm ;
reg  gcn ;
reg  GDA ;
reg  GDB ;
reg  GDC ;
reg  GDD ;
reg  GDE ;
reg  GDF ;
reg  GDG ;
reg  GDH ;
reg  GDI ;
reg  GDJ ;
reg  GDK ;
reg  GDL ;
reg  GDX ;
reg  GDY ;
reg  haa ;
reg  hab ;
reg  hac ;
reg  had ;
reg  HAE ;
reg  HAF ;
reg  HAG ;
reg  HAH ;
reg  hba ;
reg  hbb ;
reg  hbc ;
reg  hbd ;
reg  hbe ;
reg  hbf ;
reg  hbg ;
reg  hbh ;
reg  hca ;
reg  hcb ;
reg  hcc ;
reg  hcd ;
reg  hce ;
reg  hcf ;
reg  hcg ;
reg  hch ;
reg  hda ;
reg  hdb ;
reg  hdc ;
reg  hdd ;
reg  hde ;
reg  hdf ;
reg  hdh ;
reg  HDI ;
reg  HDJ ;
reg  HDK ;
reg  HDL ;
reg  hea ;
reg  heb ;
reg  heh ;
reg  HEI ;
reg  HEJ ;
reg  HEO ;
reg  HEP ;
reg  HFM ;
reg  HFN ;
reg  HIA ;
reg  HIB ;
reg  HIC ;
reg  HJA ;
reg  HJB ;
reg  HJC ;
reg  HKA ;
reg  HKB ;
reg  HKC ;
reg  HLA ;
reg  HLB ;
reg  HLC ;
reg  HMA ;
reg  HMB ;
reg  HMC ;
reg  HNA ;
reg  HNB ;
reg  HNC ;
reg  HOA ;
reg  HOB ;
reg  HOC ;
reg  HPA ;
reg  HPB ;
reg  HPC ;
reg  KAA ;
reg  KAB ;
reg  KAC ;
reg  KAD ;
reg  KAE ;
reg  KAF ;
reg  LAA ;
reg  LAB ;
reg  LAC ;
reg  LAD ;
reg  LAE ;
reg  LAF ;
reg  LBA ;
reg  LBB ;
reg  LBC ;
reg  LBD ;
reg  LBE ;
reg  LBF ;
reg  MAA ;
reg  MAB ;
reg  MAC ;
reg  NAA ;
reg  NAB ;
reg  NAC ;
reg  NAD ;
reg  NAE ;
reg  NBA ;
reg  NBB ;
reg  NBC ;
reg  NBD ;
reg  NCA ;
reg  NCB ;
reg  OAA ;
reg  OAB ;
reg  OAC ;
reg  OAD ;
reg  OAE ;
reg  OAF ;
reg  OAG ;
reg  OAH ;
reg  OAI ;
reg  OAJ ;
reg  OAK ;
reg  OAL ;
reg  OAM ;
reg  OAN ;
reg  OAO ;
reg  OAP ;
reg  OBA ;
reg  OBB ;
reg  OBC ;
reg  OBD ;
reg  OBE ;
reg  OBF ;
reg  OBG ;
reg  OBH ;
reg  OBI ;
reg  OBJ ;
reg  OBK ;
reg  OBL ;
reg  OBM ;
reg  OBN ;
reg  OBO ;
reg  OBP ;
reg  oca ;
reg  ocb ;
reg  occ ;
reg  ocd ;
reg  oce ;
reg  ocf ;
reg  ocg ;
reg  och ;
reg  oci ;
reg  ocj ;
reg  ock ;
reg  ocl ;
reg  ocm ;
reg  ocn ;
reg  oco ;
reg  ocp ;
reg  oda ;
reg  odb ;
reg  odc ;
reg  odd ;
reg  ode ;
reg  odf ;
reg  odg ;
reg  odh ;
reg  odi ;
reg  odj ;
reg  odk ;
reg  odl ;
reg  odm ;
reg  odn ;
reg  odo ;
reg  odp ;
reg  OEA ;
reg  OEB ;
reg  OEC ;
reg  OED ;
reg  OEE ;
reg  OEF ;
reg  OEG ;
reg  OEH ;
reg  oei ;
reg  OEJ ;
reg  OEK ;
reg  OEL ;
reg  OEM ;
reg  OEN ;
reg  OEO ;
reg  OEP ;
reg  oeq ;
reg  oer ;
reg  OES ;
reg  OET ;
reg  OEU ;
reg  OEV ;
reg  OEW ;
reg  OEX ;
reg  OEY ;
reg  OFA ;
reg  ofb ;
reg  OFC ;
reg  OGA ;
reg  OGB ;
reg  OGC ;
reg  OGD ;
reg  OGE ;
reg  OGF ;
reg  OGG ;
reg  OGH ;
reg  OGI ;
reg  OGJ ;
reg  OHA ;
reg  OHB ;
reg  OHC ;
reg  OHD ;
reg  OHE ;
reg  OIA ;
reg  oib ;
reg  OIC ;
reg  OID ;
reg  OIE ;
reg  oig ;
reg  OJA ;
reg  OJB ;
reg  OJC ;
reg  OJD ;
reg  OJE ;
reg  OKA ;
reg  OKB ;
reg  OLA ;
reg  OLB ;
reg  OLC ;
reg  old ;
reg  OLF ;
reg  OMA ;
reg  OMB ;
reg  oqa ;
reg  OQB ;
reg  ora ;
reg  orb ;
reg  orc ;
reg  ord ;
reg  ore ;
reg  orf ;
reg  OTA ;
reg  OTB ;
reg  OTC ;
reg  otd ;
reg  ote ;
reg  otf ;
reg  PAA ;
reg  PAB ;
reg  PAC ;
reg  PAD ;
reg  PAE ;
reg  PAF ;
reg  PAG ;
reg  PAH ;
reg  PAI ;
reg  PAJ ;
reg  PAK ;
reg  PAL ;
reg  PAM ;
reg  PAN ;
reg  PAO ;
reg  PAP ;
reg  PBA ;
reg  PBB ;
reg  PBC ;
reg  PBD ;
reg  PBE ;
reg  PBF ;
reg  PBG ;
reg  PBH ;
reg  PBI ;
reg  PBJ ;
reg  PBK ;
reg  PBL ;
reg  PBM ;
reg  PBN ;
reg  PBO ;
reg  PBP ;
reg  PCA ;
reg  PCB ;
reg  PCC ;
reg  PCD ;
reg  PCE ;
reg  PCF ;
reg  PCG ;
reg  PCH ;
reg  PCI ;
reg  PCJ ;
reg  PCK ;
reg  PCL ;
reg  PCM ;
reg  PCN ;
reg  PCO ;
reg  PCP ;
reg  PDA ;
reg  PDB ;
reg  PDC ;
reg  PDD ;
reg  PDE ;
reg  PDF ;
reg  PDG ;
reg  PDH ;
reg  PDI ;
reg  PDJ ;
reg  PDK ;
reg  PDL ;
reg  PDM ;
reg  PDN ;
reg  PDO ;
reg  PDP ;
reg  PEB ;
reg  PEC ;
reg  PED ;
reg  PEE ;
reg  PEF ;
reg  PEG ;
reg  PEH ;
reg  PEI ;
reg  PEJ ;
reg  PEK ;
reg  PEL ;
reg  PEM ;
reg  PEN ;
reg  PEO ;
reg  PEP ;
reg  PFA ;
reg  PFB ;
reg  PFC ;
reg  PFD ;
reg  PFE ;
reg  PFF ;
reg  PFG ;
reg  PFH ;
reg  PFI ;
reg  PFJ ;
reg  PFK ;
reg  PFL ;
reg  QAA ;
reg  QAB ;
reg  QAC ;
reg  QAD ;
reg  QBA ;
reg  QCD ;
reg  QCH ;
reg  QCI ;
reg  QCJ ;
reg  qck ;
reg  QCX ;
reg  QCY ;
reg  QCZ ;
reg  QEA ;
reg  QEB ;
reg  QFA ;
reg  QFB ;
reg  QFC ;
reg  QGA ;
reg  QGB ;
reg  qgd ;
reg  QGE ;
reg  QHA ;
reg  QHC ;
reg  QHD ;
reg  QHE ;
reg  QHF ;
reg  qia ;
reg  qib ;
reg  qic ;
reg  qid ;
reg  QKA ;
reg  QKB ;
reg  QKC ;
reg  QKD ;
reg  QKE ;
reg  QKF ;
reg  QKG ;
reg  QKH ;
reg  QKJ ;
reg  QKK ;
reg  QKL ;
reg  QKM ;
reg  QKN ;
reg  QKO ;
reg  QKP ;
reg  QKQ ;
reg  QKR ;
reg  QKS ;
reg  QKT ;
reg  QKW ;
reg  QKX ;
reg  QKY ;
reg  QLA ;
reg  QLB ;
reg  QLC ;
reg  QLD ;
reg  QLE ;
reg  QLF ;
reg  QLG ;
reg  QLI ;
reg  QLJ ;
reg  QLK ;
reg  QLL ;
reg  QLM ;
reg  QLN ;
reg  QLO ;
reg  QLP ;
reg  QLQ ;
reg  QLR ;
reg  QLS ;
reg  qlx ;
reg  QMA ;
reg  qmb ;
reg  qmc ;
reg  QME ;
reg  qmf ;
reg  qmg ;
reg  QMI ;
reg  qmj ;
reg  QMK ;
reg  QML ;
reg  qna ;
reg  qnb ;
reg  qnc ;
reg  QND ;
reg  qne ;
reg  qnf ;
reg  qng ;
reg  QNI ;
reg  qnj ;
reg  QNM ;
reg  qnn ;
reg  QNQ ;
reg  qnr ;
reg  QNU ;
reg  qnv ;
reg  qoa ;
reg  QPA ;
reg  QPB ;
reg  QPC ;
reg  QPD ;
reg  QQA ;
reg  QQB ;
reg  QQC ;
reg  QQD ;
reg  QQE ;
reg  QQF ;
reg  QQG ;
reg  QQH ;
reg  QQI ;
reg  QQJ ;
reg  QQK ;
reg  QQL ;
reg  QQM ;
reg  QQN ;
reg  QQO ;
reg  QQP ;
reg  QQQ ;
reg  QQR ;
reg  QQS ;
reg  QQT ;
reg  QQW ;
reg  qqx ;
reg  QQY ;
reg  QQZ ;
reg  QRA ;
reg  QRB ;
reg  QRC ;
reg  QRD ;
reg  QRE ;
reg  QRF ;
reg  QSA ;
reg  QSB ;
reg  QSC ;
reg  QSD ;
reg  QSE ;
reg  QSF ;
reg  QSG ;
reg  QSH ;
reg  qsi ;
reg  QTA ;
reg  qtb ;
reg  QTC ;
reg  QTD ;
reg  QTE ;
reg  QTF ;
reg  QTG ;
reg  QTH ;
reg  QTI ;
reg  QTJ ;
reg  QTM ;
reg  QTN ;
reg  QTO ;
reg  QTP ;
reg  qtq ;
reg  qtr ;
reg  QTW ;
reg  QTX ;
reg  QUA ;
reg  QUB ;
reg  QUC ;
reg  QUD ;
reg  QUE ;
reg  QUF ;
reg  qva ;
reg  qvb ;
reg  qvc ;
reg  qvd ;
reg  qve ;
reg  qvf ;
reg  qvg ;
reg  qvh ;
reg  qvi ;
reg  qvj ;
reg  QWA ;
reg  QWB ;
reg  QWC ;
reg  qwd ;
reg  qwe ;
reg  qwf ;
reg  qwg ;
reg  qwh ;
reg  qwi ;
reg  QWJ ;
reg  QXA ;
reg  QXB ;
reg  QXC ;
reg  QXD ;
reg  QXE ;
reg  QXF ;
reg  QYA ;
reg  QYB ;
reg  QYC ;
reg  QYD ;
reg  qza ;
reg  qzd ;
reg  QZE ;
reg  QZF ;
reg  raa ;
reg  RAB ;
reg  RAC ;
reg  RAD ;
reg  RAE ;
reg  RAF ;
reg  RAG ;
reg  rat ;
reg  RAX ;
reg  rba ;
reg  RBB ;
reg  RBC ;
reg  RBD ;
reg  RBE ;
reg  RBF ;
reg  RBG ;
reg  RBH ;
reg  RBI ;
reg  RBX ;
reg  REC ;
reg  RFA ;
reg  RFB ;
reg  RGA ;
reg  RGB ;
reg  RGC ;
reg  RGD ;
reg  RHA ;
reg  RHB ;
reg  RHC ;
reg  RHD ;
reg  RHE ;
reg  RHF ;
reg  RHG ;
reg  RHH ;
reg  RHI ;
reg  RHJ ;
reg  RIA ;
reg  RIB ;
reg  RIC ;
reg  RID ;
reg  RIE ;
reg  RIF ;
reg  RIX ;
reg  RJA ;
reg  RJB ;
reg  RJC ;
reg  RJD ;
reg  rje ;
reg  RJF ;
reg  RJG ;
reg  RJH ;
reg  RJI ;
reg  RJK ;
reg  RJL ;
reg  RKA ;
reg  RKB ;
reg  RKC ;
reg  RKD ;
reg  RLA ;
reg  RLB ;
reg  RLC ;
reg  RLD ;
reg  RLX ;
reg  RMA ;
reg  RMB ;
reg  RMC ;
reg  RMD ;
reg  RME ;
reg  RMF ;
reg  RMG ;
reg  RMH ;
reg  RMI ;
reg  RMJ ;
reg  RMK ;
reg  RML ;
reg  RMM ;
reg  RMN ;
reg  RMO ;
reg  RMP ;
reg  RMQ ;
reg  RMR ;
reg  RMS ;
reg  RMT ;
reg  RMU ;
reg  rmv ;
reg  RNA ;
reg  RNB ;
reg  RNC ;
reg  RND ;
reg  RNK ;
reg  RNL ;
reg  RNM ;
reg  RNN ;
reg  RNO ;
reg  RNP ;
reg  rqa ;
reg  RQB ;
reg  rqc ;
reg  RRA ;
reg  RRB ;
reg  RRC ;
reg  RRD ;
reg  RRE ;
reg  RRF ;
reg  rrg ;
reg  RRH ;
reg  RSA ;
reg  RSB ;
reg  RSC ;
wire  aaa ;
wire  aab ;
wire  aac ;
wire  aad ;
wire  aae ;
wire  aaf ;
wire  aag ;
wire  aah ;
wire  aai ;
wire  aaj ;
wire  aak ;
wire  aal ;
wire  aam ;
wire  aan ;
wire  aao ;
wire  aap ;
wire  aba ;
wire  abb ;
wire  abc ;
wire  abd ;
wire  abe ;
wire  abf ;
wire  abg ;
wire  abh ;
wire  abi ;
wire  abj ;
wire  abk ;
wire  abl ;
wire  abm ;
wire  abn ;
wire  abo ;
wire  abp ;
wire  ACH ;
wire  ACI ;
wire  ACJ ;
wire  ACK ;
wire  ACL ;
wire  ACM ;
wire  ACN ;
wire  ACO ;
wire  ACP ;
wire  ADA ;
wire  ADB ;
wire  ADC ;
wire  ADD ;
wire  ADE ;
wire  ADF ;
wire  ADG ;
wire  ADH ;
wire  ADI ;
wire  ADJ ;
wire  ADK ;
wire  ADL ;
wire  ADM ;
wire  ADN ;
wire  ADO ;
wire  aeh ;
wire  aei ;
wire  aej ;
wire  aek ;
wire  ael ;
wire  aem ;
wire  aen ;
wire  aeo ;
wire  aep ;
wire  afa ;
wire  afb ;
wire  afc ;
wire  afd ;
wire  afe ;
wire  aff ;
wire  afg ;
wire  afh ;
wire  afi ;
wire  afj ;
wire  afk ;
wire  afl ;
wire  afm ;
wire  afn ;
wire  afo ;
wire  agh ;
wire  agi ;
wire  agj ;
wire  agk ;
wire  agl ;
wire  agm ;
wire  agn ;
wire  ago ;
wire  agp ;
wire  aha ;
wire  ahb ;
wire  ahc ;
wire  ahd ;
wire  ahe ;
wire  ahf ;
wire  ahg ;
wire  ahh ;
wire  ahi ;
wire  ahj ;
wire  ahk ;
wire  ahl ;
wire  ahm ;
wire  ahn ;
wire  aho ;
wire  aih ;
wire  aii ;
wire  aij ;
wire  aik ;
wire  ail ;
wire  aim ;
wire  ain ;
wire  aio ;
wire  aip ;
wire  aja ;
wire  ajb ;
wire  ajc ;
wire  ajd ;
wire  aje ;
wire  ajf ;
wire  ajg ;
wire  ajh ;
wire  aji ;
wire  ajj ;
wire  ajk ;
wire  ajl ;
wire  ajm ;
wire  ajn ;
wire  ajo ;
wire  akh ;
wire  aki ;
wire  akj ;
wire  akk ;
wire  akl ;
wire  akm ;
wire  akn ;
wire  ako ;
wire  akp ;
wire  ala ;
wire  alb ;
wire  alc ;
wire  ald ;
wire  ale ;
wire  alf ;
wire  alg ;
wire  alh ;
wire  ali ;
wire  alj ;
wire  alk ;
wire  all ;
wire  alm ;
wire  aln ;
wire  alo ;
wire  amh ;
wire  ami ;
wire  amj ;
wire  amk ;
wire  aml ;
wire  amm ;
wire  amn ;
wire  amo ;
wire  amp ;
wire  ana ;
wire  anb ;
wire  anc ;
wire  andd  ;
wire  ane ;
wire  anf ;
wire  ang ;
wire  anh ;
wire  ani ;
wire  anj ;
wire  ank ;
wire  anl ;
wire  anm ;
wire  ann ;
wire  ano ;
wire  aoh ;
wire  aoi ;
wire  aoj ;
wire  aok ;
wire  aol ;
wire  aom ;
wire  aon ;
wire  aoo ;
wire  aop ;
wire  apa ;
wire  apb ;
wire  apc ;
wire  apd ;
wire  ape ;
wire  apf ;
wire  apg ;
wire  aph ;
wire  api ;
wire  apj ;
wire  apk ;
wire  apl ;
wire  apm ;
wire  apn ;
wire  apo ;
wire  aqh ;
wire  aqi ;
wire  aqj ;
wire  aqk ;
wire  aql ;
wire  aqm ;
wire  aqn ;
wire  aqo ;
wire  aqp ;
wire  ara ;
wire  arb ;
wire  arc ;
wire  ard ;
wire  are ;
wire  arf ;
wire  arg ;
wire  arh ;
wire  ari ;
wire  arj ;
wire  ark ;
wire  arl ;
wire  arm ;
wire  arn ;
wire  aro ;
wire  ash ;
wire  asi ;
wire  asj ;
wire  ask ;
wire  asl ;
wire  asm ;
wire  asn ;
wire  aso ;
wire  asp ;
wire  ata ;
wire  atb ;
wire  atc ;
wire  atd ;
wire  ate ;
wire  atf ;
wire  atg ;
wire  ath ;
wire  ati ;
wire  atj ;
wire  atk ;
wire  atl ;
wire  atm ;
wire  atn ;
wire  ato ;
wire  atp ;
wire  bah ;
wire  bai ;
wire  baj ;
wire  bak ;
wire  bal ;
wire  bam ;
wire  ban ;
wire  bao ;
wire  bap ;
wire  bba ;
wire  bbb ;
wire  bbc ;
wire  bbd ;
wire  bbe ;
wire  bbf ;
wire  bbg ;
wire  bbh ;
wire  bbi ;
wire  bbj ;
wire  bbk ;
wire  bbl ;
wire  bbm ;
wire  bbn ;
wire  bbo ;
wire  bbp ;
wire  bci ;
wire  bcj ;
wire  bck ;
wire  bcm ;
wire  bcn ;
wire  bco ;
wire  bda ;
wire  bdb ;
wire  bdc ;
wire  bde ;
wire  bdf ;
wire  bdg ;
wire  bdi ;
wire  bdj ;
wire  bdk ;
wire  bdm ;
wire  bdn ;
wire  bdo ;
wire  beh ;
wire  bei ;
wire  bej ;
wire  bek ;
wire  bel ;
wire  bem ;
wire  ben ;
wire  beo ;
wire  bep ;
wire  bfa ;
wire  bfb ;
wire  bfc ;
wire  bfd ;
wire  bfe ;
wire  bff ;
wire  bfg ;
wire  bfh ;
wire  bfi ;
wire  bfj ;
wire  bfk ;
wire  bfl ;
wire  bga ;
wire  BGA ;
wire  bgb ;
wire  BGB ;
wire  bgc ;
wire  BGC ;
wire  bgd ;
wire  BGD ;
wire  bge ;
wire  BGE ;
wire  bgf ;
wire  BGF ;
wire  bgg ;
wire  BGG ;
wire  bgh ;
wire  BGH ;
wire  bha ;
wire  BHA ;
wire  bhb ;
wire  BHB ;
wire  bhc ;
wire  BHC ;
wire  bhd ;
wire  BHD ;
wire  bhe ;
wire  BHE ;
wire  bhf ;
wire  BHF ;
wire  bhg ;
wire  BHG ;
wire  bhh ;
wire  BHH ;
wire  bia ;
wire  BIA ;
wire  bib ;
wire  BIB ;
wire  bic ;
wire  BIC ;
wire  bid ;
wire  BID ;
wire  bie ;
wire  BIE ;
wire  bif ;
wire  BIF ;
wire  big ;
wire  BIG ;
wire  bih ;
wire  BIH ;
wire  bja ;
wire  BJA ;
wire  bjb ;
wire  BJB ;
wire  bjc ;
wire  BJC ;
wire  bjd ;
wire  BJD ;
wire  bje ;
wire  BJE ;
wire  bjf ;
wire  BJF ;
wire  bjg ;
wire  BJG ;
wire  bjh ;
wire  BJH ;
wire  bka ;
wire  BKA ;
wire  bkb ;
wire  BKB ;
wire  bkc ;
wire  BKC ;
wire  bkd ;
wire  BKD ;
wire  bke ;
wire  BKE ;
wire  bkf ;
wire  BKF ;
wire  bkg ;
wire  BKG ;
wire  bkh ;
wire  BKH ;
wire  bla ;
wire  BLA ;
wire  blb ;
wire  BLB ;
wire  blc ;
wire  BLC ;
wire  bld ;
wire  BLD ;
wire  ble ;
wire  BLE ;
wire  blf ;
wire  BLF ;
wire  blg ;
wire  BLG ;
wire  blh ;
wire  BLH ;
wire  bma ;
wire  BMA ;
wire  bmb ;
wire  BMB ;
wire  bmc ;
wire  BMC ;
wire  bmd ;
wire  BMD ;
wire  bme ;
wire  BME ;
wire  bmf ;
wire  BMF ;
wire  bmg ;
wire  BMG ;
wire  bmh ;
wire  BMH ;
wire  bna ;
wire  BNA ;
wire  bnb ;
wire  BNB ;
wire  bnc ;
wire  BNC ;
wire  bnd ;
wire  BND ;
wire  bne ;
wire  BNE ;
wire  bnf ;
wire  BNF ;
wire  bng ;
wire  BNG ;
wire  bnh ;
wire  BNH ;
wire  caa ;
wire  cab ;
wire  cac ;
wire  cca ;
wire  ccb ;
wire  cda ;
wire  cdb ;
wire  cea ;
wire  ceb ;
wire  cfa ;
wire  cfb ;
wire  cga ;
wire  cgb ;
wire  cha ;
wire  chb ;
wire  cia ;
wire  cib ;
wire  cja ;
wire  cjb ;
wire  daa ;
wire  dab ;
wire  dac ;
wire  dad ;
wire  dae ;
wire  daf ;
wire  dag ;
wire  dah ;
wire  dai ;
wire  daj ;
wire  dak ;
wire  dal ;
wire  dam ;
wire  dan ;
wire  dao ;
wire  dap ;
wire  dba ;
wire  dbb ;
wire  dbc ;
wire  dbd ;
wire  dbe ;
wire  dbf ;
wire  dbg ;
wire  dbh ;
wire  dbi ;
wire  dbj ;
wire  dbk ;
wire  dbl ;
wire  dbm ;
wire  dbn ;
wire  dbo ;
wire  dbp ;
wire  EAA ;
wire  EAB ;
wire  EAC ;
wire  EAD ;
wire  EAE ;
wire  EAF ;
wire  EAG ;
wire  EAH ;
wire  EAI ;
wire  EAJ ;
wire  EAK ;
wire  EAL ;
wire  EAM ;
wire  EAN ;
wire  EAO ;
wire  EAP ;
wire  EBJ ;
wire  EBK ;
wire  EBL ;
wire  EBP ;
wire  ECI ;
wire  ECJ ;
wire  ECK ;
wire  ECL ;
wire  ECM ;
wire  ECN ;
wire  ECO ;
wire  eda ;
wire  edb ;
wire  edc ;
wire  edd ;
wire  ede ;
wire  edf ;
wire  edg ;
wire  edh ;
wire  edi ;
wire  edj ;
wire  edk ;
wire  edl ;
wire  edm ;
wire  edn ;
wire  edo ;
wire  edp ;
wire  faa ;
wire  FAA ;
wire  fab ;
wire  FAB ;
wire  fac ;
wire  FAC ;
wire  fad ;
wire  FAD ;
wire  fae ;
wire  FAE ;
wire  faf ;
wire  FAF ;
wire  fag ;
wire  FAG ;
wire  fah ;
wire  FAH ;
wire  fai ;
wire  FAI ;
wire  faj ;
wire  FAJ ;
wire  fak ;
wire  FAK ;
wire  fal ;
wire  FAL ;
wire  fap ;
wire  FAP ;
wire  fba ;
wire  FBA ;
wire  fbb ;
wire  FBB ;
wire  fbc ;
wire  FBC ;
wire  fbd ;
wire  FBD ;
wire  fbe ;
wire  FBE ;
wire  fbg ;
wire  FBG ;
wire  fbh ;
wire  FBH ;
wire  GAA ;
wire  GAB ;
wire  GAC ;
wire  gae ;
wire  GAF ;
wire  GAG ;
wire  GAH ;
wire  GAI ;
wire  GAL ;
wire  GAM ;
wire  GAN ;
wire  GAO ;
wire  GAP ;
wire  GBA ;
wire  GBC ;
wire  GBD ;
wire  GBE ;
wire  GBF ;
wire  GBG ;
wire  GBH ;
wire  GBI ;
wire  GBJ ;
wire  GBK ;
wire  GBM ;
wire  GBN ;
wire  GBO ;
wire  GBP ;
wire  GCA ;
wire  GCB ;
wire  GCC ;
wire  GCD ;
wire  GCH ;
wire  GCI ;
wire  GCJ ;
wire  GCK ;
wire  GCL ;
wire  GCM ;
wire  GCN ;
wire  gda ;
wire  gdb ;
wire  gdc ;
wire  gdd ;
wire  gde ;
wire  gdf ;
wire  gdg ;
wire  gdh ;
wire  gdi ;
wire  gdj ;
wire  gdk ;
wire  gdl ;
wire  gdx ;
wire  gdy ;
wire  HAA ;
wire  HAB ;
wire  HAC ;
wire  HAD ;
wire  hae ;
wire  haf ;
wire  hag ;
wire  hah ;
wire  HBA ;
wire  HBB ;
wire  HBC ;
wire  HBD ;
wire  HBE ;
wire  HBF ;
wire  HBG ;
wire  HBH ;
wire  HCA ;
wire  HCB ;
wire  HCC ;
wire  HCD ;
wire  HCE ;
wire  HCF ;
wire  HCG ;
wire  HCH ;
wire  HDA ;
wire  HDB ;
wire  HDC ;
wire  HDD ;
wire  HDE ;
wire  HDF ;
wire  HDH ;
wire  hdi ;
wire  hdj ;
wire  hdk ;
wire  hdl ;
wire  HEA ;
wire  HEB ;
wire  HEH ;
wire  hei ;
wire  hej ;
wire  heo ;
wire  hep ;
wire  hfm ;
wire  hfn ;
wire  hia ;
wire  hib ;
wire  hic ;
wire  hja ;
wire  hjb ;
wire  hjc ;
wire  hka ;
wire  hkb ;
wire  hkc ;
wire  hla ;
wire  hlb ;
wire  hlc ;
wire  hma ;
wire  hmb ;
wire  hmc ;
wire  hna ;
wire  hnb ;
wire  hnc ;
wire  hoa ;
wire  hob ;
wire  hoc ;
wire  hpa ;
wire  hpb ;
wire  hpc ;
wire  iaa ;
wire  iab ;
wire  iac ;
wire  iad ;
wire  iae ;
wire  iaf ;
wire  iag ;
wire  iah ;
wire  iai ;
wire  iaj ;
wire  iak ;
wire  ial ;
wire  iam ;
wire  ian ;
wire  iao ;
wire  iap ;
wire  iba ;
wire  ibb ;
wire  ibc ;
wire  ibd ;
wire  ibe ;
wire  ibf ;
wire  ibg ;
wire  ibh ;
wire  ibi ;
wire  ibj ;
wire  ibk ;
wire  ibl ;
wire  ibm ;
wire  ibn ;
wire  ibo ;
wire  ibp ;
wire  ica ;
wire  icb ;
wire  icc ;
wire  icd ;
wire  ice ;
wire  icf ;
wire  icg ;
wire  ich ;
wire  ici ;
wire  icj ;
wire  ick ;
wire  icl ;
wire  icm ;
wire  icn ;
wire  ico ;
wire  icp ;
wire  ida ;
wire  idb ;
wire  idc ;
wire  idd ;
wire  ide ;
wire  idf ;
wire  idg ;
wire  idh ;
wire  idi ;
wire  idj ;
wire  idk ;
wire  idl ;
wire  idm ;
wire  idn ;
wire  ido ;
wire  idp ;
wire  iea ;
wire  ieb ;
wire  iec ;
wire  ied ;
wire  iee ;
wire  ief ;
wire  ieg ;
wire  ieh ;
wire  iei ;
wire  iej ;
wire  iek ;
wire  iel ;
wire  iem ;
wire  ien ;
wire  ieo ;
wire  iep ;
wire  ifa ;
wire  ifb ;
wire  ifc ;
wire  ifd ;
wire  ife ;
wire  ifff  ;
wire  ifg ;
wire  ifh ;
wire  ifi ;
wire  iga ;
wire  igb ;
wire  igc ;
wire  ihb ;
wire  ihc ;
wire  ija ;
wire  ijb ;
wire  ijc ;
wire  ijd ;
wire  ika ;
wire  ikb ;
wire  ila ;
wire  ilb ;
wire  ilc ;
wire  ima ;
wire  imb ;
wire  imc ;
wire  imd ;
wire  ime ;
wire  imf ;
wire  img ;
wire  ina ;
wire  ioa ;
wire  iob ;
wire  ioc ;
wire  iod ;
wire  ipa ;
wire  ipb ;
wire  ipc ;
wire  ipd ;
wire  ipe ;
wire  ipf ;
wire  iqa ;
wire  iqb ;
wire  iqc ;
wire  iqd ;
wire  iqe ;
wire  iqf ;
wire  iqg ;
wire  iqh ;
wire  iqi ;
wire  izz ;
wire  jaa ;
wire  JAA ;
wire  jab ;
wire  JAB ;
wire  jac ;
wire  JAC ;
wire  jad ;
wire  JAD ;
wire  jae ;
wire  JAE ;
wire  jaf ;
wire  JAF ;
wire  jag ;
wire  JAG ;
wire  jam ;
wire  JAM ;
wire  jan ;
wire  JAN ;
wire  jao ;
wire  JAO ;
wire  jap ;
wire  JAP ;
wire  jaq ;
wire  JAQ ;
wire  jbb ;
wire  JBB ;
wire  jbc ;
wire  JBC ;
wire  jbd ;
wire  JBD ;
wire  jbe ;
wire  JBE ;
wire  jbg ;
wire  JBG ;
wire  jbo ;
wire  JBO ;
wire  jbx ;
wire  JBX ;
wire  jby ;
wire  JBY ;
wire  jca ;
wire  JCA ;
wire  jcb ;
wire  JCB ;
wire  jcc ;
wire  JCC ;
wire  jcd ;
wire  JCD ;
wire  jce ;
wire  JCE ;
wire  jcf ;
wire  JCF ;
wire  jcg ;
wire  JCG ;
wire  jch ;
wire  JCH ;
wire  jci ;
wire  JCI ;
wire  jcj ;
wire  JCJ ;
wire  jck ;
wire  JCK ;
wire  jcl ;
wire  JCL ;
wire  jcm ;
wire  JCM ;
wire  jcn ;
wire  JCN ;
wire  jco ;
wire  JCO ;
wire  jcp ;
wire  JCP ;
wire  jcq ;
wire  JCQ ;
wire  jcr ;
wire  JCR ;
wire  jcs ;
wire  JCS ;
wire  jct ;
wire  JCT ;
wire  jcu ;
wire  JCU ;
wire  jcv ;
wire  JCV ;
wire  jcw ;
wire  JCW ;
wire  jcx ;
wire  JCX ;
wire  jcy ;
wire  JCY ;
wire  jcz ;
wire  JCZ ;
wire  jda ;
wire  JDA ;
wire  jdb ;
wire  JDB ;
wire  jdc ;
wire  JDC ;
wire  jdd ;
wire  JDD ;
wire  jde ;
wire  JDE ;
wire  jdf ;
wire  JDF ;
wire  jdh ;
wire  JDH ;
wire  jdi ;
wire  JDI ;
wire  jdj ;
wire  JDJ ;
wire  jdk ;
wire  JDK ;
wire  jdl ;
wire  JDL ;
wire  jdm ;
wire  JDM ;
wire  jdn ;
wire  JDN ;
wire  jdo ;
wire  JDO ;
wire  jdp ;
wire  JDP ;
wire  jea ;
wire  JEA ;
wire  jeb ;
wire  JEB ;
wire  jec ;
wire  JEC ;
wire  jed ;
wire  JED ;
wire  jee ;
wire  JEE ;
wire  jef ;
wire  JEF ;
wire  jeg ;
wire  JEG ;
wire  jeh ;
wire  JEH ;
wire  jei ;
wire  JEI ;
wire  jej ;
wire  JEJ ;
wire  jek ;
wire  JEK ;
wire  jel ;
wire  JEL ;
wire  jem ;
wire  JEM ;
wire  jen ;
wire  JEN ;
wire  jeo ;
wire  JEO ;
wire  jep ;
wire  JEP ;
wire  jfa ;
wire  JFA ;
wire  jfb ;
wire  JFB ;
wire  jfc ;
wire  JFC ;
wire  jfd ;
wire  JFD ;
wire  jfe ;
wire  JFE ;
wire  jff ;
wire  JFF ;
wire  jfg ;
wire  JFG ;
wire  jfh ;
wire  JFH ;
wire  jfi ;
wire  JFI ;
wire  jfj ;
wire  JFJ ;
wire  jfx ;
wire  JFX ;
wire  jfy ;
wire  JFY ;
wire  jga ;
wire  JGA ;
wire  jgb ;
wire  JGB ;
wire  jgc ;
wire  JGC ;
wire  jgd ;
wire  JGD ;
wire  jge ;
wire  JGE ;
wire  jgf ;
wire  JGF ;
wire  jgg ;
wire  JGG ;
wire  jgh ;
wire  JGH ;
wire  jgi ;
wire  JGI ;
wire  jgj ;
wire  JGJ ;
wire  jgk ;
wire  JGK ;
wire  jgl ;
wire  JGL ;
wire  jgm ;
wire  JGM ;
wire  jgn ;
wire  JGN ;
wire  jgo ;
wire  JGO ;
wire  jgp ;
wire  JGP ;
wire  jha ;
wire  JHA ;
wire  jhb ;
wire  JHB ;
wire  jhc ;
wire  JHC ;
wire  jhd ;
wire  JHD ;
wire  jhe ;
wire  JHE ;
wire  jhf ;
wire  JHF ;
wire  jhg ;
wire  JHG ;
wire  jhh ;
wire  JHH ;
wire  jhi ;
wire  JHI ;
wire  jhj ;
wire  JHJ ;
wire  jhk ;
wire  JHK ;
wire  jhl ;
wire  JHL ;
wire  jhm ;
wire  JHM ;
wire  jhn ;
wire  JHN ;
wire  jho ;
wire  JHO ;
wire  jhp ;
wire  JHP ;
wire  jia ;
wire  JIA ;
wire  jic ;
wire  JIC ;
wire  jid ;
wire  JID ;
wire  jie ;
wire  JIE ;
wire  jjb ;
wire  JJB ;
wire  jjc ;
wire  JJC ;
wire  jjd ;
wire  JJD ;
wire  jje ;
wire  JJE ;
wire  jjg ;
wire  JJG ;
wire  jjh ;
wire  JJH ;
wire  jjk ;
wire  JJK ;
wire  jjl ;
wire  JJL ;
wire  jjp ;
wire  JJP ;
wire  jka ;
wire  JKA ;
wire  jkb ;
wire  JKB ;
wire  jkc ;
wire  JKC ;
wire  jkd ;
wire  JKD ;
wire  jke ;
wire  JKE ;
wire  jla ;
wire  JLA ;
wire  jlb ;
wire  JLB ;
wire  jlc ;
wire  JLC ;
wire  jld ;
wire  JLD ;
wire  jle ;
wire  JLE ;
wire  jlf ;
wire  JLF ;
wire  jlg ;
wire  JLG ;
wire  jma ;
wire  JMA ;
wire  jmb ;
wire  JMB ;
wire  jna ;
wire  JNA ;
wire  jnb ;
wire  JNB ;
wire  jnc ;
wire  JNC ;
wire  jnd ;
wire  JND ;
wire  jne ;
wire  JNE ;
wire  joa ;
wire  JOA ;
wire  job ;
wire  JOB ;
wire  joc ;
wire  JOC ;
wire  jod ;
wire  JOD ;
wire  joe ;
wire  JOE ;
wire  jof ;
wire  JOF ;
wire  jog ;
wire  JOG ;
wire  joh ;
wire  JOH ;
wire  joj ;
wire  JOJ ;
wire  jok ;
wire  JOK ;
wire  jol ;
wire  JOL ;
wire  joo ;
wire  JOO ;
wire  jop ;
wire  JOP ;
wire  jox ;
wire  JOX ;
wire  jpa ;
wire  JPA ;
wire  jqa ;
wire  JQA ;
wire  jqb ;
wire  JQB ;
wire  jqc ;
wire  JQC ;
wire  jqe ;
wire  JQE ;
wire  jqf ;
wire  JQF ;
wire  jqh ;
wire  JQH ;
wire  jqi ;
wire  JQI ;
wire  jqj ;
wire  JQJ ;
wire  jra ;
wire  JRA ;
wire  jrb ;
wire  JRB ;
wire  jrc ;
wire  JRC ;
wire  jrd ;
wire  JRD ;
wire  jre ;
wire  JRE ;
wire  jrf ;
wire  JRF ;
wire  jsa ;
wire  JSA ;
wire  jsb ;
wire  JSB ;
wire  jsc ;
wire  JSC ;
wire  jsd ;
wire  JSD ;
wire  jse ;
wire  JSE ;
wire  jtb ;
wire  JTB ;
wire  jua ;
wire  JUA ;
wire  jva ;
wire  JVA ;
wire  jvb ;
wire  JVB ;
wire  jvc ;
wire  JVC ;
wire  jvd ;
wire  JVD ;
wire  jxa ;
wire  JXA ;
wire  jxb ;
wire  JXB ;
wire  kaa ;
wire  kab ;
wire  kac ;
wire  kad ;
wire  kae ;
wire  kaf ;
wire  laa ;
wire  lab ;
wire  lac ;
wire  lad ;
wire  lae ;
wire  laf ;
wire  lba ;
wire  lbb ;
wire  lbc ;
wire  lbd ;
wire  lbe ;
wire  lbf ;
wire  maa ;
wire  mab ;
wire  mac ;
wire  naa ;
wire  nab ;
wire  nac ;
wire  nad ;
wire  nae ;
wire  nba ;
wire  nbb ;
wire  nbc ;
wire  nbd ;
wire  nca ;
wire  ncb ;
wire  oaa ;
wire  oab ;
wire  oac ;
wire  oad ;
wire  oae ;
wire  oaf ;
wire  oag ;
wire  oah ;
wire  oai ;
wire  oaj ;
wire  oak ;
wire  oal ;
wire  oam ;
wire  oan ;
wire  oao ;
wire  oap ;
wire  oba ;
wire  obb ;
wire  obc ;
wire  obd ;
wire  obe ;
wire  obf ;
wire  obg ;
wire  obh ;
wire  obi ;
wire  obj ;
wire  obk ;
wire  obl ;
wire  obm ;
wire  obn ;
wire  obo ;
wire  obp ;
wire  OCA ;
wire  OCB ;
wire  OCC ;
wire  OCD ;
wire  OCE ;
wire  OCF ;
wire  OCG ;
wire  OCH ;
wire  OCI ;
wire  OCJ ;
wire  OCK ;
wire  OCL ;
wire  OCM ;
wire  OCN ;
wire  OCO ;
wire  OCP ;
wire  ODA ;
wire  ODB ;
wire  ODC ;
wire  ODD ;
wire  ODE ;
wire  ODF ;
wire  ODG ;
wire  ODH ;
wire  ODI ;
wire  ODJ ;
wire  ODK ;
wire  ODL ;
wire  ODM ;
wire  ODN ;
wire  ODO ;
wire  ODP ;
wire  oea ;
wire  oeb ;
wire  oec ;
wire  oed ;
wire  oee ;
wire  oef ;
wire  oeg ;
wire  oeh ;
wire  OEI ;
wire  oej ;
wire  oek ;
wire  oel ;
wire  oem ;
wire  oen ;
wire  oeo ;
wire  oep ;
wire  OEQ ;
wire  OER ;
wire  oes ;
wire  oet ;
wire  oeu ;
wire  oev ;
wire  oew ;
wire  oex ;
wire  oey ;
wire  ofa ;
wire  OFB ;
wire  ofc ;
wire  oga ;
wire  ogb ;
wire  ogc ;
wire  ogd ;
wire  oge ;
wire  ogf ;
wire  ogg ;
wire  ogh ;
wire  ogi ;
wire  ogj ;
wire  oha ;
wire  ohb ;
wire  ohc ;
wire  ohd ;
wire  ohe ;
wire  oia ;
wire  OIB ;
wire  oic ;
wire  oid ;
wire  oie ;
wire  OIG ;
wire  oja ;
wire  ojb ;
wire  ojc ;
wire  ojd ;
wire  oje ;
wire  oka ;
wire  okb ;
wire  ola ;
wire  olb ;
wire  olc ;
wire  OLD ;
wire  olf ;
wire  oma ;
wire  omb ;
wire  OQA ;
wire  oqb ;
wire  ORA ;
wire  ORB ;
wire  ORC ;
wire  ORD ;
wire  ORE ;
wire  ORF ;
wire  ota ;
wire  otb ;
wire  otc ;
wire  OTD ;
wire  OTE ;
wire  OTF ;
wire  paa ;
wire  pab ;
wire  pac ;
wire  pad ;
wire  pae ;
wire  paf ;
wire  pag ;
wire  pah ;
wire  pai ;
wire  paj ;
wire  pak ;
wire  pal ;
wire  pam ;
wire  pan ;
wire  pao ;
wire  pap ;
wire  pba ;
wire  pbb ;
wire  pbc ;
wire  pbd ;
wire  pbe ;
wire  pbf ;
wire  pbg ;
wire  pbh ;
wire  pbi ;
wire  pbj ;
wire  pbk ;
wire  pbl ;
wire  pbm ;
wire  pbn ;
wire  pbo ;
wire  pbp ;
wire  pca ;
wire  pcb ;
wire  pcc ;
wire  pcd ;
wire  pce ;
wire  pcf ;
wire  pcg ;
wire  pch ;
wire  pci ;
wire  pcj ;
wire  pck ;
wire  pcl ;
wire  pcm ;
wire  pcn ;
wire  pco ;
wire  pcp ;
wire  pda ;
wire  pdb ;
wire  pdc ;
wire  pdd ;
wire  pde ;
wire  pdf ;
wire  pdg ;
wire  pdh ;
wire  pdi ;
wire  pdj ;
wire  pdk ;
wire  pdl ;
wire  pdm ;
wire  pdn ;
wire  pdo ;
wire  pdp ;
wire  peb ;
wire  pec ;
wire  ped ;
wire  pee ;
wire  pef ;
wire  peg ;
wire  peh ;
wire  pei ;
wire  pej ;
wire  pek ;
wire  pel ;
wire  pem ;
wire  pen ;
wire  peo ;
wire  pep ;
wire  pfa ;
wire  pfb ;
wire  pfc ;
wire  pfd ;
wire  pfe ;
wire  pff ;
wire  pfg ;
wire  pfh ;
wire  pfi ;
wire  pfj ;
wire  pfk ;
wire  pfl ;
wire  qaa ;
wire  qab ;
wire  qac ;
wire  qad ;
wire  qba ;
wire  qcd ;
wire  qch ;
wire  qci ;
wire  qcj ;
wire  QCK ;
wire  qcx ;
wire  qcy ;
wire  qcz ;
wire  qea ;
wire  qeb ;
wire  qfa ;
wire  qfb ;
wire  qfc ;
wire  qga ;
wire  qgb ;
wire  QGD ;
wire  qge ;
wire  qha ;
wire  qhc ;
wire  qhd ;
wire  qhe ;
wire  qhf ;
wire  QIA ;
wire  QIB ;
wire  QIC ;
wire  QID ;
wire  qka ;
wire  qkb ;
wire  qkc ;
wire  qkd ;
wire  qke ;
wire  qkf ;
wire  qkg ;
wire  qkh ;
wire  qkj ;
wire  qkk ;
wire  qkl ;
wire  qkm ;
wire  qkn ;
wire  qko ;
wire  qkp ;
wire  qkq ;
wire  qkr ;
wire  qks ;
wire  qkt ;
wire  qkw ;
wire  qkx ;
wire  qky ;
wire  qla ;
wire  qlb ;
wire  qlc ;
wire  qld ;
wire  qle ;
wire  qlf ;
wire  qlg ;
wire  qli ;
wire  qlj ;
wire  qlk ;
wire  qll ;
wire  qlm ;
wire  qln ;
wire  qlo ;
wire  qlp ;
wire  qlq ;
wire  qlr ;
wire  qls ;
wire  QLX ;
wire  qma ;
wire  QMB ;
wire  QMC ;
wire  qme ;
wire  QMF ;
wire  QMG ;
wire  qmi ;
wire  QMJ ;
wire  qmk ;
wire  qml ;
wire  QNA ;
wire  QNB ;
wire  QNC ;
wire  qnd ;
wire  QNE ;
wire  QNF ;
wire  QNG ;
wire  qni ;
wire  QNJ ;
wire  qnm ;
wire  QNN ;
wire  qnq ;
wire  QNR ;
wire  qnu ;
wire  QNV ;
wire  QOA ;
wire  qpa ;
wire  qpb ;
wire  qpc ;
wire  qpd ;
wire  qqa ;
wire  qqb ;
wire  qqc ;
wire  qqd ;
wire  qqe ;
wire  qqf ;
wire  qqg ;
wire  qqh ;
wire  qqi ;
wire  qqj ;
wire  qqk ;
wire  qql ;
wire  qqm ;
wire  qqn ;
wire  qqo ;
wire  qqp ;
wire  qqq ;
wire  qqr ;
wire  qqs ;
wire  qqt ;
wire  qqw ;
wire  QQX ;
wire  qqy ;
wire  qqz ;
wire  qra ;
wire  qrb ;
wire  qrc ;
wire  qrd ;
wire  qre ;
wire  qrf ;
wire  qsa ;
wire  qsb ;
wire  qsc ;
wire  qsd ;
wire  qse ;
wire  qsf ;
wire  qsg ;
wire  qsh ;
wire  QSI ;
wire  qta ;
wire  QTB ;
wire  qtc ;
wire  qtd ;
wire  qte ;
wire  qtf ;
wire  qtg ;
wire  qth ;
wire  qti ;
wire  qtj ;
wire  qtm ;
wire  qtn ;
wire  qto ;
wire  qtp ;
wire  QTQ ;
wire  QTR ;
wire  qtw ;
wire  qtx ;
wire  qua ;
wire  qub ;
wire  quc ;
wire  qud ;
wire  que ;
wire  quf ;
wire  QVA ;
wire  QVB ;
wire  QVC ;
wire  QVD ;
wire  QVE ;
wire  QVF ;
wire  QVG ;
wire  QVH ;
wire  QVI ;
wire  QVJ ;
wire  qwa ;
wire  qwb ;
wire  qwc ;
wire  QWD ;
wire  QWE ;
wire  QWF ;
wire  QWG ;
wire  QWH ;
wire  QWI ;
wire  qwj ;
wire  qxa ;
wire  qxb ;
wire  qxc ;
wire  qxd ;
wire  qxe ;
wire  qxf ;
wire  qya ;
wire  qyb ;
wire  qyc ;
wire  qyd ;
wire  QZA ;
wire  QZD ;
wire  qze ;
wire  qzf ;
wire  RAA ;
wire  rab ;
wire  rac ;
wire  rad ;
wire  rae ;
wire  raf ;
wire  rag ;
wire  RAT ;
wire  rax ;
wire  RBA ;
wire  rbb ;
wire  rbc ;
wire  rbd ;
wire  rbe ;
wire  rbf ;
wire  rbg ;
wire  rbh ;
wire  rbi ;
wire  rbx ;
wire  rec ;
wire  rfa ;
wire  rfb ;
wire  rga ;
wire  rgb ;
wire  rgc ;
wire  rgd ;
wire  rha ;
wire  rhb ;
wire  rhc ;
wire  rhd ;
wire  rhe ;
wire  rhf ;
wire  rhg ;
wire  rhh ;
wire  rhi ;
wire  rhj ;
wire  ria ;
wire  rib ;
wire  ric ;
wire  rid ;
wire  rie ;
wire  rif ;
wire  rix ;
wire  rja ;
wire  rjb ;
wire  rjc ;
wire  rjd ;
wire  RJE ;
wire  rjf ;
wire  rjg ;
wire  rjh ;
wire  rji ;
wire  rjk ;
wire  rjl ;
wire  rka ;
wire  rkb ;
wire  rkc ;
wire  rkd ;
wire  rla ;
wire  rlb ;
wire  rlc ;
wire  rld ;
wire  rlx ;
wire  rma ;
wire  rmb ;
wire  rmc ;
wire  rmd ;
wire  rme ;
wire  rmf ;
wire  rmg ;
wire  rmh ;
wire  rmi ;
wire  rmj ;
wire  rmk ;
wire  rml ;
wire  rmm ;
wire  rmn ;
wire  rmo ;
wire  rmp ;
wire  rmq ;
wire  rmr ;
wire  rms ;
wire  rmt ;
wire  rmu ;
wire  RMV ;
wire  rna ;
wire  rnb ;
wire  rnc ;
wire  rnd ;
wire  rnk ;
wire  rnl ;
wire  rnm ;
wire  rnn ;
wire  rno ;
wire  rnp ;
wire  RQA ;
wire  rqb ;
wire  RQC ;
wire  rra ;
wire  rrb ;
wire  rrc ;
wire  rrd ;
wire  rre ;
wire  rrf ;
wire  RRG ;
wire  rrh ;
wire  rsa ;
wire  rsb ;
wire  rsc ;
wire  taa ;
wire  TAA ;
wire  tab ;
wire  TAB ;
wire  tac ;
wire  TAC ;
wire  tad ;
wire  TAD ;
wire  tba ;
wire  TBA ;
wire  tbb ;
wire  TBB ;
wire  tbc ;
wire  TBC ;
wire  tbd ;
wire  TBD ;
wire  tca ;
wire  TCA ;
wire  tcb ;
wire  TCB ;
wire  tcc ;
wire  TCC ;
wire  tcd ;
wire  TCD ;
wire  tda ;
wire  TDA ;
wire  tdb ;
wire  TDB ;
wire  tdc ;
wire  TDC ;
wire  tdd ;
wire  TDD ;
wire  tea ;
wire  TEA ;
wire  teb ;
wire  TEB ;
wire  tec ;
wire  TEC ;
wire  ted ;
wire  TED ;
wire  tee ;
wire  TEE ;
wire  tef ;
wire  TEF ;
wire  tfa ;
wire  TFA ;
wire  tfb ;
wire  TFB ;
wire  tfc ;
wire  TFC ;
wire  tfd ;
wire  TFD ;
wire  tga ;
wire  TGA ;
wire  tgb ;
wire  TGB ;
wire  tgc ;
wire  TGC ;
wire  tgd ;
wire  TGD ;
wire  tge ;
wire  TGE ;
wire  tgf ;
wire  TGF ;
wire  tha ;
wire  THA ;
wire  tla ;
wire  TLA ;
wire  tlb ;
wire  TLB ;
wire  tlc ;
wire  TLC ;
wire  tld ;
wire  TLD ;
wire  tma ;
wire  TMA ;
wire  tmb ;
wire  TMB ;
wire  tmc ;
wire  TMC ;
wire  tmd ;
wire  TMD ;
wire  tme ;
wire  TME ;
wire  tpa ;
wire  TPA ;
wire  tpb ;
wire  TPB ;
wire  tpc ;
wire  TPC ;
wire  tpd ;
wire  TPD ;
wire  waa ;
wire  WAA ;
wire  wab ;
wire  WAB ;
wire  wac ;
wire  WAC ;
wire  wad ;
wire  WAD ;
wire  wae ;
wire  WAE ;
wire  waf ;
wire  WAF ;
wire  wag ;
wire  WAG ;
wire  wah ;
wire  WAH ;
wire  wai ;
wire  WAI ;
wire  waj ;
wire  WAJ ;
wire  wak ;
wire  WAK ;
wire  wal ;
wire  WAL ;
wire  wam ;
wire  WAM ;
wire  wan ;
wire  WAN ;
wire  wao ;
wire  WAO ;
wire  wap ;
wire  WAP ;
wire  wba ;
wire  WBA ;
wire  wbb ;
wire  WBB ;
wire  wbc ;
wire  WBC ;
wire  wbd ;
wire  WBD ;
wire  wbe ;
wire  WBE ;
wire  wbf ;
wire  WBF ;
wire  wbg ;
wire  WBG ;
wire  wbh ;
wire  WBH ;
wire  wbi ;
wire  WBI ;
wire  wbj ;
wire  WBJ ;
wire  wbk ;
wire  WBK ;
wire  wbl ;
wire  WBL ;
wire  wbm ;
wire  WBM ;
wire  wbn ;
wire  WBN ;
wire  wbo ;
wire  WBO ;
wire  wbp ;
wire  WBP ;
wire  wca ;
wire  WCA ;
wire  wcb ;
wire  WCB ;
wire  wcc ;
wire  WCC ;
wire  wcd ;
wire  WCD ;
wire  wce ;
wire  WCE ;
wire  wcf ;
wire  WCF ;
wire  wcg ;
wire  WCG ;
wire  wch ;
wire  WCH ;
wire  wci ;
wire  WCI ;
wire  wcj ;
wire  WCJ ;
wire  wck ;
wire  WCK ;
wire  wcl ;
wire  WCL ;
wire  wcm ;
wire  WCM ;
wire  wcn ;
wire  WCN ;
wire  wco ;
wire  WCO ;
wire  wcp ;
wire  WCP ;
wire  wda ;
wire  WDA ;
wire  wdb ;
wire  WDB ;
wire  wdc ;
wire  WDC ;
wire  wdd ;
wire  WDD ;
wire  wde ;
wire  WDE ;
wire  wdf ;
wire  WDF ;
wire  wdg ;
wire  WDG ;
wire  wdh ;
wire  WDH ;
wire  wdi ;
wire  WDI ;
wire  wdj ;
wire  WDJ ;
wire  wdk ;
wire  WDK ;
wire  wdl ;
wire  WDL ;
wire  wdm ;
wire  WDM ;
wire  wdn ;
wire  WDN ;
wire  wdo ;
wire  WDO ;
wire  wdp ;
wire  WDP ;
wire  ZZI ;
wire  ZZO ;
assign ZZI = 1'b1;
assign ZZO = 1'b0;
assign paa = ~PAA;  //complement 
assign pca = ~PCA;  //complement 
assign JGA =  ZZI & ZZI & QVA  ; 
assign jga = ~JGA;  //complement 
assign JPA =  ZZI & paa & QVA  |  qva & PAA  ; 
assign jpa = ~JPA;  //complement 
assign JGI = QVD; 
assign jgi = ~JGI; //complement 
assign JDI = QWD; 
assign jdi = ~JDI;  //complement 
assign pai = ~PAI;  //complement 
assign pci = ~PCI;  //complement 
assign pei = ~PEI;  //complement 
assign QVA = ~qva;  //complement 
assign QVJ = ~qvj;  //complement 
assign bai = ~BAI;  //complement 
assign bci = ~BCI;  //complement 
assign bei = ~BEI;  //complement 
assign HAA = ~haa;  //complement 
assign HAB = ~hab;  //complement 
assign pba = ~PBA;  //complement 
assign pda = ~PDA;  //complement 
assign pfa = ~PFA;  //complement 
assign TPC = QWJ; 
assign tpc = ~TPC; //complement 
assign TPD = QWJ; 
assign tpd = ~TPD;  //complement 
assign TPA = QWJ; 
assign tpa = ~TPA;  //complement 
assign TPB = QWJ; 
assign tpb = ~TPB;  //complement 
assign bba = ~BBA;  //complement 
assign bda = ~BDA;  //complement 
assign bfa = ~BFA;  //complement 
assign HAC = ~hac;  //complement 
assign HAD = ~had;  //complement 
assign pbi = ~PBI;  //complement 
assign pdi = ~PDI;  //complement 
assign pfi = ~PFI;  //complement 
assign JHI =  QVG & QVI  ; 
assign jhi = ~JHI;  //complement  
assign JHA =  QVF  ; 
assign jha = ~JHA;  //complement 
assign bbi = ~BBI;  //complement 
assign bdi = ~BDI;  //complement 
assign bfi = ~BFI;  //complement 
assign JEA = QWF; 
assign jea = ~JEA; //complement 
assign jei = qwh; 
assign JEI = ~jei;  //complement 
assign HBA = ~hba;  //complement 
assign HCA = ~hca;  //complement 
assign HDA = ~hda;  //complement 
assign HEA = ~hea;  //complement 
assign HBB = ~hbb;  //complement 
assign HCB = ~hcb;  //complement 
assign HDB = ~hdb;  //complement 
assign HEB = ~heb;  //complement 
assign HBC = ~hbc;  //complement 
assign HCC = ~hcc;  //complement 
assign HDC = ~hdc;  //complement 
assign HBH = ~hbh;  //complement 
assign HBE = ~hbe;  //complement 
assign HCE = ~hce;  //complement 
assign HDE = ~hde;  //complement 
assign HBD = ~hbd;  //complement 
assign HBF = ~hbf;  //complement 
assign HCF = ~hcf;  //complement 
assign HDF = ~hdf;  //complement 
assign HCD = ~hcd;  //complement 
assign HBG = ~hbg;  //complement 
assign HCG = ~hcg;  //complement 
assign HDD = ~hdd;  //complement 
assign HCH = ~hch;  //complement 
assign HDH = ~hdh;  //complement 
assign HEH = ~heh;  //complement 
assign hae = ~HAE;  //complement 
assign haf = ~HAF;  //complement 
assign hag = ~HAG;  //complement 
assign hah = ~HAH;  //complement 
assign JAD = HDE & HDD ; 
assign jad = ~JAD ; //complement 
assign JAE = HDF & HDA ; 
assign jae = ~JAE ;  //complement 
assign JAF = HDF & HDB; 
assign jaf = ~JAF; 
assign lba = ~LBA;  //complement 
assign ACI = ~aci;  //complement 
assign ADA = ~ada;  //complement 
assign ADI = ~adi;  //complement 
assign BGA =  ach & ASH  |  aai & ACI  |  AAI & aci  |  asj & ACJ  |  ASJ & acj  |  ash & ACH  ;
assign bga = ~BGA;  //complement 
assign cca = ~CCA;  //complement 
assign BGC =  acn & ASN  |  asn & ACN  |  ASO & aco  |  aso & ACO  |  ASP & acp  |  asp & ACP  ;
assign bgc = ~BGC;  //complement 
assign ccb = ~CCB;  //complement 
assign BGE =  add & ATD  |  atd & ADD  |  ATE & ade  |  ate & ADE  |  ATF & adf  |  atf & ADF  ;
assign bge = ~BGE;  //complement 
assign GAA = ~gaa;  //complement 
assign GAI = ~gai;  //complement 
assign GAB = ~gab;  //complement 
assign BGG =  adj & ATJ  |  atj & ADJ  |  ATK & adk  |  atk & ADK  |  ATL & adl  |  atl & ADL  ;
assign bgg = ~BGG;  //complement 
assign GAO = ~gao;  //complement 
assign GBH = ~gbh;  //complement 
assign FAI =  eal & eak & eaj  ; 
assign fai = ~FAI;  //complement  
assign FBA =  ebl & ebk  ; 
assign fba = ~FBA;  //complement 
assign GCI = ~gci;  //complement 
assign GAM = ~gam;  //complement 
assign hdi = ~HDI;  //complement 
assign hdj = ~HDJ;  //complement 
assign hdk = ~HDK;  //complement 
assign hdl = ~HDL;  //complement 
assign qqi = ~QQI;  //complement 
assign qta = ~QTA;  //complement 
assign rja = ~RJA;  //complement 
assign JMA = QOA & ZZI ; 
assign jma = ~JMA ; //complement 
assign JMB = QOA & KAA ; 
assign jmb = ~JMB ;  //complement 
assign qnd = ~QND;  //complement 
assign QOA = ~qoa;  //complement 
assign jaq =  hdf & qtm  ; 
assign JAQ = ~jaq;  //complement 
assign BGB =  ASK & ack  |  ask & ACK  |  ASL & acl  |  asl & ACL  |  ASM & acm  |  asm & ACM  ;
assign bgb = ~BGB;  //complement 
assign aaa = ~AAA;  //complement 
assign WAA =  ZZO & ZZI & qxa  |  AAA & ZZI & QXA  ; 
assign waa = ~WAA;  //complement 
assign WAI =  BAI & ZZI & qxa  |  AAI & ZZI & QXA  ; 
assign wai = ~WAI;  //complement 
assign oaa = ~OAA;  //complement 
assign oai = ~OAI;  //complement 
assign BGD =  ABA & ada  |  aba & ADA  |  ATB & adb  |  atb & ADB  |  ATC & adc  |  atc & ADC  ;
assign bgd = ~BGD;  //complement 
assign asi = ~ASI;  //complement 
assign aai = ~AAI;  //complement 
assign TBA = QZA; 
assign tba = ~TBA; //complement 
assign TBB = QZA; 
assign tbb = ~TBB;  //complement 
assign tbc = qza; 
assign TBC = ~tbc;  //complement 
assign tbd = qza; 
assign TBD = ~tbd;  //complement 
assign wca = aaa; 
assign WCA = ~wca; //complement 
assign wci = aai; 
assign WCI = ~wci;  //complement 
assign wda = aba; 
assign WDA = ~wda;  //complement 
assign wdi = abi; 
assign WDI = ~wdi;  //complement 
assign BGF =  ATG & adg  |  atg & ADG  |  ATH & adh  |  ath & ADH  |  ABI & adi  |  abi & ADI  ;
assign bgf = ~BGF;  //complement 
assign ata = ~ATA;  //complement 
assign aba = ~ABA;  //complement 
assign daa = ~DAA;  //complement 
assign dai = ~DAI;  //complement 
assign dba = ~DBA;  //complement 
assign dbi = ~DBI;  //complement 
assign ORA = ~ora;  //complement 
assign otb = ~OTB;  //complement 
assign edi = ~EDI;  //complement 
assign QZA = ~qza;  //complement 
assign BGH =  ATM & adm  |  atm & ADM  |  ATN & adn  |  atn & ADN  |  ATO & ado  |  ato & ADO  ;
assign bgh = ~BGH;  //complement 
assign ati = ~ATI;  //complement 
assign abi = ~ABI;  //complement 
assign WBA =  BBA & ZZI & qxb  |  ABA & ZZI & QXB  ; 
assign wba = ~WBA;  //complement 
assign WBI =  BBI & ZZI & qxb  |  ABI & ZZI & QXB  ; 
assign wbi = ~WBI;  //complement 
assign oba = ~OBA;  //complement 
assign obi = ~OBI;  //complement 
assign EAA = ~eaa;  //complement 
assign EAI = ~eai;  //complement 
assign ECI = ~eci;  //complement 
assign naa = ~NAA;  //complement 
assign nba = ~NBA;  //complement 
assign nca = ~NCA;  //complement 
assign qze = ~QZE;  //complement 
assign RJE = ~rje;  //complement 
assign qya = ~QYA;  //complement 
assign qyb = ~QYB;  //complement 
assign qyc = ~QYC;  //complement 
assign qyd = ~QYD;  //complement 
assign eda = ~EDA;  //complement 
assign rjd = ~RJD;  //complement 
assign JSC =  QQI & NBA & NBB  ; 
assign jsc = ~JSC;  //complement 
assign JSB =  QQI & NBA  ; 
assign jsb = ~JSB;  //complement 
assign JSA =  QQI  ; 
assign jsa = ~JSA;  //complement 
assign jbx = heo; 
assign JBX = ~jbx; //complement 
assign jby = hep; 
assign JBY = ~jby;  //complement 
assign OCA = ~oca;  //complement 
assign OCI = ~oci;  //complement 
assign ODA = ~oda;  //complement 
assign ODI = ~odi;  //complement 
assign heo = ~HEO;  //complement 
assign hep = ~HEP;  //complement 
assign qge = ~QGE;  //complement 
assign QGD = ~qgd;  //complement 
assign rjk = ~RJK;  //complement 
assign oea = ~OEA;  //complement 
assign QZD = ~qzd;  //complement 
assign rjb = ~RJB;  //complement 
assign qtm = ~QTM;  //complement 
assign kaa = ~KAA;  //complement 
assign JNA =  MAA & ZZI & QNG  |  NCA & ZZI & RQC  ; 
assign jna = ~JNA;  //complement 
assign JNB =  MAB & ZZI & QNG  |  NCB & ZZI & RQC  ; 
assign jnb = ~JNB;  //complement 
assign rjf = ~RJF;  //complement 
assign rjg = ~RJG;  //complement 
assign rjh = ~RJH;  //complement 
assign rji = ~RJI;  //complement 
assign laa = ~LAA;  //complement 
assign pab = ~PAB;  //complement 
assign pcb = ~PCB;  //complement 
assign peb = ~PEB;  //complement 
assign JGB =  QVB  ; 
assign jgb = ~JGB;  //complement  
assign JGJ =  QVD & PCI  ; 
assign jgj = ~JGJ;  //complement 
assign JDJ =  QWD & BCI  ; 
assign jdj = ~JDJ;  //complement 
assign paj = ~PAJ;  //complement 
assign pcj = ~PCJ;  //complement 
assign pej = ~PEJ;  //complement 
assign QVH = ~qvh;  //complement 
assign QVI = ~qvi;  //complement 
assign baj = ~BAJ;  //complement 
assign bcj = ~BCJ;  //complement 
assign bej = ~BEJ;  //complement 
assign pbb = ~PBB;  //complement 
assign pdb = ~PDB;  //complement 
assign pfb = ~PFB;  //complement 
assign JFE =  PFA & PFB & PFC & PFD  ; 
assign jfe = ~JFE;  //complement  
assign JFG =  PFI & PFJ & PFK & PFL  ; 
assign jfg = ~JFG;  //complement 
assign bbb = ~BBB;  //complement 
assign bdb = ~BDB;  //complement 
assign bfb = ~BFB;  //complement 
assign pbj = ~PBJ;  //complement 
assign pdj = ~PDJ;  //complement 
assign pfj = ~PFJ;  //complement 
assign JHJ =  QVG & QVI & PDI  ; 
assign jhj = ~JHJ;  //complement  
assign JHB =  QVF & PDA  ; 
assign jhb = ~JHB;  //complement 
assign bbj = ~BBJ;  //complement 
assign bdj = ~BDJ;  //complement 
assign bfj = ~BFJ;  //complement 
assign JEB =  QWF & BDA  ; 
assign jeb = ~JEB;  //complement 
assign jfi =  gbh & gbi & gbj  ; 
assign JFI = ~jfi;  //complement 
assign JEJ =  QWH & BDI & gbj  ; 
assign jej = ~JEJ;  //complement 
assign rha = ~RHA;  //complement 
assign rhb = ~RHB;  //complement 
assign rhc = ~RHC;  //complement 
assign rhd = ~RHD;  //complement 
assign rhe = ~RHE;  //complement 
assign rhf = ~RHF;  //complement 
assign rhg = ~RHG;  //complement 
assign rhh = ~RHH;  //complement 
assign rhi = ~RHI;  //complement 
assign rhj = ~RHJ;  //complement 
assign qha = ~QHA;  //complement 
assign jid =  rhf & rhg & rhh & rhi & rhj & qhc  ; 
assign JID = ~jid;  //complement  
assign jic =  qha & rha & rhb & rhc & rhd & rhe  ; 
assign JIC = ~jic;  //complement  
assign qkk = ~QKK;  //complement 
assign rid = ~RID;  //complement 
assign rie = ~RIE;  //complement 
assign rif = ~RIF;  //complement 
assign jrb =  ria & rib & ric & rid & rie & rif  ; 
assign JRB = ~jrb;  //complement  
assign qtw = ~QTW;  //complement 
assign qkl = ~QKL;  //complement 
assign qkm = ~QKM;  //complement 
assign qkn = ~QKN;  //complement 
assign ria = ~RIA;  //complement 
assign rib = ~RIB;  //complement 
assign ric = ~RIC;  //complement 
assign lbb = ~LBB;  //complement 
assign aeh = ~AEH;  //complement 
assign aei = ~AEI;  //complement 
assign aej = ~AEJ;  //complement 
assign aek = ~AEK;  //complement 
assign ACJ = ~acj;  //complement 
assign ADB = ~adb;  //complement 
assign ADJ = ~adj;  //complement 
assign BHA =  aeh & ASH  |  asi & AEI  |  ASI & aei  |  aaj & AEJ  |  AAJ & aej  |  ash & AEH  ;
assign bha = ~BHA;  //complement 
assign ael = ~AEL;  //complement 
assign aem = ~AEM;  //complement 
assign aen = ~AEN;  //complement 
assign aeo = ~AEO;  //complement 
assign cda = ~CDA;  //complement 
assign BHC =  aen & ASN  |  asn & AEN  |  ASO & aeo  |  aso & AEO  |  ASP & aep  |  asp & AEP  ;
assign bhc = ~BHC;  //complement 
assign aep = ~AEP;  //complement 
assign afa = ~AFA;  //complement 
assign afb = ~AFB;  //complement 
assign afc = ~AFC;  //complement 
assign cdb = ~CDB;  //complement 
assign BHE =  afd & ATD  |  atd & AFD  |  ATE & afe  |  ate & AFE  |  ATF & aff  |  atf & AFF  ;
assign bhe = ~BHE;  //complement 
assign afd = ~AFD;  //complement 
assign afe = ~AFE;  //complement 
assign aff = ~AFF;  //complement 
assign afg = ~AFG;  //complement 
assign afh = ~AFH;  //complement 
assign afi = ~AFI;  //complement 
assign afj = ~AFJ;  //complement 
assign afk = ~AFK;  //complement 
assign JOA =  cca & ccb  ; 
assign joa = ~JOA;  //complement 
assign JOB =  cda & cdb  ; 
assign job = ~JOB;  //complement 
assign JOC =  cea & ceb  ; 
assign joc = ~JOC;  //complement 
assign BHG =  ABJ & afj  |  abj & AFJ  |  ATK & afk  |  atk & AFK  |  ATL & afl  |  atl & AFL  ;
assign bhg = ~BHG;  //complement 
assign afl = ~AFL;  //complement 
assign afm = ~AFM;  //complement 
assign afn = ~AFN;  //complement 
assign afo = ~AFO;  //complement 
assign GBJ = ~gbj;  //complement 
assign GBI = ~gbi;  //complement 
assign FBB = EBK & ebl ; 
assign fbb = ~FBB ; //complement 
assign FBH = EBK & ZZI ; 
assign fbh = ~FBH ;  //complement 
assign FBG = EBJ; 
assign fbg = ~FBG;  //complement 
assign GBP = ~gbp;  //complement 
assign GBE = ~gbe;  //complement 
assign FAJ =  eal & eak & EAJ  ; 
assign faj = ~FAJ;  //complement 
assign qkg = ~QKG;  //complement 
assign qkh = ~QKH;  //complement 
assign JCZ = QKJ & ZZI ; 
assign jcz = ~JCZ ; //complement 
assign JCY = QKJ & ZZI ; 
assign jcy = ~JCY ;  //complement 
assign jco = qkj & rbd ; 
assign JCO = ~jco ;  //complement 
assign jcp = qkj & ZZI; 
assign JCP = ~jcp; 
assign JLB = QLE & lba ; 
assign jlb = ~JLB ; //complement 
assign JLA = QLE & ZZI ; 
assign jla = ~JLA ;  //complement 
assign qkf = ~QKF;  //complement 
assign hei = ~HEI;  //complement 
assign hej = ~HEJ;  //complement 
assign BHB =  ASK & aek  |  ask & AEK  |  ASL & ael  |  asl & AEL  |  ASM & aem  |  asm & AEM  ;
assign bhb = ~BHB;  //complement 
assign aab = ~AAB;  //complement 
assign WAB =  ZZO & ZZI & qxa  |  AAB & ZZI & QXA  ; 
assign wab = ~WAB;  //complement 
assign WAJ =  BAJ & ZZI & qxa  |  AAJ & ZZI & QXA  ; 
assign waj = ~WAJ;  //complement 
assign oab = ~OAB;  //complement 
assign oaj = ~OAJ;  //complement 
assign BHD =  ATA & afa  |  ata & AFA  |  ABB & afb  |  abb & AFB  |  ATC & afc  |  atc & AFC  ;
assign bhd = ~BHD;  //complement 
assign asj = ~ASJ;  //complement 
assign aaj = ~AAJ;  //complement 
assign tda = QXF; 
assign TDA = ~tda; //complement 
assign tdb = QXF; 
assign TDB = ~tdb;  //complement 
assign TDC = qxf; 
assign tdc = ~TDC;  //complement 
assign TDD = qxf; 
assign tdd = ~TDD;  //complement 
assign wcb = aab; 
assign WCB = ~wcb; //complement 
assign wcj = aaj; 
assign WCJ = ~wcj;  //complement 
assign wdb = abb; 
assign WDB = ~wdb;  //complement 
assign wdj = abj; 
assign WDJ = ~wdj;  //complement 
assign BHF =  ATG & afg  |  atg & AFG  |  ATH & afh  |  ath & AFH  |  ATI & afi  |  ati & AFI  ;
assign bhf = ~BHF;  //complement 
assign atb = ~ATB;  //complement 
assign abb = ~ABB;  //complement 
assign dab = ~DAB;  //complement 
assign daj = ~DAJ;  //complement 
assign dbb = ~DBB;  //complement 
assign dbj = ~DBJ;  //complement 
assign ORB = ~orb;  //complement 
assign edb = ~EDB;  //complement 
assign edj = ~EDJ;  //complement 
assign BHH =  ATM & afm  |  atm & AFM  |  ATN & afn  |  atn & AFN  |  ATO & afo  |  ato & AFO  ;
assign bhh = ~BHH;  //complement 
assign atj = ~ATJ;  //complement 
assign abj = ~ABJ;  //complement 
assign WBB =  BBB & ZZI & qxb  |  ABB & ZZI & QXB  ; 
assign wbb = ~WBB;  //complement 
assign WBJ =  BBJ & ZZI & qxb  |  ABJ & ZZI & QXB  ; 
assign wbj = ~WBJ;  //complement 
assign obb = ~OBB;  //complement 
assign obj = ~OBJ;  //complement 
assign EAB = ~eab;  //complement 
assign EAJ = ~eaj;  //complement 
assign EBJ = ~ebj;  //complement 
assign ECJ = ~ecj;  //complement 
assign nab = ~NAB;  //complement 
assign nbb = ~NBB;  //complement 
assign ncb = ~NCB;  //complement 
assign qxe = ~QXE;  //complement 
assign qxf = ~QXF;  //complement 
assign OCB = ~ocb;  //complement 
assign OCJ = ~ocj;  //complement 
assign ODB = ~odb;  //complement 
assign ODJ = ~odj;  //complement 
assign qkx = ~QKX;  //complement 
assign JSE =  QQI & NBA & NBB & NBC & NBD  ; 
assign jse = ~JSE;  //complement  
assign JSD =  QQI & NBA & NBB & NBC  ; 
assign jsd = ~JSD;  //complement 
assign qkj = ~QKJ;  //complement 
assign oje = ~OJE;  //complement 
assign qga = ~QGA;  //complement 
assign JBB =  QGE  |  qgd & HEI  |  QGD & HEJ  |  qkf & QKG  |  QKF & QKH  |  QKX  ;
assign jbb = ~JBB;  //complement 
assign rfb = ~RFB;  //complement 
assign ojb = ~OJB;  //complement 
assign JBC = RGA & ~cab & ~caa  |  RGB & ~cab & caa  |  RGC & cab & ~caa  |  RGD & cab & caa; 
assign jbc = ~JBC;  //complement 
assign JBD = RGA & ~cab & ~caa  |         RGB & ~cab & caa  |  RGC & cab & ~caa  |  RGD & cab & caa ; 
assign jbd = ~JBD;  //complement 
assign oeb = ~OEB;  //complement 
assign caa = ~CAA;  //complement 
assign cab = ~CAB;  //complement 
assign cac = ~CAC;  //complement 
assign kab = ~KAB;  //complement 
assign rfa = ~RFA;  //complement 
assign oja = ~OJA;  //complement 
assign rga = ~RGA;  //complement 
assign rgb = ~RGB;  //complement 
assign rgc = ~RGC;  //complement 
assign rgd = ~RGD;  //complement 
assign lab = ~LAB;  //complement 
assign pac = ~PAC;  //complement 
assign pcc = ~PCC;  //complement 
assign pec = ~PEC;  //complement 
assign JGC =  QVB & PCB  ; 
assign jgc = ~JGC;  //complement  
assign JGK =  QVD & PCI & PCJ  ; 
assign jgk = ~JGK;  //complement 
assign JDK =  QWD & BCI & BCJ  ; 
assign jdk = ~JDK;  //complement 
assign jfj =  gbc & gbd & gbe & gbf & gbg & gae  ; 
assign JFJ = ~jfj;  //complement  
assign pak = ~PAK;  //complement 
assign pck = ~PCK;  //complement 
assign pek = ~PEK;  //complement 
assign qub = ~QUB;  //complement 
assign quc = ~QUC;  //complement 
assign que = ~QUE;  //complement 
assign QVB = ~qvb;  //complement 
assign bak = ~BAK;  //complement 
assign bck = ~BCK;  //complement 
assign bek = ~BEK;  //complement 
assign qpa = ~QPA;  //complement 
assign qpb = ~QPB;  //complement 
assign qpc = ~QPC;  //complement 
assign qpd = ~QPD;  //complement 
assign pbc = ~PBC;  //complement 
assign pdc = ~PDC;  //complement 
assign pfc = ~PFC;  //complement 
assign qua = ~QUA;  //complement 
assign quf = ~QUF;  //complement 
assign bbc = ~BBC;  //complement 
assign bdc = ~BDC;  //complement 
assign bfc = ~BFC;  //complement 
assign qud = ~QUD;  //complement 
assign pbk = ~PBK;  //complement 
assign pdk = ~PDK;  //complement 
assign pfk = ~PFK;  //complement 
assign JHK =  QVG & QVI & PDI & PDJ  ; 
assign jhk = ~JHK;  //complement  
assign JHC =  QVF & PDA & PDB  ; 
assign jhc = ~JHC;  //complement 
assign bbk = ~BBK;  //complement 
assign bdk = ~BDK;  //complement 
assign bfk = ~BFK;  //complement 
assign JEC =  QWF & BDA & BDB  ; 
assign jec = ~JEC;  //complement 
assign JEK =  QWH & BDI & BDJ  ; 
assign jek = ~JEK;  //complement 
assign rma = ~RMA;  //complement 
assign rmc = ~RMC;  //complement 
assign rmd = ~RMD;  //complement 
assign rnm = ~RNM;  //complement 
assign rnn = ~RNN;  //complement 
assign rno = ~RNO;  //complement 
assign rnp = ~RNP;  //complement 
assign rna = ~RNA;  //complement 
assign rnk = ~RNK;  //complement 
assign rmn = ~RMN;  //complement 
assign rmg = ~RMG;  //complement 
assign rmh = ~RMH;  //complement 
assign rmi = ~RMI;  //complement 
assign rmj = ~RMJ;  //complement 
assign jrc =  rna & rnb & rnc & rnd  ; 
assign JRC = ~jrc;  //complement  
assign JKB =  QLL & QLM  ; 
assign jkb = ~JKB;  //complement 
assign rmk = ~RMK;  //complement 
assign rme = ~RME;  //complement 
assign rml = ~RML;  //complement 
assign rmm = ~RMM;  //complement 
assign rmo = ~RMO;  //complement 
assign rmp = ~RMP;  //complement 
assign rnb = ~RNB;  //complement 
assign rnc = ~RNC;  //complement 
assign rnd = ~RND;  //complement 
assign rnl = ~RNL;  //complement 
assign rmr = ~RMR;  //complement 
assign rmf = ~RMF;  //complement 
assign rmq = ~RMQ;  //complement 
assign rms = ~RMS;  //complement 
assign rmt = ~RMT;  //complement 
assign rmu = ~RMU;  //complement 
assign rmb = ~RMB;  //complement 
assign lbc = ~LBC;  //complement 
assign agh = ~AGH;  //complement 
assign agi = ~AGI;  //complement 
assign agj = ~AGJ;  //complement 
assign agk = ~AGK;  //complement 
assign ACK = ~ack;  //complement 
assign ADC = ~adc;  //complement 
assign ADK = ~adk;  //complement 
assign BIA =  agh & ASH  |  asi & AGI  |  ASI & agi  |  asj & AGJ  |  ASJ & agj  |  ash & AGH  ;
assign bia = ~BIA;  //complement 
assign agl = ~AGL;  //complement 
assign agm = ~AGM;  //complement 
assign agn = ~AGN;  //complement 
assign ago = ~AGO;  //complement 
assign cea = ~CEA;  //complement 
assign BIC =  agn & ASN  |  asn & AGN  |  ASO & ago  |  aso & AGO  |  ASP & agp  |  asp & AGP  ;
assign bic = ~BIC;  //complement 
assign agp = ~AGP;  //complement 
assign aha = ~AHA;  //complement 
assign ahb = ~AHB;  //complement 
assign ahc = ~AHC;  //complement 
assign ceb = ~CEB;  //complement 
assign BIE =  ahd & ATD  |  atd & AHD  |  ATE & ahe  |  ate & AHE  |  ATF & ahf  |  atf & AHF  ;
assign bie = ~BIE;  //complement 
assign ahd = ~AHD;  //complement 
assign ahe = ~AHE;  //complement 
assign ahf = ~AHF;  //complement 
assign ahg = ~AHG;  //complement 
assign ahh = ~AHH;  //complement 
assign ahi = ~AHI;  //complement 
assign ahj = ~AHJ;  //complement 
assign ahk = ~AHK;  //complement 
assign GAC = ~gac;  //complement 
assign GCK = ~gck;  //complement 
assign gae = ~GAE;  //complement 
assign BIG =  ahj & ATJ  |  atj & AHJ  |  ABK & ahk  |  abk & AHK  |  ATL & ahl  |  atl & AHL  ;
assign big = ~BIG;  //complement 
assign ahl = ~AHL;  //complement 
assign ahm = ~AHM;  //complement 
assign ahn = ~AHN;  //complement 
assign aho = ~AHO;  //complement 
assign GAG = ~gag;  //complement 
assign GCH = ~gch;  //complement 
assign GAL = ~gal;  //complement 
assign GAN = ~gan;  //complement 
assign FAD =  eap & eao & ean & eam  ; 
assign fad = ~FAD;  //complement  
assign FAA =  eap & eao & ean & eam  ; 
assign faa = ~FAA;  //complement 
assign GBC = ~gbc;  //complement 
assign GBD = ~gbd;  //complement 
assign GBG = ~gbg;  //complement 
assign GBA = ~gba;  //complement 
assign FAC =  ebp & eao & ean  ; 
assign fac = ~FAC;  //complement 
assign FAK =  eal & EAK & eaj  ; 
assign fak = ~FAK;  //complement 
assign FBC =  EBL & ebk & eaj  ; 
assign fbc = ~FBC;  //complement 
assign GBK = ~gbk;  //complement 
assign GBF = ~gbf;  //complement 
assign qkb = ~QKB;  //complement 
assign hfm = ~HFM;  //complement 
assign hfn = ~HFN;  //complement 
assign qka = ~QKA;  //complement 
assign JLC =  QLE & lba & lbb  ; 
assign jlc = ~JLC;  //complement 
assign maa = ~MAA;  //complement 
assign mab = ~MAB;  //complement 
assign mac = ~MAC;  //complement 
assign JAA =  QAA & GAN & gab  ; 
assign jaa = ~JAA;  //complement 
assign JCI =  gal & GAN  ; 
assign jci = ~JCI;  //complement 
assign BIB =  AAK & agk  |  aak & AGK  |  ASL & agl  |  asl & AGL  |  ASM & agm  |  asm & AGM  ;
assign bib = ~BIB;  //complement 
assign aac = ~AAC;  //complement 
assign oha = ~OHA;  //complement 
assign WAC =  ZZO & ZZI & qxa  |  AAC & ZZI & QXA  ; 
assign wac = ~WAC;  //complement 
assign WAK =  BAK & ZZI & qxa  |  AAK & ZZI & QXA  ; 
assign wak = ~WAK;  //complement 
assign oac = ~OAC;  //complement 
assign oak = ~OAK;  //complement 
assign BID =  ATA & aha  |  ata & AHA  |  ATB & ahb  |  atb & AHB  |  ABC & ahc  |  abc & AHC  ;
assign bid = ~BID;  //complement 
assign ask = ~ASK;  //complement 
assign aak = ~AAK;  //complement 
assign tca = qxe; 
assign TCA = ~tca; //complement 
assign tcb = qxe; 
assign TCB = ~tcb;  //complement 
assign TCC = QXE; 
assign tcc = ~TCC;  //complement 
assign TCD = QXE; 
assign tcd = ~TCD;  //complement 
assign wcc = aac; 
assign WCC = ~wcc; //complement 
assign wck = aak; 
assign WCK = ~wck;  //complement 
assign wdc = abc; 
assign WDC = ~wdc;  //complement 
assign wdk = abk; 
assign WDK = ~wdk;  //complement 
assign BIF =  ATG & ahg  |  atg & AHG  |  ATH & ahh  |  ath & AHH  |  ATI & ahi  |  ati & AHI  ;
assign bif = ~BIF;  //complement 
assign atc = ~ATC;  //complement 
assign abc = ~ABC;  //complement 
assign dac = ~DAC;  //complement 
assign dak = ~DAK;  //complement 
assign dbc = ~DBC;  //complement 
assign dbk = ~DBK;  //complement 
assign ORC = ~orc;  //complement 
assign edc = ~EDC;  //complement 
assign qzf = ~QZF;  //complement 
assign BIH =  ATM & ahm  |  atm & AHM  |  ATN & ahn  |  atn & AHN  |  ATO & aho  |  ato & AHO  ;
assign bih = ~BIH;  //complement 
assign atk = ~ATK;  //complement 
assign abk = ~ABK;  //complement 
assign WBC =  BBC & ZZI & qxb  |  ABC & ZZI & QXB  ; 
assign wbc = ~WBC;  //complement 
assign WBK =  BBK & ZZI & qxb  |  ABK & ZZI & QXB  ; 
assign wbk = ~WBK;  //complement 
assign obc = ~OBC;  //complement 
assign obk = ~OBK;  //complement 
assign EBK = ~ebk;  //complement 
assign EAK = ~eak;  //complement 
assign EAC = ~eac;  //complement 
assign ECK = ~eck;  //complement 
assign nac = ~NAC;  //complement 
assign nbc = ~NBC;  //complement 
assign jac = gac; 
assign JAC = ~jac;  //complement 
assign OCC = ~occ;  //complement 
assign OCK = ~ock;  //complement 
assign ODC = ~odc;  //complement 
assign ODK = ~odk;  //complement 
assign JNC = QNG & MAC ; 
assign jnc = ~JNC ; //complement 
assign JND = QNG & ZZI ; 
assign jnd = ~JND ;  //complement 
assign jne = qng & rqc ; 
assign JNE = ~jne ;  //complement 
assign JAN =  QCZ & HFN & QGA  |  QCZ & HFN & QGB  ; 
assign jan = ~JAN;  //complement 
assign JBE =  HFM & qga & qgb  |  HFN & QGA  |  HFN & QGB  ; 
assign jbe = ~JBE; //complement 
assign qgb = ~QGB;  //complement 
assign qkc = ~QKC;  //complement 
assign qfa = ~QFA;  //complement 
assign RMV = ~rmv;  //complement 
assign rag = ~RAG;  //complement 
assign oka = ~OKA;  //complement 
assign oec = ~OEC;  //complement 
assign edk = ~EDK;  //complement 
assign kac = ~KAC;  //complement 
assign kae = ~KAE;  //complement 
assign qkd = ~QKD;  //complement 
assign qke = ~QKE;  //complement 
assign okb = ~OKB;  //complement 
assign lac = ~LAC;  //complement 
assign pad = ~PAD;  //complement 
assign pcd = ~PCD;  //complement 
assign ped = ~PED;  //complement 
assign JGD =  QVB & PCB & PCC  ; 
assign jgd = ~JGD;  //complement  
assign JGL =  QVD & PCI & PCJ & PCK  ; 
assign jgl = ~JGL;  //complement 
assign JDB =  BEI & BEJ & BEK & BEL  ; 
assign jdb = ~JDB;  //complement  
assign JDL =  QWD & BCI & BCJ & BCK  ; 
assign jdl = ~JDL;  //complement 
assign JDD =  BFA & BFB & BFC & BFD  ; 
assign jdd = ~JDD;  //complement  
assign JDF =  BFI & BFJ & BFK & BFL  ; 
assign jdf = ~JDF;  //complement 
assign pal = ~PAL;  //complement 
assign pcl = ~PCL;  //complement 
assign pel = ~PEL;  //complement 
assign JFA =  ZZI & PEB & PEC & PED  ; 
assign jfa = ~JFA;  //complement  
assign JFC =  PEI & PEJ & PEK & PEL  ; 
assign jfc = ~JFC;  //complement 
assign bal = ~BAL;  //complement 
assign bel = ~BEL;  //complement 
assign qwb = ~QWB;  //complement 
assign qwc = ~QWC;  //complement 
assign QWI = ~qwi;  //complement 
assign QWD = ~qwd;  //complement 
assign pbd = ~PBD;  //complement 
assign pdd = ~PDD;  //complement 
assign pfd = ~PFD;  //complement 
assign tfc = qwa; 
assign TFC = ~tfc; //complement 
assign tfd = qwa; 
assign TFD = ~tfd;  //complement 
assign tfa = qwa; 
assign TFA = ~tfa;  //complement 
assign tfb = qwa; 
assign TFB = ~tfb;  //complement 
assign bbd = ~BBD;  //complement 
assign bfd = ~BFD;  //complement 
assign qwa = ~QWA;  //complement 
assign qwj = ~QWJ;  //complement 
assign pbl = ~PBL;  //complement 
assign pdl = ~PDL;  //complement 
assign pfl = ~PFL;  //complement 
assign JHL =  QVG & QVI & PDI & PDJ & PDK  ; 
assign jhl = ~JHL;  //complement  
assign JHD =  QVF & PDA & PDB & PDC  ; 
assign jhd = ~JHD;  //complement 
assign bbl = ~BBL;  //complement 
assign bfl = ~BFL;  //complement 
assign JED =  QWF & BDA & BDB & BDC  ; 
assign jed = ~JED;  //complement  
assign JEL =  QWH & BDI & BDJ & BDK  ; 
assign jel = ~JEL;  //complement 
assign qll = ~QLL;  //complement 
assign rkb = ~RKB;  //complement 
assign rkc = ~RKC;  //complement 
assign rkd = ~RKD;  //complement 
assign rlb = ~RLB;  //complement 
assign rld = ~RLD;  //complement 
assign rla = ~RLA;  //complement 
assign qlm = ~QLM;  //complement 
assign qla = ~QLA;  //complement 
assign qlb = ~QLB;  //complement 
assign qlc = ~QLC;  //complement 
assign rlc = ~RLC;  //complement 
assign jka =  qlf & rka & rkb & rkc & rkd  ; 
assign JKA = ~jka;  //complement  
assign qlf = ~QLF;  //complement 
assign qlg = ~QLG;  //complement 
assign qld = ~QLD;  //complement 
assign qln = ~QLN;  //complement 
assign qlo = ~QLO;  //complement 
assign qli = ~QLI;  //complement 
assign qlk = ~QLK;  //complement 
assign jqa =  qln & qqm & qqk  ; 
assign JQA = ~jqa;  //complement 
assign jjg =  ZZI & ZZI & qln  ; 
assign JJG = ~jjg;  //complement 
assign lbd = ~LBD;  //complement 
assign aih = ~AIH;  //complement 
assign aii = ~AII;  //complement 
assign aij = ~AIJ;  //complement 
assign aik = ~AIK;  //complement 
assign ACL = ~acl;  //complement 
assign ADD = ~add;  //complement 
assign ADL = ~adl;  //complement 
assign BJA =  aih & ASH  |  asi & AII  |  ASI & aii  |  asj & AIJ  |  ASJ & aij  |  ash & AIH  ;
assign bja = ~BJA;  //complement 
assign ail = ~AIL;  //complement 
assign aim = ~AIM;  //complement 
assign ain = ~AIN;  //complement 
assign aio = ~AIO;  //complement 
assign cfa = ~CFA;  //complement 
assign BJC =  ain & ASN  |  asn & AIN  |  ASO & aio  |  aso & AIO  |  ASP & aip  |  asp & AIP  ;
assign bjc = ~BJC;  //complement 
assign aip = ~AIP;  //complement 
assign aja = ~AJA;  //complement 
assign ajb = ~AJB;  //complement 
assign ajc = ~AJC;  //complement 
assign cfb = ~CFB;  //complement 
assign BJE =  ABD & ajd  |  abd & AJD  |  ATE & aje  |  ate & AJE  |  ATF & ajf  |  atf & AJF  ;
assign bje = ~BJE;  //complement 
assign ajd = ~AJD;  //complement 
assign aje = ~AJE;  //complement 
assign ajf = ~AJF;  //complement 
assign ajg = ~AJG;  //complement 
assign ajh = ~AJH;  //complement 
assign aji = ~AJI;  //complement 
assign ajj = ~AJJ;  //complement 
assign ajk = ~AJK;  //complement 
assign GCL = ~gcl;  //complement 
assign GAH = ~gah;  //complement 
assign GAF = ~gaf;  //complement 
assign BJG =  ajj & ATJ  |  atj & AJJ  |  ATK & ajk  |  atk & AJK  |  ABL & ajl  |  abl & AJL  ;
assign bjg = ~BJG;  //complement 
assign ajl = ~AJL;  //complement 
assign ajm = ~AJM;  //complement 
assign ajn = ~AJN;  //complement 
assign ajo = ~AJO;  //complement 
assign jfy =  rbd & rld  ; 
assign JFY = ~jfy;  //complement 
assign jfx =  gaf  ; 
assign JFX = ~jfx;  //complement 
assign GCA = ~gca;  //complement 
assign GCB = ~gcb;  //complement 
assign FAG =  eap & EAO & EAN & eam  ; 
assign fag = ~FAG;  //complement  
assign FBD =  EBL & EBK  ; 
assign fbd = ~FBD;  //complement 
assign qlp = ~QLP;  //complement 
assign qlq = ~QLQ;  //complement 
assign GCC = ~gcc;  //complement 
assign GCD = ~gcd;  //complement 
assign FBE =  EBL  ; 
assign fbe = ~FBE;  //complement  
assign FAL =  eal & EAK & EAJ  ; 
assign fal = ~FAL;  //complement 
assign rka = ~RKA;  //complement 
assign qlj = ~QLJ;  //complement 
assign qrb = ~QRB;  //complement 
assign qrc = ~QRC;  //complement 
assign qrd = ~QRD;  //complement 
assign qre = ~QRE;  //complement 
assign JAG =  QAD  ; 
assign jag = ~JAG;  //complement 
assign jrd =  qia & qib & qic  ; 
assign JRD = ~jrd;  //complement 
assign jjk =  rlc & qic  ; 
assign JJK = ~jjk;  //complement 
assign JLD =  QLE & lba & lbb & lbc  ; 
assign jld = ~JLD;  //complement  
assign QNA = ~qna;  //complement 
assign QNE = ~qne;  //complement 
assign jra =  qia & qib & qic & qid  ; 
assign JRA = ~jra;  //complement  
assign tld =  qma & qne  ; 
assign TLD = ~tld;  //complement 
assign BJB =  ASK & aik  |  ask & AIK  |  AAL & ail  |  aal & AIL  |  ASM & aim  |  asm & AIM  ;
assign bjb = ~BJB;  //complement 
assign aad = ~AAD;  //complement 
assign ohb = ~OHB;  //complement 
assign WAD =  ZZO & ZZI & qxa  |  AAD & ZZI & QXA  ; 
assign wad = ~WAD;  //complement 
assign WAL =  BAL & ZZI & qxa  |  AAL & ZZI & QXA  ; 
assign wal = ~WAL;  //complement 
assign oad = ~OAD;  //complement 
assign oal = ~OAL;  //complement 
assign BJD =  ATA & aja  |  ata & AJA  |  ATB & ajb  |  atb & AJB  |  ATC & ajc  |  atc & AJC  ;
assign bjd = ~BJD;  //complement 
assign asl = ~ASL;  //complement 
assign aal = ~AAL;  //complement 
assign taa = rjl; 
assign TAA = ~taa; //complement 
assign tab = rjl; 
assign TAB = ~tab;  //complement 
assign TAC = RJL; 
assign tac = ~TAC;  //complement 
assign TAD = RJL; 
assign tad = ~TAD;  //complement 
assign wcd = aad; 
assign WCD = ~wcd; //complement 
assign wcl = aal; 
assign WCL = ~wcl;  //complement 
assign wdd = abd; 
assign WDD = ~wdd;  //complement 
assign wdl = abl; 
assign WDL = ~wdl;  //complement 
assign BJF =  ATG & ajg  |  atg & AJG  |  ATH & ajh  |  ath & AJH  |  ATI & aji  |  ati & AJI  ;
assign bjf = ~BJF;  //complement 
assign atd = ~ATD;  //complement 
assign abd = ~ABD;  //complement 
assign dad = ~DAD;  //complement 
assign dal = ~DAL;  //complement 
assign dbd = ~DBD;  //complement 
assign dbl = ~DBL;  //complement 
assign ORD = ~ord;  //complement 
assign edd = ~EDD;  //complement 
assign edl = ~EDL;  //complement 
assign rjl = ~RJL;  //complement 
assign BJH =  ATM & ajm  |  atm & AJM  |  ATN & ajn  |  atn & AJN  |  ATO & ajo  |  ato & AJO  ;
assign bjh = ~BJH;  //complement 
assign atl = ~ATL;  //complement 
assign abl = ~ABL;  //complement 
assign WBD =  BBD & ZZI & qxb  |  ABD & ZZI & QXB  ; 
assign wbd = ~WBD;  //complement 
assign WBL =  BBL & ZZI & qxb  |  ABL & ZZI & QXB  ; 
assign wbl = ~WBL;  //complement 
assign obd = ~OBD;  //complement 
assign obl = ~OBL;  //complement 
assign EBL = ~ebl;  //complement 
assign EAL = ~eal;  //complement 
assign EAD = ~ead;  //complement 
assign ECL = ~ecl;  //complement 
assign nad = ~NAD;  //complement 
assign nbd = ~NBD;  //complement 
assign qfb = ~QFB;  //complement 
assign olf = ~OLF;  //complement 
assign OCD = ~ocd;  //complement 
assign OCL = ~ocl;  //complement 
assign ODD = ~odd;  //complement 
assign ODL = ~odl;  //complement 
assign qni = ~QNI;  //complement 
assign qnm = ~QNM;  //complement 
assign qnq = ~QNQ;  //complement 
assign qnu = ~QNU;  //complement 
assign qra = ~QRA;  //complement 
assign ojc = ~OJC;  //complement 
assign oma = ~OMA;  //complement 
assign omb = ~OMB;  //complement 
assign jjc =  rjc  ; 
assign JJC = ~jjc;  //complement 
assign jjb =  rae & raf & rjk  ; 
assign JJB = ~jjb;  //complement 
assign jkc =  qlg & qli & rjk  ; 
assign JKC = ~jkc;  //complement 
assign qlr = ~QLR;  //complement 
assign qls = ~QLS;  //complement 
assign rjc = ~RJC;  //complement 
assign rix = ~RIX;  //complement 
assign ojd = ~OJD;  //complement 
assign oed = ~OED;  //complement 
assign OEI = ~oei;  //complement 
assign kad = ~KAD;  //complement 
assign QIB = ~qib;  //complement 
assign QIC = ~qic;  //complement 
assign QID = ~qid;  //complement 
assign otc = ~OTC;  //complement 
assign QIA = ~qia;  //complement 
assign lad = ~LAD;  //complement 
assign pae = ~PAE;  //complement 
assign pce = ~PCE;  //complement 
assign pee = ~PEE;  //complement 
assign JGE =  QVC  ; 
assign jge = ~JGE;  //complement  
assign JGM =  QVE  ; 
assign jgm = ~JGM;  //complement 
assign JDM =  QWE  ; 
assign jdm = ~JDM;  //complement 
assign pam = ~PAM;  //complement 
assign pcm = ~PCM;  //complement 
assign pem = ~PEM;  //complement 
assign QVC = ~qvc;  //complement 
assign QVD = ~qvd;  //complement 
assign bam = ~BAM;  //complement 
assign bcm = ~BCM;  //complement 
assign bem = ~BEM;  //complement 
assign QWH = ~qwh;  //complement 
assign pbe = ~PBE;  //complement 
assign pde = ~PDE;  //complement 
assign pfe = ~PFE;  //complement 
assign bbe = ~BBE;  //complement 
assign bde = ~BDE;  //complement 
assign bfe = ~BFE;  //complement 
assign pbm = ~PBM;  //complement 
assign pdm = ~PDM;  //complement 
assign JHM =  QVG & QVJ  ; 
assign jhm = ~JHM;  //complement  
assign JHE =  QVF & QVH  ; 
assign jhe = ~JHE;  //complement 
assign bbm = ~BBM;  //complement 
assign bdm = ~BDM;  //complement 
assign JEE =  QWG  ; 
assign jee = ~JEE;  //complement 
assign JEM =  QWI & QWH  ; 
assign jem = ~JEM;  //complement 
assign jcx = rbf & qcz ; 
assign JCX = ~jcx ; //complement 
assign rbx = ~RBX;  //complement 
assign jck =  gbm & gbn & gbp  ; 
assign JCK = ~jck;  //complement  
assign jcl =  gbm & gbn & gbo & gbp  ; 
assign JCL = ~jcl;  //complement 
assign QNJ = ~qnj;  //complement 
assign QNN = ~qnn;  //complement 
assign QNR = ~qnr;  //complement 
assign QNV = ~qnv;  //complement 
assign qmk = ~QMK;  //complement 
assign qml = ~QML;  //complement 
assign lbe = ~LBE;  //complement 
assign akh = ~AKH;  //complement 
assign aki = ~AKI;  //complement 
assign akj = ~AKJ;  //complement 
assign akk = ~AKK;  //complement 
assign ACM = ~acm;  //complement 
assign ADE = ~ade;  //complement 
assign ADM = ~adm;  //complement 
assign BKA =  akh & ASH  |  asi & AKI  |  ASI & aki  |  asj & AKJ  |  ASJ & akj  |  ash & AKH  ;
assign bka = ~BKA;  //complement 
assign akl = ~AKL;  //complement 
assign akm = ~AKM;  //complement 
assign akn = ~AKN;  //complement 
assign ako = ~AKO;  //complement 
assign cga = ~CGA;  //complement 
assign BKC =  akn & ASN  |  asn & AKN  |  ASO & ako  |  aso & AKO  |  ASP & akp  |  asp & AKP  ;
assign bkc = ~BKC;  //complement 
assign akp = ~AKP;  //complement 
assign ala = ~ALA;  //complement 
assign alb = ~ALB;  //complement 
assign alc = ~ALC;  //complement 
assign cgb = ~CGB;  //complement 
assign BKE =  ald & ATD  |  atd & ALD  |  ABE & ale  |  abe & ALE  |  ATF & alf  |  atf & ALF  ;
assign bke = ~BKE;  //complement 
assign ald = ~ALD;  //complement 
assign ale = ~ALE;  //complement 
assign alf = ~ALF;  //complement 
assign alg = ~ALG;  //complement 
assign alh = ~ALH;  //complement 
assign ali = ~ALI;  //complement 
assign alj = ~ALJ;  //complement 
assign alk = ~ALK;  //complement 
assign GCM = ~gcm;  //complement 
assign GCJ = ~gcj;  //complement 
assign GCN = ~gcn;  //complement 
assign BKG =  alj & ATJ  |  atj & ALJ  |  ATK & alk  |  atk & ALK  |  ATL & all  |  atl & ALL  ;
assign bkg = ~BKG;  //complement 
assign all = ~ALL;  //complement 
assign alm = ~ALM;  //complement 
assign aln = ~ALN;  //complement 
assign alo = ~ALO;  //complement 
assign rbb = ~RBB;  //complement 
assign rbc = ~RBC;  //complement 
assign rbd = ~RBD;  //complement 
assign rbe = ~RBE;  //complement 
assign GBN = ~gbn;  //complement 
assign GBM = ~gbm;  //complement 
assign FAE =  eap & EAO & ean & eam  ; 
assign fae = ~FAE;  //complement  
assign FAB =  ebp & eao & ean & EAM  ; 
assign fab = ~FAB;  //complement 
assign jfh = gbm & gbn ; 
assign JFH = ~jfh ; //complement 
assign jcj = gbm & gbo ; 
assign JCJ = ~jcj ;  //complement 
assign JOX = qqs & RBD ; 
assign jox = ~JOX ;  //complement 
assign JCM =  QKS & RAE  ; 
assign jcm = ~JCM;  //complement  
assign JCW =  qks & RAE & heo & hep  ; 
assign jcw = ~JCW;  //complement 
assign GAP = ~gap;  //complement 
assign GBO = ~gbo;  //complement 
assign jcg =  rae & raf & qkj  |  ZZI & ZZI & QCY  ; 
assign JCG = ~jcg;  //complement 
assign jbg =  ZZI & ZZI & qkj  |  ZZI & ZZI & QCY  ; 
assign JBG = ~jbg;  //complement 
assign qle = ~QLE;  //complement 
assign raf = ~RAF;  //complement 
assign qko = ~QKO;  //complement 
assign qks = ~QKS;  //complement 
assign jcc =  rja & rat  ; 
assign JCC = ~jcc;  //complement 
assign jre =  qlp & qsi  ; 
assign JRE = ~jre;  //complement 
assign jol =  rae & rbc  ; 
assign JOL = ~jol;  //complement 
assign JLE =  QLE & lba & lbb & lbc & lbd  ; 
assign jle = ~JLE;  //complement  
assign rab = ~RAB;  //complement 
assign rac = ~RAC;  //complement 
assign rad = ~RAD;  //complement 
assign rae = ~RAE;  //complement 
assign qcx = ~QCX;  //complement 
assign qcz = ~QCZ;  //complement 
assign qcy = ~QCY;  //complement 
assign BKB =  ASK & akk  |  ask & AKK  |  ASL & akl  |  asl & AKL  |  AAM & akm  |  aam & AKM  ;
assign bkb = ~BKB;  //complement 
assign aae = ~AAE;  //complement 
assign ohc = ~OHC;  //complement 
assign WAE =  ZZO & ZZI & qxa  |  AAE & ZZI & QXA  ; 
assign wae = ~WAE;  //complement 
assign WAM =  BAM & ZZI & qxa  |  AAM & ZZI & QXA  ; 
assign wam = ~WAM;  //complement 
assign oae = ~OAE;  //complement 
assign oam = ~OAM;  //complement 
assign BKD =  ATA & ala  |  ata & ALA  |  ATB & alb  |  atb & ALB  |  ATC & alc  |  atc & ALC  ;
assign bkd = ~BKD;  //complement 
assign asm = ~ASM;  //complement 
assign aam = ~AAM;  //complement 
assign qxa = ~QXA;  //complement 
assign qxb = ~QXB;  //complement 
assign wce = aae; 
assign WCE = ~wce; //complement 
assign wcm = aam; 
assign WCM = ~wcm;  //complement 
assign wde = abe; 
assign WDE = ~wde;  //complement 
assign wdm = abm; 
assign WDM = ~wdm;  //complement 
assign BKF =  ATG & alg  |  atg & ALG  |  ATH & alh  |  ath & ALH  |  ATI & ali  |  ati & ALI  ;
assign bkf = ~BKF;  //complement 
assign ate = ~ATE;  //complement 
assign abe = ~ABE;  //complement 
assign dae = ~DAE;  //complement 
assign dam = ~DAM;  //complement 
assign dbe = ~DBE;  //complement 
assign dbm = ~DBM;  //complement 
assign ORE = ~ore;  //complement 
assign ede = ~EDE;  //complement 
assign edm = ~EDM;  //complement 
assign OIG = ~oig;  //complement 
assign BKH =  ABM & alm  |  abm & ALM  |  ATN & aln  |  atn & ALN  |  ATO & alo  |  ato & ALO  ;
assign bkh = ~BKH;  //complement 
assign atm = ~ATM;  //complement 
assign abm = ~ABM;  //complement 
assign WBE =  BBE & ZZI & qxb  |  ABE & ZZI & QXB  ; 
assign wbe = ~WBE;  //complement 
assign WBM =  BBM & ZZI & qxb  |  ABM & ZZI & QXB  ; 
assign wbm = ~WBM;  //complement 
assign obe = ~OBE;  //complement 
assign obm = ~OBM;  //complement 
assign EAE = ~eae;  //complement 
assign EAM = ~eam;  //complement 
assign ECM = ~ecm;  //complement 
assign EAO = ~eao;  //complement 
assign JAO =  HEO & QCY  ; 
assign jao = ~JAO;  //complement 
assign jcb =  rba & rbb & rbx  ; 
assign JCB = ~jcb;  //complement 
assign JAP =  HEP & QCY & rbx  ; 
assign jap = ~JAP;  //complement 
assign rec = ~REC;  //complement 
assign oia = ~OIA;  //complement 
assign OCE = ~oce;  //complement 
assign OCM = ~ocm;  //complement 
assign ODE = ~ode;  //complement 
assign ODM = ~odm;  //complement 
assign jce =  gac & rax & qqp & rlx & gaf  ; 
assign JCE = ~jce;  //complement  
assign jcd =  rja & raa & rax & qqz  ; 
assign JCD = ~jcd;  //complement 
assign jca =  raa & rab & rac & rad & rag  ; 
assign JCA = ~jca;  //complement  
assign JAM =  QCZ & HFM & qga & qgb  ; 
assign jam = ~JAM;  //complement 
assign oic = ~OIC;  //complement 
assign qqz = ~QQZ;  //complement 
assign oid = ~OID;  //complement 
assign qqo = ~QQO;  //complement 
assign qci = ~QCI;  //complement 
assign qkw = ~QKW;  //complement 
assign jcu =  qqz & qkw & qky  ; 
assign JCU = ~jcu;  //complement  
assign jkd =  qmj & qnm & qnq & qnj  ; 
assign JKD = ~jkd;  //complement 
assign joo = rba & rac ; 
assign JOO = ~joo ; //complement 
assign jop = rba & rac ; 
assign JOP = ~jop ;  //complement 
assign joj = rba & rac ; 
assign JOJ = ~joj ;  //complement 
assign jok = rba & rac; 
assign JOK = ~jok; 
assign oie = ~OIE;  //complement 
assign qky = ~QKY;  //complement 
assign oee = ~OEE;  //complement 
assign qrf = ~QRF;  //complement 
assign olc = ~OLC;  //complement 
assign ota = ~OTA;  //complement 
assign QMB = ~qmb;  //complement 
assign QMC = ~qmc;  //complement 
assign QMF = ~qmf;  //complement 
assign QMG = ~qmg;  //complement 
assign OTD = ~otd;  //complement 
assign QMJ = ~qmj;  //complement 
assign OIB = ~oib;  //complement 
assign QCK = ~qck;  //complement 
assign JCR = RQB; 
assign jcr = ~JCR; //complement 
assign JCT = QTP; 
assign jct = ~JCT;  //complement 
assign jrf = rix & qsa ; 
assign JRF = ~jrf ;  //complement 
assign lae = ~LAE;  //complement 
assign paf = ~PAF;  //complement 
assign pcf = ~PCF;  //complement 
assign pef = ~PEF;  //complement 
assign JGF =  QVC & PCE  ; 
assign jgf = ~JGF;  //complement  
assign JGN =  QVE & PCM  ; 
assign jgn = ~JGN;  //complement 
assign JDN =  QWE & BCM  ; 
assign jdn = ~JDN;  //complement 
assign pan = ~PAN;  //complement 
assign pcn = ~PCN;  //complement 
assign pen = ~PEN;  //complement 
assign ban = ~BAN;  //complement 
assign bcn = ~BCN;  //complement 
assign ben = ~BEN;  //complement 
assign QWF = ~qwf;  //complement 
assign QWE = ~qwe;  //complement 
assign pbf = ~PBF;  //complement 
assign pdf = ~PDF;  //complement 
assign pff = ~PFF;  //complement 
assign bbf = ~BBF;  //complement 
assign bdf = ~BDF;  //complement 
assign bff = ~BFF;  //complement 
assign pbn = ~PBN;  //complement 
assign pdn = ~PDN;  //complement 
assign JHN =  QVG & QVJ & PDM  ; 
assign jhn = ~JHN;  //complement  
assign JHF =  QVF & QVH & PDE  ; 
assign jhf = ~JHF;  //complement 
assign bbn = ~BBN;  //complement 
assign bdn = ~BDN;  //complement 
assign JEF =  QWG & BDE  ; 
assign jef = ~JEF;  //complement 
assign JEN =  QWH & QWI & BDM  ; 
assign jen = ~JEN;  //complement 
assign hia = ~HIA;  //complement 
assign hib = ~HIB;  //complement 
assign hic = ~HIC;  //complement 
assign hka = ~HKA;  //complement 
assign hkb = ~HKB;  //complement 
assign hkc = ~HKC;  //complement 
assign JJP = QQC & QQL ; 
assign jjp = ~JJP ; //complement 
assign JJH = QQC & QQC ; 
assign jjh = ~JJH ;  //complement 
assign qqc = ~QQC;  //complement 
assign qqp = ~QQP;  //complement 
assign qqq = ~QQQ;  //complement 
assign hja = ~HJA;  //complement 
assign hjb = ~HJB;  //complement 
assign hjc = ~HJC;  //complement 
assign hla = ~HLA;  //complement 
assign hlb = ~HLB;  //complement 
assign hlc = ~HLC;  //complement 
assign hma = ~HMA;  //complement 
assign hmb = ~HMB;  //complement 
assign hmc = ~HMC;  //complement 
assign gdy = ~GDY;  //complement 
assign JLG =  LBA & lbb & lbc & lbd & lbe & lbf  ; 
assign jlg = ~JLG;  //complement  
assign jje =  qqe  ; 
assign JJE = ~jje;  //complement 
assign lbf = ~LBF;  //complement 
assign amh = ~AMH;  //complement 
assign ami = ~AMI;  //complement 
assign amj = ~AMJ;  //complement 
assign amk = ~AMK;  //complement 
assign ACN = ~acn;  //complement 
assign ADF = ~adf;  //complement 
assign ADN = ~adn;  //complement 
assign BLA =  amh & ASH  |  asi & AMI  |  ASI & ami  |  asj & AMJ  |  ASJ & amj  |  ash & AMH  ;
assign bla = ~BLA;  //complement 
assign aml = ~AML;  //complement 
assign amm = ~AMM;  //complement 
assign amn = ~AMN;  //complement 
assign amo = ~AMO;  //complement 
assign cha = ~CHA;  //complement 
assign BLC =  AAN & amn  |  aan & AMN  |  ASO & amo  |  aso & AMO  |  ASP & amp  |  asp & AMP  ;
assign blc = ~BLC;  //complement 
assign amp = ~AMP;  //complement 
assign ana = ~ANA;  //complement 
assign anb = ~ANB;  //complement 
assign anc = ~ANC;  //complement 
assign chb = ~CHB;  //complement 
assign BLE =  andd  & ATD  |  atd & ANDD   |  ATE & ane  |  ate & ANE  |  ABF & anf  |  abf & ANF  ;
assign ble = ~BLE;  //complement 
assign andd  = ~ANDD ;  //complement 
assign ane = ~ANE;  //complement 
assign anf = ~ANF;  //complement 
assign ang = ~ANG;  //complement 
assign anh = ~ANH;  //complement 
assign ani = ~ANI;  //complement 
assign anj = ~ANJ;  //complement 
assign ank = ~ANK;  //complement 
assign TGF = QBA; 
assign tgf = ~TGF; //complement 
assign TGA = QBA; 
assign tga = ~TGA;  //complement 
assign BLG =  anj & ATJ  |  atj & ANJ  |  ATK & ank  |  atk & ANK  |  ATL & anl  |  atl & ANL  ;
assign blg = ~BLG;  //complement 
assign anl = ~ANL;  //complement 
assign anm = ~ANM;  //complement 
assign ann = ~ANN;  //complement 
assign ano = ~ANO;  //complement 
assign tge = qba; 
assign TGE = ~tge; //complement 
assign tgc = qba; 
assign TGC = ~tgc;  //complement 
assign tgb = qba; 
assign TGB = ~tgb;  //complement 
assign tgd = qba; 
assign TGD = ~tgd;  //complement 
assign FAF =  ebp & EAO & ean & EAM  ; 
assign faf = ~FAF;  //complement  
assign FAH =  ebp & EAO & EAN & EAM  ; 
assign fah = ~FAH;  //complement 
assign JTB =  qqa & qlq & qtw & qqb  ; 
assign jtb = ~JTB;  //complement  
assign jjl =  qql & qtr & qqc & qqz  ; 
assign JJL = ~jjl;  //complement 
assign qqb = ~QQB;  //complement 
assign qqw = ~QQW;  //complement 
assign jcn =  qka & qkj & qkt & qta & qtx  ; 
assign JCN = ~jcn;  //complement  
assign jcf =  qqt & qqp & qkj  ; 
assign JCF = ~jcf;  //complement 
assign qqd = ~QQD;  //complement 
assign qqe = ~QQE;  //complement 
assign qqf = ~QQF;  //complement 
assign qqg = ~QQG;  //complement 
assign JQE =  QQA & qko & qqb  |  QQY & qqb & QKO  ; 
assign jqe = ~JQE;  //complement 
assign jcv = qqt & qqp ; 
assign JCV = ~jcv ; //complement 
assign jcq = qqt & ZZI ; 
assign JCQ = ~jcq ;  //complement 
assign jjd = qqd; 
assign JJD = ~jjd;  //complement 
assign JLF =  QLE & lba & lbb & lbc & lbd & lbe  ; 
assign jlf = ~JLF;  //complement  
assign JXB =  QSC & qlq & qqa  ; 
assign jxb = ~JXB;  //complement 
assign qhe = ~QHE;  //complement 
assign qhf = ~QHF;  //complement 
assign QTQ = ~qtq;  //complement 
assign QTR = ~qtr;  //complement 
assign rlx = ~RLX;  //complement 
assign BLB =  ASK & amk  |  ask & AMK  |  ASL & aml  |  asl & AML  |  ASM & amm  |  asm & AMM  ;
assign blb = ~BLB;  //complement 
assign aaf = ~AAF;  //complement 
assign ohd = ~OHD;  //complement 
assign WAF =  ZZO & ZZI & qxc  |  AAF & ZZI & QXC  ; 
assign waf = ~WAF;  //complement 
assign WAN =  BAN & ZZI & qxc  |  AAN & ZZI & QXC  ; 
assign wan = ~WAN;  //complement 
assign oaf = ~OAF;  //complement 
assign oan = ~OAN;  //complement 
assign BLD =  ATA & ana  |  ata & ANA  |  ATB & anb  |  atb & ANB  |  ATC & anc  |  atc & ANC  ;
assign bld = ~BLD;  //complement 
assign asn = ~ASN;  //complement 
assign aan = ~AAN;  //complement 
assign qxc = ~QXC;  //complement 
assign qxd = ~QXD;  //complement 
assign wcf = aaf; 
assign WCF = ~wcf; //complement 
assign wcn = aan; 
assign WCN = ~wcn;  //complement 
assign wdf = abf; 
assign WDF = ~wdf;  //complement 
assign wdn = abn; 
assign WDN = ~wdn;  //complement 
assign BLF =  ATG & ang  |  atg & ANG  |  ATH & anh  |  ath & ANH  |  ATI & ani  |  ati & ANI  ;
assign blf = ~BLF;  //complement 
assign atf = ~ATF;  //complement 
assign abf = ~ABF;  //complement 
assign daf = ~DAF;  //complement 
assign dan = ~DAN;  //complement 
assign dbf = ~DBF;  //complement 
assign dbn = ~DBN;  //complement 
assign ORF = ~orf;  //complement 
assign edf = ~EDF;  //complement 
assign edn = ~EDN;  //complement 
assign BLH =  ATM & anm  |  atm & ANM  |  ABN & ann  |  abn & ANN  |  ATO & ano  |  ato & ANO  ;
assign blh = ~BLH;  //complement 
assign atn = ~ATN;  //complement 
assign abn = ~ABN;  //complement 
assign WBF =  BBF & ZZI & qxd  |  ABF & ZZI & QXD  ; 
assign wbf = ~WBF;  //complement 
assign WBN =  BBN & ZZI & qxd  |  ABN & ZZI & QXD  ; 
assign wbn = ~WBN;  //complement 
assign obf = ~OBF;  //complement 
assign obn = ~OBN;  //complement 
assign EAF = ~eaf;  //complement 
assign qba = ~QBA;  //complement 
assign EAN = ~ean;  //complement 
assign ECN = ~ecn;  //complement 
assign nae = ~NAE;  //complement 
assign RBA = ~rba;  //complement 
assign OCF = ~ocf;  //complement 
assign OCN = ~ocn;  //complement 
assign ODF = ~odf;  //complement 
assign ODN = ~odn;  //complement 
assign oga = ~OGA;  //complement 
assign ogb = ~OGB;  //complement 
assign qhc = ~QHC;  //complement 
assign qhd = ~QHD;  //complement 
assign oej = ~OEJ;  //complement 
assign ogc = ~OGC;  //complement 
assign ogd = ~OGD;  //complement 
assign qcd = ~QCD;  //complement 
assign oem = ~OEM;  //complement 
assign oef = ~OEF;  //complement 
assign OTE = ~ote;  //complement 
assign qqy = ~QQY;  //complement 
assign gdx = ~GDX;  //complement 
assign ogi = ~OGI;  //complement 
assign qqt = ~QQT;  //complement 
assign qqa = ~QQA;  //complement 
assign oep = ~OEP;  //complement 
assign laf = ~LAF;  //complement 
assign pag = ~PAG;  //complement 
assign pcg = ~PCG;  //complement 
assign peg = ~PEG;  //complement 
assign JGG =  QVC & PCE & PCF  ; 
assign jgg = ~JGG;  //complement  
assign JGO =  QVE & PCM & PCN  ; 
assign jgo = ~JGO;  //complement 
assign JDO =  QWE & BCM & BCN  ; 
assign jdo = ~JDO;  //complement 
assign pao = ~PAO;  //complement 
assign pco = ~PCO;  //complement 
assign peo = ~PEO;  //complement 
assign QVE = ~qve;  //complement 
assign bao = ~BAO;  //complement 
assign bco = ~BCO;  //complement 
assign beo = ~BEO;  //complement 
assign QWG = ~qwg;  //complement 
assign pbg = ~PBG;  //complement 
assign pdg = ~PDG;  //complement 
assign pfg = ~PFG;  //complement 
assign JFF =  PFE & PFF & PFG & PFH  ; 
assign jff = ~JFF;  //complement  
assign JFD =  PEM & PEN & PEO & PEP  ; 
assign jfd = ~JFD;  //complement 
assign bbg = ~BBG;  //complement 
assign bdg = ~BDG;  //complement 
assign bfg = ~BFG;  //complement 
assign JDC =  BEM & BEN & BEO & BEP  ; 
assign jdc = ~JDC;  //complement  
assign JUA =  GDA & GDB  ; 
assign jua = ~JUA;  //complement 
assign pbo = ~PBO;  //complement 
assign pdo = ~PDO;  //complement 
assign JHO =  QVG & QVJ & PDM & PDN  ; 
assign jho = ~JHO;  //complement  
assign JHG =  QVF & QVH & PDE & PDF  ; 
assign jhg = ~JHG;  //complement 
assign bbo = ~BBO;  //complement 
assign bdo = ~BDO;  //complement 
assign JEG =  QWG & BDE & BDF  ; 
assign jeg = ~JEG;  //complement  
assign JEO =  QWH & QWI & BDM & BDN  ; 
assign jeo = ~JEO;  //complement 
assign gda = ~GDA;  //complement 
assign gdb = ~GDB;  //complement 
assign gdd = ~GDD;  //complement 
assign gdg = ~GDG;  //complement 
assign gde = ~GDE;  //complement 
assign gdh = ~GDH;  //complement 
assign gdc = ~GDC;  //complement 
assign JVC =  GDY & GDD & GDE  ; 
assign jvc = ~JVC;  //complement 
assign JVB =  GDY & GDD  ; 
assign jvb = ~JVB;  //complement 
assign JVA =  GDY  ; 
assign jva = ~JVA;  //complement 
assign gdf = ~GDF;  //complement 
assign gdi = ~GDI;  //complement 
assign jvd =  GDD & hma  |  gdd & HMA  |  GDE & hmb  |  gde & HMB  |  GDF & hmc  |  gdf & HMC  ;
assign JVD = ~jvd;  //complement 
assign qkp = ~QKP;  //complement 
assign qkq = ~QKQ;  //complement 
assign qtf = ~QTF;  //complement 
assign qtg = ~QTG;  //complement 
assign qth = ~QTH;  //complement 
assign qti = ~QTI;  //complement 
assign aoh = ~AOH;  //complement 
assign aoi = ~AOI;  //complement 
assign aoj = ~AOJ;  //complement 
assign aok = ~AOK;  //complement 
assign ACO = ~aco;  //complement 
assign ADO = ~ado;  //complement 
assign ADG = ~adg;  //complement 
assign BMA =  aoh & ASH  |  asi & AOI  |  ASI & aoi  |  asj & AOJ  |  ASJ & aoj  |  ash & AOH  ;
assign bma = ~BMA;  //complement 
assign aol = ~AOL;  //complement 
assign aom = ~AOM;  //complement 
assign aon = ~AON;  //complement 
assign aoo = ~AOO;  //complement 
assign cia = ~CIA;  //complement 
assign BMC =  aon & ASN  |  asn & AON  |  AAO & aoo  |  aao & AOO  |  ASP & aop  |  asp & AOP  ;
assign bmc = ~BMC;  //complement 
assign aop = ~AOP;  //complement 
assign apa = ~APA;  //complement 
assign apb = ~APB;  //complement 
assign apc = ~APC;  //complement 
assign cib = ~CIB;  //complement 
assign BME =  apd & ATD  |  atd & APD  |  ATE & ape  |  ate & APE  |  ATF & apf  |  atf & APF  ;
assign bme = ~BME;  //complement 
assign apd = ~APD;  //complement 
assign ape = ~APE;  //complement 
assign apf = ~APF;  //complement 
assign apg = ~APG;  //complement 
assign aph = ~APH;  //complement 
assign api = ~API;  //complement 
assign apj = ~APJ;  //complement 
assign apk = ~APK;  //complement 
assign JOG =  cia & cib  ; 
assign jog = ~JOG;  //complement 
assign JOH =  cja & cjb  ; 
assign joh = ~JOH;  //complement 
assign JBO =  ADO  ; 
assign jbo = ~JBO;  //complement 
assign BMG =  apj & ATJ  |  atj & APJ  |  ATK & apk  |  atk & APK  |  ATL & apl  |  atl & APL  ;
assign bmg = ~BMG;  //complement 
assign apl = ~APL;  //complement 
assign apm = ~APM;  //complement 
assign apn = ~APN;  //complement 
assign apo = ~APO;  //complement 
assign rax = ~RAX;  //complement 
assign RAA = ~raa;  //complement 
assign RAT = ~rat;  //complement 
assign FAP =  EAL & EAK & EAJ  ; 
assign fap = ~FAP;  //complement 
assign QTB = ~qtb;  //complement 
assign qtc = ~QTC;  //complement 
assign qtd = ~QTD;  //complement 
assign qte = ~QTE;  //complement 
assign JIA =  QAA & GAC & gba  |  RJC  |  QYD  ; 
assign jia = ~JIA; //complement 
assign jch =  qqq & qqn & qta & qtx  ; 
assign JCH = ~jch;  //complement  
assign jke =  qnj & qnr & qnv  ; 
assign JKE = ~jke;  //complement 
assign qkr = ~QKR;  //complement 
assign QNB = ~qnb;  //complement 
assign QNC = ~qnc;  //complement 
assign QNF = ~qnf;  //complement 
assign QNG = ~qng;  //complement 
assign tme =  qto  ; 
assign TME = ~tme;  //complement 
assign tha =  rqb  ; 
assign THA = ~tha;  //complement 
assign JCS =  RQC  ; 
assign jcs = ~JCS;  //complement 
assign qma = ~QMA;  //complement 
assign qme = ~QME;  //complement 
assign qmi = ~QMI;  //complement 
assign tla =  qma & rsb & rqc  ; 
assign TLA = ~tla;  //complement  
assign tlc =  qmc & qnc & rsc & rqc  ; 
assign TLC = ~tlc;  //complement 
assign rqb = ~RQB;  //complement 
assign RQC = ~rqc;  //complement 
assign BMB =  ASK & aok  |  ask & AOK  |  ASL & aol  |  asl & AOL  |  ASM & aom  |  asm & AOM  ;
assign bmb = ~BMB;  //complement 
assign aag = ~AAG;  //complement 
assign ohe = ~OHE;  //complement 
assign WAG =  ZZO & ZZI & qxc  |  AAG & ZZI & QXC  ; 
assign wag = ~WAG;  //complement 
assign WAO =  BAO & ZZI & qxc  |  AAO & ZZI & QXC  ; 
assign wao = ~WAO;  //complement 
assign oag = ~OAG;  //complement 
assign oao = ~OAO;  //complement 
assign BMD =  ATA & apa  |  ata & APA  |  ATB & apb  |  atb & APB  |  ATC & apc  |  atc & APC  ;
assign bmd = ~BMD;  //complement 
assign aso = ~ASO;  //complement 
assign aao = ~AAO;  //complement 
assign tec = qeb; 
assign TEC = ~tec; //complement 
assign ted = qeb; 
assign TED = ~ted;  //complement 
assign tea = qea; 
assign TEA = ~tea;  //complement 
assign teb = qea; 
assign TEB = ~teb;  //complement 
assign wcg = aag; 
assign WCG = ~wcg; //complement 
assign wco = aao; 
assign WCO = ~wco;  //complement 
assign wdg = abg; 
assign WDG = ~wdg;  //complement 
assign wdo = abo; 
assign WDO = ~wdo;  //complement 
assign BMF =  ABG & apg  |  abg & APG  |  ATH & aph  |  ath & APH  |  ATI & api  |  ati & API  ;
assign bmf = ~BMF;  //complement 
assign atg = ~ATG;  //complement 
assign abg = ~ABG;  //complement 
assign dag = ~DAG;  //complement 
assign dao = ~DAO;  //complement 
assign dbg = ~DBG;  //complement 
assign dbo = ~DBO;  //complement 
assign QSI = ~qsi;  //complement 
assign QQX = ~qqx;  //complement 
assign qto = ~QTO;  //complement 
assign qtn = ~QTN;  //complement 
assign BMH =  ATM & apm  |  atm & APM  |  ATN & apn  |  atn & APN  |  ABO & apo  |  abo & APO  ;
assign bmh = ~BMH;  //complement 
assign ato = ~ATO;  //complement 
assign abo = ~ABO;  //complement 
assign WBG =  BBG & ZZI & qxd  |  ABG & ZZI & QXD  ; 
assign wbg = ~WBG;  //complement 
assign WBO =  BBO & ZZI & qxd  |  ABO & ZZI & QXD  ; 
assign wbo = ~WBO;  //complement 
assign obg = ~OBG;  //complement 
assign obo = ~OBO;  //complement 
assign edg = ~EDG;  //complement 
assign edo = ~EDO;  //complement 
assign EAG = ~eag;  //complement 
assign ECO = ~eco;  //complement 
assign qaa = ~QAA;  //complement 
assign qab = ~QAB;  //complement 
assign qac = ~QAC;  //complement 
assign qad = ~QAD;  //complement 
assign qea = ~QEA;  //complement 
assign qeb = ~QEB;  //complement 
assign OCG = ~ocg;  //complement 
assign OCO = ~oco;  //complement 
assign ODG = ~odg;  //complement 
assign ODO = ~odo;  //complement 
assign JXA =  QLN & QSD  ; 
assign jxa = ~JXA;  //complement 
assign jab =  qad  ; 
assign JAB = ~jab;  //complement 
assign JQF =  QQB & qtp  ; 
assign jqf = ~JQF;  //complement 
assign qsa = ~QSA;  //complement 
assign oes = ~OES;  //complement 
assign OLD = ~old;  //complement 
assign ofc = ~OFC;  //complement 
assign oqb = ~OQB;  //complement 
assign olb = ~OLB;  //complement 
assign OTF = ~otf;  //complement 
assign gdj = ~GDJ;  //complement 
assign gdk = ~GDK;  //complement 
assign gdl = ~GDL;  //complement 
assign qcj = ~QCJ;  //complement 
assign qsb = ~QSB;  //complement 
assign oet = ~OET;  //complement 
assign oeh = ~OEH;  //complement 
assign OEQ = ~oeq;  //complement 
assign OER = ~oer;  //complement 
assign qtj = ~QTJ;  //complement 
assign kaf = ~KAF;  //complement 
assign qtx = ~QTX;  //complement 
assign qtp = ~QTP;  //complement 
assign ofa = ~OFA;  //complement 
assign OFB = ~ofb;  //complement 
assign OQA = ~oqa;  //complement 
assign pah = ~PAH;  //complement 
assign pch = ~PCH;  //complement 
assign peh = ~PEH;  //complement 
assign JGH =  QVC & PCE & PCF & PCG  ; 
assign jgh = ~JGH;  //complement  
assign JGP =  QVE & PCM & PCN & PCO  ; 
assign jgp = ~JGP;  //complement 
assign bah = ~BAH;  //complement 
assign beh = ~BEH;  //complement 
assign JDH =  QWC  ; 
assign jdh = ~JDH;  //complement  
assign JDP =  QWE & BCM & BCN & BCO  ; 
assign jdp = ~JDP;  //complement 
assign pap = ~PAP;  //complement 
assign pcp = ~PCP;  //complement 
assign pep = ~PEP;  //complement 
assign QVF = ~qvf;  //complement 
assign QVG = ~qvg;  //complement 
assign bap = ~BAP;  //complement 
assign bep = ~BEP;  //complement 
assign ola = ~OLA;  //complement 
assign pbh = ~PBH;  //complement 
assign pdh = ~PDH;  //complement 
assign pfh = ~PFH;  //complement 
assign JHH =  QVF & QVH & PDE & PDF & PDG  ; 
assign jhh = ~JHH;  //complement  
assign JFB =  PEE & PEF & PEG & PEH  ; 
assign jfb = ~JFB;  //complement 
assign bbh = ~BBH;  //complement 
assign bfh = ~BFH;  //complement 
assign JDA =  BEH & QWB  ; 
assign jda = ~JDA;  //complement  
assign JDE =  BFE & BFF & BFG & BFH  ; 
assign jde = ~JDE;  //complement 
assign pbp = ~PBP;  //complement 
assign pdp = ~PDP;  //complement 
assign JHP =  QVG & QVJ & PDM & PDN & PDO  ; 
assign jhp = ~JHP;  //complement  
assign bbp = ~BBP;  //complement 
assign JEP =  QWH & QWI & BDM & BDN & BDO  ; 
assign jep = ~JEP;  //complement  
assign JEH =  QWG & BDE & BDF & BDG  ; 
assign jeh = ~JEH;  //complement 
assign JQI =  QQH & qqc  ; 
assign jqi = ~JQI;  //complement 
assign JQJ =  QQJ & qqk  ; 
assign jqj = ~JQJ;  //complement 
assign hna = ~HNA;  //complement 
assign hnb = ~HNB;  //complement 
assign hnc = ~HNC;  //complement 
assign qsc = ~QSC;  //complement 
assign qsd = ~QSD;  //complement 
assign hpa = ~HPA;  //complement 
assign hpb = ~HPB;  //complement 
assign hpc = ~HPC;  //complement 
assign qsf = ~QSF;  //complement 
assign rsb = ~RSB;  //complement 
assign qsg = ~QSG;  //complement 
assign qqk = ~QQK;  //complement 
assign qqr = ~QQR;  //complement 
assign hoa = ~HOA;  //complement 
assign hob = ~HOB;  //complement 
assign hoc = ~HOC;  //complement 
assign rre = ~RRE;  //complement 
assign rrf = ~RRF;  //complement 
assign RRG = ~rrg;  //complement 
assign rrh = ~RRH;  //complement 
assign rrb = ~RRB;  //complement 
assign rsc = ~RSC;  //complement 
assign rrc = ~RRC;  //complement 
assign rrd = ~RRD;  //complement 
assign aqh = ~AQH;  //complement 
assign aqi = ~AQI;  //complement 
assign aqj = ~AQJ;  //complement 
assign aqk = ~AQK;  //complement 
assign ACH = ~ach;  //complement 
assign ACP = ~acp;  //complement 
assign ADH = ~adh;  //complement 
assign BNA =  AAH & aqh  |  asi & AQI  |  ASI & aqi  |  asj & AQJ  |  ASJ & aqj  |  aah & AQH  ;
assign bna = ~BNA;  //complement 
assign aql = ~AQL;  //complement 
assign aqm = ~AQM;  //complement 
assign aqn = ~AQN;  //complement 
assign aqo = ~AQO;  //complement 
assign cja = ~CJA;  //complement 
assign BNC =  aqn & ASN  |  asn & AQN  |  ASO & aqo  |  aso & AQO  |  AAP & aqp  |  aap & AQP  ;
assign bnc = ~BNC;  //complement 
assign aqp = ~AQP;  //complement 
assign ara = ~ARA;  //complement 
assign arb = ~ARB;  //complement 
assign arc = ~ARC;  //complement 
assign cjb = ~CJB;  //complement 
assign BNE =  ard & ATD  |  atd & ARD  |  ATE & are  |  ate & ARE  |  ATF & arf  |  atf & ARF  ;
assign bne = ~BNE;  //complement 
assign ard = ~ARD;  //complement 
assign are = ~ARE;  //complement 
assign arf = ~ARF;  //complement 
assign arg = ~ARG;  //complement 
assign arh = ~ARH;  //complement 
assign ari = ~ARI;  //complement 
assign arj = ~ARJ;  //complement 
assign ark = ~ARK;  //complement 
assign JOD =  cfa & cfb  ; 
assign jod = ~JOD;  //complement 
assign JOE =  cga & cgb  ; 
assign joe = ~JOE;  //complement 
assign JOF =  cha & chb  ; 
assign jof = ~JOF;  //complement 
assign BNG =  arj & ATJ  |  atj & ARJ  |  ATK & ark  |  atk & ARK  |  ATL & arl  |  atl & ARL  ;
assign bng = ~BNG;  //complement 
assign arl = ~ARL;  //complement 
assign arm = ~ARM;  //complement 
assign arn = ~ARN;  //complement 
assign aro = ~ARO;  //complement 
assign JQH =  RBE & QQF  |  RBI  ; 
assign jqh = ~JQH;  //complement 
assign qqj = ~QQJ;  //complement 
assign qqh = ~QQH;  //complement 
assign rbf = ~RBF;  //complement 
assign rbg = ~RBG;  //complement 
assign rbh = ~RBH;  //complement 
assign rbi = ~RBI;  //complement 
assign qsh = ~QSH;  //complement 
assign qse = ~QSE;  //complement 
assign qqn = ~QQN;  //complement 
assign qqm = ~QQM;  //complement 
assign JQC =  qql & qlx  ; 
assign jqc = ~JQC;  //complement  
assign JQB =  qql & qlp & qqw  ; 
assign jqb = ~JQB;  //complement 
assign qql = ~QQL;  //complement 
assign qqs = ~QQS;  //complement 
assign RQA = ~rqa;  //complement 
assign BNB =  ASK & aqk  |  ask & AQK  |  ASL & aql  |  asl & AQL  |  ASM & aqm  |  asm & AQM  ;
assign bnb = ~BNB;  //complement 
assign ash = ~ASH;  //complement 
assign aah = ~AAH;  //complement 
assign WAH =  BAH & ZZI & qxc  |  AAH & ZZI & QXC  ; 
assign wah = ~WAH;  //complement 
assign WAP =  BAP & ZZI & qxc  |  AAP & ZZI & QXC  ; 
assign wap = ~WAP;  //complement 
assign oah = ~OAH;  //complement 
assign oap = ~OAP;  //complement 
assign BND =  ATA & ara  |  ata & ARA  |  ATB & arb  |  atb & ARB  |  ATC & arc  |  atc & ARC  ;
assign bnd = ~BND;  //complement 
assign asp = ~ASP;  //complement 
assign aap = ~AAP;  //complement 
assign tma = qtn; 
assign TMA = ~tma; //complement 
assign tmb = qtn; 
assign TMB = ~tmb;  //complement 
assign tmc = qtn; 
assign TMC = ~tmc;  //complement 
assign tmd = qtn; 
assign TMD = ~tmd;  //complement 
assign wch = aah; 
assign WCH = ~wch; //complement 
assign wcp = aap; 
assign WCP = ~wcp;  //complement 
assign wdh = abh; 
assign WDH = ~wdh;  //complement 
assign wdp = abp; 
assign WDP = ~wdp;  //complement 
assign BNF =  ATG & arg  |  atg & ARG  |  ABH & arh  |  abh & ARH  |  ATI & ari  |  ati & ARI  ;
assign bnf = ~BNF;  //complement 
assign ath = ~ATH;  //complement 
assign abh = ~ABH;  //complement 
assign dah = ~DAH;  //complement 
assign dap = ~DAP;  //complement 
assign dbh = ~DBH;  //complement 
assign dbp = ~DBP;  //complement 
assign TEE = QQX; 
assign tee = ~TEE; //complement 
assign TEF = QQX; 
assign tef = ~TEF;  //complement 
assign BNH =  ATM & arm  |  atm & ARM  |  ATN & arn  |  atn & ARN  |  ATO & aro  |  ato & ARO  ;
assign bnh = ~BNH;  //complement 
assign abp = ~ABP;  //complement 
assign atp = ~ATP;  //complement 
assign WBH =  BBH & ZZI & qxd  |  ABH & ZZI & QXD  ; 
assign wbh = ~WBH;  //complement 
assign WBP =  BBP & ZZI & qxd  |  ABP & ZZI & QXD  ; 
assign wbp = ~WBP;  //complement 
assign obh = ~OBH;  //complement 
assign obp = ~OBP;  //complement 
assign EAH = ~eah;  //complement 
assign EAP = ~eap;  //complement 
assign EBP = ~ebp;  //complement 
assign ogj = ~OGJ;  //complement 
assign edh = ~EDH;  //complement 
assign edp = ~EDP;  //complement 
assign qkt = ~QKT;  //complement 
assign OCH = ~och;  //complement 
assign OCP = ~ocp;  //complement 
assign ODH = ~odh;  //complement 
assign ODP = ~odp;  //complement 
assign oge = ~OGE;  //complement 
assign ogf = ~OGF;  //complement 
assign JIE = qcy & RLD ; 
assign jie = ~JIE ; //complement 
assign oeg = ~OEG;  //complement 
assign qfc = ~QFC;  //complement 
assign ogg = ~OGG;  //complement 
assign ogh = ~OGH;  //complement 
assign qch = ~QCH;  //complement 
assign oev = ~OEV;  //complement 
assign oel = ~OEL;  //complement 
assign oen = ~OEN;  //complement 
assign oeo = ~OEO;  //complement 
assign oex = ~OEX;  //complement 
assign oey = ~OEY;  //complement 
assign rra = ~RRA;  //complement 
assign rsa = ~RSA;  //complement 
assign QLX = ~qlx;  //complement 
assign tlb = rsa; 
assign TLB = ~tlb;  //complement 
assign oek = ~OEK;  //complement 
assign oeu = ~OEU;  //complement 
assign oew = ~OEW;  //complement 
assign iaa = ~IAA; //complement 
assign iab = ~IAB; //complement 
assign iac = ~IAC; //complement 
assign iad = ~IAD; //complement 
assign iae = ~IAE; //complement 
assign iaf = ~IAF; //complement 
assign iag = ~IAG; //complement 
assign iah = ~IAH; //complement 
assign iai = ~IAI; //complement 
assign iaj = ~IAJ; //complement 
assign iak = ~IAK; //complement 
assign ial = ~IAL; //complement 
assign iam = ~IAM; //complement 
assign ian = ~IAN; //complement 
assign iao = ~IAO; //complement 
assign iap = ~IAP; //complement 
assign iba = ~IBA; //complement 
assign ibb = ~IBB; //complement 
assign ibc = ~IBC; //complement 
assign ibd = ~IBD; //complement 
assign ibe = ~IBE; //complement 
assign ibf = ~IBF; //complement 
assign ibg = ~IBG; //complement 
assign ibh = ~IBH; //complement 
assign ibi = ~IBI; //complement 
assign ibj = ~IBJ; //complement 
assign ibk = ~IBK; //complement 
assign ibl = ~IBL; //complement 
assign ibm = ~IBM; //complement 
assign ibn = ~IBN; //complement 
assign ibo = ~IBO; //complement 
assign ibp = ~IBP; //complement 
assign ica = ~ICA; //complement 
assign icb = ~ICB; //complement 
assign icc = ~ICC; //complement 
assign icd = ~ICD; //complement 
assign ice = ~ICE; //complement 
assign icf = ~ICF; //complement 
assign icg = ~ICG; //complement 
assign ich = ~ICH; //complement 
assign ici = ~ICI; //complement 
assign icj = ~ICJ; //complement 
assign ick = ~ICK; //complement 
assign icl = ~ICL; //complement 
assign icm = ~ICM; //complement 
assign icn = ~ICN; //complement 
assign ico = ~ICO; //complement 
assign icp = ~ICP; //complement 
assign ida = ~IDA; //complement 
assign idb = ~IDB; //complement 
assign idc = ~IDC; //complement 
assign idd = ~IDD; //complement 
assign ide = ~IDE; //complement 
assign idf = ~IDF; //complement 
assign idg = ~IDG; //complement 
assign idh = ~IDH; //complement 
assign idi = ~IDI; //complement 
assign idj = ~IDJ; //complement 
assign idk = ~IDK; //complement 
assign idl = ~IDL; //complement 
assign idm = ~IDM; //complement 
assign idn = ~IDN; //complement 
assign ido = ~IDO; //complement 
assign idp = ~IDP; //complement 
assign iea = ~IEA; //complement 
assign ieb = ~IEB; //complement 
assign iec = ~IEC; //complement 
assign ied = ~IED; //complement 
assign iee = ~IEE; //complement 
assign ief = ~IEF; //complement 
assign ieg = ~IEG; //complement 
assign ieh = ~IEH; //complement 
assign iei = ~IEI; //complement 
assign iej = ~IEJ; //complement 
assign iek = ~IEK; //complement 
assign iel = ~IEL; //complement 
assign iem = ~IEM; //complement 
assign ien = ~IEN; //complement 
assign ieo = ~IEO; //complement 
assign iep = ~IEP; //complement 
assign ifa = ~IFA; //complement 
assign ifb = ~IFB; //complement 
assign ifc = ~IFC; //complement 
assign ifd = ~IFD; //complement 
assign ife = ~IFE; //complement 
assign ifff  = ~IFFF ; //complement 
assign ifg = ~IFG; //complement 
assign ifh = ~IFH; //complement 
assign ifi = ~IFI; //complement 
assign iga = ~IGA; //complement 
assign igb = ~IGB; //complement 
assign igc = ~IGC; //complement 
assign ihb = ~IHB; //complement 
assign ihc = ~IHC; //complement 
assign ija = ~IJA; //complement 
assign ijb = ~IJB; //complement 
assign ijc = ~IJC; //complement 
assign ijd = ~IJD; //complement 
assign ika = ~IKA; //complement 
assign ikb = ~IKB; //complement 
assign ila = ~ILA; //complement 
assign ilb = ~ILB; //complement 
assign ilc = ~ILC; //complement 
assign ima = ~IMA; //complement 
assign imb = ~IMB; //complement 
assign imc = ~IMC; //complement 
assign imd = ~IMD; //complement 
assign ime = ~IME; //complement 
assign imf = ~IMF; //complement 
assign img = ~IMG; //complement 
assign ina = ~INA; //complement 
assign ioa = ~IOA; //complement 
assign iob = ~IOB; //complement 
assign ioc = ~IOC; //complement 
assign iod = ~IOD; //complement 
assign ipa = ~IPA; //complement 
assign ipb = ~IPB; //complement 
assign ipc = ~IPC; //complement 
assign ipd = ~IPD; //complement 
assign ipe = ~IPE; //complement 
assign ipf = ~IPF; //complement 
assign iqa = ~IQA; //complement 
assign iqb = ~IQB; //complement 
assign iqc = ~IQC; //complement 
assign iqd = ~IQD; //complement 
assign iqe = ~IQE; //complement 
assign iqf = ~IQF; //complement 
assign iqg = ~IQG; //complement 
assign iqh = ~IQH; //complement 
assign iqi = ~IQI; //complement 
assign izz = ~IZZ; //complement 
always@(posedge IZZ )
   begin 
 PAA <=  PAA & jga & tpa  |  paa & JGA  |  AAA & TPA  ; 
 PCA <=  PAA & jga & tpa  |  paa & JGA  |  AAA & TPA  ; 
 PAI <=  PAI & jgi & tpb  |  pai & JGI  |  AAI & TPB  ; 
 PCI <=  PAI & jgi & tpb  |  pai & JGI  |  AAI & TPB  ; 
 PEI <=  PAI & jgi & tpb  |  pai & JGI  |  AAI & TPB  ; 
 qva <=  qua  ; 
 qvj <=  jfe  |  jff  |  jfg  ; 
 BAI <=  BAI & jdi & tfb  |  bai & JDI  |  AAI & TFB  ; 
 BCI <=  BAI & jdi & tfb  |  bai & JDI  |  AAI & TFB  ; 
 BEI <=  BAI & jdi & tfb  |  bai & JDI  |  AAI & TFB  ; 
 haa <=  GAB  |  GAA  ; 
 hab <=  GAB  |  gaa  ; 
 PBA <=  PBA & jha & tpc  |  pba & JHA  |  ABA & TPC  ; 
 PDA <=  PBA & jha & tpc  |  pba & JHA  |  ABA & TPC  ; 
 PFA <=  PBA & jha & tpc  |  pba & JHA  |  ABA & TPC  ; 
 BBA <=  BBA & jea & tfc  |  bba & JEA  |  ABA & TFC  ; 
 BDA <=  BBA & jea & tfc  |  bba & JEA  |  ABA & TFC  ; 
 BFA <=  BBA & jea & tfc  |  bba & JEA  |  ABA & TFC  ; 
 hac <=  gab  |  GAA  ; 
 had <=  gab  |  gaa  ; 
 PBI <=  PBI & jhi & tpd  |  pbi & JHI  |  ABI & TPD  ; 
 PDI <=  PBI & jhi & tpd  |  pbi & JHI  |  ABI & TPD  ; 
 PFI <=  PBI & jhi & tpd  |  pbi & JHI  |  ABI & TPD  ; 
 BBI <=  BBI & jei & tfd  |  bbi & JEI  |  ABI & TFD  ; 
 BDI <=  BBI & jei & tfd  |  bbi & JEI  |  ABI & TFD  ; 
 BFI <=  BBI & jei & tfd  |  bbi & JEI  |  ABI & TFD  ; 
 hba <= haa ; 
 hca <= hba ; 
 hda <= hca ; 
 hea <= hda ; 
 hbb <= hab ; 
 hcb <= hbb ; 
 hdb <= hcb ; 
 heb <= hdb ; 
 hbc <= hac ; 
 hcc <= hbc ; 
 hdc <= hcc ; 
 hbh <= hah ; 
 hbe <= hae ; 
 hce <= hbe ; 
 hde <= hce ; 
 hbd <= had ; 
 hbf <= haf ; 
 hcf <= hbf ; 
 hdf <= hcf ; 
 hcd <= hbd ; 
 hbg <= hag ; 
 hcg <= hbg ; 
 hdd <= hcd ; 
 hch <= hbh ; 
 hdh <= hch ; 
 heh <= hdh ; 
 HAE <= QAD & GAM ; 
 HAF <= QAD & GAN ; 
 HAG <= QAD & GAO ; 
 HAH <= QAD & GAP ; 
 LBA <=  LBA & jla & tla  |  lba & JLA  |  LAA & TLA  ; 
 aci <= wci & QKR |  aqi & qkr ; 
 ada <= wda & QKR |  ara & qkr ; 
 adi <= wdi & QKR |  ari & qkr ; 
 CCA <=  BGD  |  ZZI & BGB  |  BGA  |  ZZO & ZZI  |  BGC  ; 
 CCB <=  BGH  |  BGE  |  BGF  |  ZZO & ZZI  |  BGG  ; 
 gaa <= fbg & TGA |  gaa & tga ; 
 gai <= eai & TGA |  gai & tga ; 
 gab <= fbh & TGA |  gab & tga ; 
 gao <=  fab & TGB  |  FBE & TGD  |  gao & tgb  ; 
 gbh <=  fae & TGB  |  fba & TGD  |  gbh & tgb  ; 
 gci <=  eaa & TGC  |  ZZO & TGE  |  gci & tgc  ; 
 gam <=  fad & TGC  |  FBE & TGE  |  gam & tgc  ; 
 HDI <= HCG & HCA ; 
 HDJ <= HCG & HCB ; 
 HDK <= HCG & HCC ; 
 HDL <= HCG & HCD ; 
 QQI <= JJD & RLA ; 
 QTA <=  QTA & qtx  |  GCH & QAD  |  IMB  ; 
 RJA <=  ZZO & qtx  |  GBA & QAD  ; 
 QND <=  QNC  ; 
 qoa <=  rld  |  QND  ; 
 AAA <=  IAA & TAA  |  DAA & TBA  |  IEA & TCA  |  WAA & TDA  |  TMA  ; 
 OAA <=  DAA & TEA  |  EAA & TEC  |  NAA & TEE  ; 
 OAI <=  DAI & TEA  |  ECI & TEC  |  WCK & TEE  ; 
 ASI <=  IAI & TAB  |  DAI & TBB  |  IEI & TCB  |  WAI & TDB  |  TMB  ; 
 AAI <=  IAI & TAB  |  DAI & TBB  |  IEI & TCB  |  WAI & TDB  |  TMB  ; 
 ATA <=  IBA & TAC  |  DBA & TBC  |  EAA & TCC  |  WBA & TDC  |  TMC  ; 
 ABA <=  IBA & TAC  |  DBA & TBC  |  EAA & TCC  |  WBA & TDC  |  TMC  ; 
 DAA <= ICA ; 
 DAI <= ICI ; 
 DBA <= IDA ; 
 DBI <= IDI ; 
 ora <= gci ; 
 OTB <= QTW ; 
 EDI <= ECI ; 
 qza <= qya ; 
 ATI <=  IBI & TAD  |  DBI & TBD  |  ECI & TCD  |  WBI & TDD  |  TMD  ; 
 ABI <=  IBI & TAD  |  DBI & TBD  |  ECI & TCD  |  WBI & TDD  |  TMD  ; 
 OBA <=  DBA & TEB  |  EDA & TED  |  WDC & TEF  ; 
 OBI <=  DBI & TEB  |  EDI & TED  |  WDK & TEF  ; 
 eaa <= iea ; 
 eai <= iei ; 
 eci <= iei ; 
 NAA <=  NAA & jsa & tha  |  naa & JSA  |  WCC & THA  ; 
 NBA <=  NAA & jsa & tha  |  naa & JSA  |  WCC & THA  ; 
 NCA <=  NAA & jsa & tha  |  naa & JSA  |  WCC & THA  ; 
 QZE <=  QZE & qzd  |  QYA  ; 
 rje <=  rjd & qzd  ; 
 QYA <= IMC ; 
 QYB <= IMD ; 
 QYC <= IME ; 
 QYD <= IMF ; 
 EDA <= EAA ; 
 RJD <= JJC ; 
 oca <= pca ; 
 oci <= pci ; 
 oda <= pda ; 
 odi <= pdi ; 
 HEO <= HDH & HDC ; 
 HEP <= HDH & HDD ; 
 QGE <=  IGC & HDL  |  igc & HDK  |  ZZO & igb  ; 
 qgd <=  ZZO & HDL  |  ZZO & HDK  |  iga & igb  ; 
 RJK <=  RJK & rjl & jct  |  RJA  ; 
 OEA <= KAA ; 
 qzd <= qyd ; 
 RJB <= RJA ; 
 QTM <= IMA ; 
 KAA <=  KAA & tlc & jma  |  kaa & JMA  |  JNA  ; 
 RJF <= RJE ; 
 RJG <= RJF ; 
 RJH <= RJG ; 
 RJI <= RJH ; 
 LAA <=  IPA & tlb & jcr  |  IQA & TLB  ; 
 PAB <=  PAB & jgb & tpa  |  pab & JGB  |  AAB & TPA  ; 
 PCB <=  PAB & jgb & tpa  |  pab & JGB  |  AAB & TPA  ; 
 PEB <=  PAB & jgb & tpa  |  pab & JGB  |  AAB & TPA  ; 
 PAJ <=  PAJ & jgj & tpb  |  paj & JGJ  |  AAJ & TPB  ; 
 PCJ <=  PAJ & jgj & tpb  |  paj & JGJ  |  AAJ & TPB  ; 
 PEJ <=  PAJ & jgj & tpb  |  paj & JGJ  |  AAJ & TPB  ; 
 qvh <=  jfe  ; 
 qvi <=  jfe  |  jff  ; 
 BAJ <=  BAJ & jdj & tfb  |  baj & JDJ  |  AAJ & TFB  ; 
 BCJ <=  BAJ & jdj & tfb  |  baj & JDJ  |  AAJ & TFB  ; 
 BEJ <=  BAJ & jdj & tfb  |  baj & JDJ  |  AAJ & TFB  ; 
 PBB <=  PBB & jhb & tpc  |  pbb & JHB  |  ABB & TPC  ; 
 PDB <=  PBB & jhb & tpc  |  pbb & JHB  |  ABB & TPC  ; 
 PFB <=  PBB & jhb & tpc  |  pbb & JHB  |  ABB & TPC  ; 
 BBB <=  BBB & jeb & tfc  |  bbb & JEB  |  ABB & TFC  ; 
 BDB <=  BBB & jeb & tfc  |  bbb & JEB  |  ABB & TFC  ; 
 BFB <=  BBB & jeb & tfc  |  bbb & JEB  |  ABB & TFC  ; 
 PBJ <=  PBJ & jhj & tpd  |  pbj & JHJ  |  ABJ & TPD  ; 
 PDJ <=  PBJ & jhj & tpd  |  pbj & JHJ  |  ABJ & TPD  ; 
 PFJ <=  PBJ & jhj & tpd  |  pbj & JHJ  |  ABJ & TPD  ; 
 BBJ <=  BBJ & jej & tfd  |  bbj & JEJ  |  ABJ & TFD  ; 
 BDJ <=  BBJ & jej & tfd  |  bbj & JEJ  |  ABJ & TFD  ; 
 BFJ <=  BBJ & jej & tfd  |  bbj & JEJ  |  ABJ & TFD  ; 
 RHA <= QHA ; 
 RHB <= RHA ; 
 RHC <= RHB ; 
 RHD <= RHC ; 
 RHE <= RHD ; 
 RHF <= RHE ; 
 RHG <= RHF ; 
 RHH <= RHG ; 
 RHI <= RHH ; 
 RHJ <= RHI ; 
 QHA <=  RHJ & QRC  |  QLD & qlk  |  JFX & QAB  |  JJH & qrc  ; 
 QKK <=  QKA & jic & jid  |  QKK & qkn  ; 
 RID <= RHC & QIC |  RIC & qic ; 
 RIE <= RHD & QIC |  RID & qic ; 
 RIF <= RHE & QIC |  RIE & qic ; 
 QTW <=  JIC  |  JID  ; 
 QKL <= QKK ; 
 QKM <= QKL ; 
 QKN <= QKM ; 
 RIA <= QHA & QIC |  ZZO & qic ; 
 RIB <= RHA & QIC |  RIA & qic ; 
 RIC <= RHB & QIC |  RIB & qic ; 
 LBB <=  LBB & jlb & tla  |  lbb & JLB  |  LAB & TLA  ; 
 AEH <= ACH ; 
 AEI <= ACI ; 
 AEJ <= ACJ ; 
 AEK <= ACK ; 
 acj <= wcj & QKR |  aqj & qkr ; 
 adb <= wdb & QKR |  arb & qkr ; 
 adj <= wdj & QKR |  arj & qkr ; 
 AEL <= ACL ; 
 AEM <= ACM ; 
 AEN <= ACN ; 
 AEO <= ACO ; 
 CDA <=  BHD  |  ZZI & BHB  |  BHA  |  ZZO & ZZI  |  BHC  ; 
 AEP <= ACP ; 
 AFA <= ADA ; 
 AFB <= ADB ; 
 AFC <= ADC ; 
 CDB <=  BHH  |  BHE  |  BHF  |  ZZO & ZZI  |  BHG  ; 
 AFD <= ADD ; 
 AFE <= ADE ; 
 AFF <= ADF ; 
 AFG <= ADG ; 
 AFH <= ADH ; 
 AFI <= ADI ; 
 AFJ <= ADJ ; 
 AFK <= ADK ; 
 AFL <= ADL ; 
 AFM <= ADM ; 
 AFN <= ADN ; 
 AFO <= JBO ; 
 gbj <=  faf & TGB  |  TGD & fbc  |  gbj & tgb  ; 
 gbi <=  fae & TGB  |  TGD & fbc  |  gbi & tgb  ; 
 gbp <=  fah & TGC  |  fal & TGE  |  gbp & tgc  ; 
 gbe <=  fae & TGC  |  fbb & TGE  |  gbe & tgc  ; 
 QKG <= JAE ; 
 QKH <= JAF ; 
 QKF <=  QKF & haf  |  QKC & QKD  ; 
 HEI <= HDI ; 
 HEJ <= HDJ ; 
 AAB <=  IAB & TAA  |  DAB & TBA  |  IEB & TCA  |  WAB & TDA  |  TMA  ; 
 OAB <=  DAB & TEA  |  EAB & TEC  |  NAB & TEE  ; 
 OAJ <=  DAJ & TEA  |  ECJ & TEC  |  WCL & TEE  ; 
 ASJ <=  IAJ & TAB  |  DAJ & TBB  |  IEJ & TCB  |  WAJ & TDB  |  TMB  ; 
 AAJ <=  IAJ & TAB  |  DAJ & TBB  |  IEJ & TCB  |  WAJ & TDB  |  TMB  ; 
 ATB <=  IBB & TAC  |  DBB & TBC  |  EAB & TCC  |  WBB & TDC  |  TMC  ; 
 ABB <=  IBB & TAC  |  DBB & TBC  |  EAB & TCC  |  WBB & TDC  |  TMC  ; 
 DAB <= ICB ; 
 DAJ <= ICJ ; 
 DBB <= IDB ; 
 DBJ <= IDJ ; 
 orb <= gcj ; 
 EDB <= EAB ; 
 EDJ <= ECJ ; 
 ATJ <=  IBJ & TAD  |  DBJ & TBD  |  ECJ & TCD  |  WBJ & TDD  |  TMD  ; 
 ABJ <=  IBJ & TAD  |  DBJ & TBD  |  ECJ & TCD  |  WBJ & TDD  |  TMD  ; 
 OBB <=  DBB & TEB  |  EDB & TED  |  WDD & TEF  ; 
 OBJ <=  DBJ & TEB  |  EDJ & TED  |  WDL & TEF  ; 
 eab <= ieb ; 
 eaj <= iej ; 
 ebj <= iej ; 
 ecj <= iej ; 
 NAB <=  NAB & jsb & tha  |  nab & JSB  |  WCD & THA  ; 
 NBB <=  NAB & jsb & tha  |  nab & JSB  |  WCD & THA  ; 
 NCB <=  NAB & jsb & tha  |  nab & JSB  |  WCD & THA  ; 
 QXE <=  JAB & JAC  ; 
 QXF <=  JAB & JAC  |  JJC  |  QYA  ; 
 ocb <= pcb ; 
 ocj <= pcj ; 
 odb <= pdb ; 
 odj <= pdj ; 
 QKX <=  JAD  |  RJG  |  RBB  ; 
 QKJ <=  ifi & JBX  |  IFI & JBY  |  JBE  |  JBB & rbc  ; 
 OJE <=  ifi & JBX  |  IFI & JBY  |  JBE  |  JBB & rbc  ; 
 QGA <=  ifa  |  ifb  |  ifc  |  ifd  ; 
 RFB <=  RFB & jcz  |  WCB & JCZ  ; 
 OJB <=  RFB & jcz  |  WCB & JCZ  ; 
 OEB <= KAB ; 
 CAA <= ILA ; 
 CAB <= ILB ; 
 CAC <= ILC ; 
 KAB <=  KAB & tlc & jmb  |  kab & JMB  |  JNB  ; 
 RFA <=  RFA & jcz  |  WCA & JCZ  ; 
 OJA <=  RFA & jcz  |  WCA & JCZ  ; 
 RGA <= INA ; 
 RGB <= RGA ; 
 RGC <= RGB ; 
 RGD <= RGC ; 
 LAB <=  IPB & tlb & jcr  |  IQB & TLB  ; 
 PAC <=  PAC & jgc & tpa  |  pac & JGC  |  AAC & TPA  ; 
 PCC <=  PAC & jgc & tpa  |  pac & JGC  |  AAC & TPA  ; 
 PEC <=  PAC & jgc & tpa  |  pac & JGC  |  AAC & TPA  ; 
 PAK <=  PAK & jgk & tpb  |  pak & JGK  |  AAK & TPB  ; 
 PCK <=  PAK & jgk & tpb  |  pak & JGK  |  AAK & TPB  ; 
 PEK <=  PAK & jgk & tpb  |  pak & JGK  |  AAK & TPB  ; 
 QUB <= QPD ; 
 QUC <= QUB ; 
 QUE <= QUD ; 
 qvb <= quf ; 
 BAK <=  BAK & jdk & tfb  |  bak & JDK  |  AAK & TFB  ; 
 BCK <=  BAK & jdk & tfb  |  bak & JDK  |  AAK & TFB  ; 
 BEK <=  BAK & jdk & tfb  |  bak & JDK  |  AAK & TFB  ; 
 QPA <= QAB & ZZI ; 
 QPB <= QAB & JFI ; 
 QPC <= QAB & JFJ ; 
 QPD <= QAB & GBK ; 
 PBC <=  PBC & jhc & tpc  |  pbc & JHC  |  ABC & TPC  ; 
 PDC <=  PBC & jhc & tpc  |  pbc & JHC  |  ABC & TPC  ; 
 PFC <=  PBC & jhc & tpc  |  pbc & JHC  |  ABC & TPC  ; 
 QUA <=  qpb & QPA  ; 
 QUF <=  JPA & QPA  |  QPB  |  QUE  ; 
 BBC <=  BBC & jec & tfc  |  bbc & JEC  |  ABC & TFC  ; 
 BDC <=  BBC & jec & tfc  |  bbc & JEC  |  ABC & TFC  ; 
 BFC <=  BBC & jec & tfc  |  bbc & JEC  |  ABC & TFC  ; 
 QUD <=  QUC  |  QPC  ; 
 PBK <=  PBK & jhk & tpd  |  pbk & JHK  |  ABK & TPD  ; 
 PDK <=  PBK & jhk & tpd  |  pbk & JHK  |  ABK & TPD  ; 
 PFK <=  PBK & jhk & tpd  |  pbk & JHK  |  ABK & TPD  ; 
 BBK <=  BBK & jek & tfd  |  bbk & JEK  |  ABK & TFD  ; 
 BDK <=  BBK & jek & tfd  |  bbk & JEK  |  ABK & TFD  ; 
 BFK <=  BBK & jek & tfd  |  bbk & JEK  |  ABK & TFD  ; 
 RMA <= JKB ; 
 RMC <= RMB ; 
 RMD <= RMC ; 
 RNM <= RNL ; 
 RNN <= RNM ; 
 RNO <= RNN ; 
 RNP <= RNO ; 
 RNA <=  JKB & QHD  |  RME  ; 
 RNK <=  RMJ & QHD  ; 
 RMN <=  RMM & jjg  ; 
 RMG <= RMF ; 
 RMH <= RMG ; 
 RMI <= RMH ; 
 RMJ <= RMI ; 
 RMK <=  RMJ & qhd  |  RMU  ; 
 RME <=  RKA & jic & jid  |  RMD  ; 
 RML <= RMK ; 
 RMM <= RML ; 
 RMO <= RMN ; 
 RMP <= RMO ; 
 RNB <= RNA ; 
 RNC <= RNB ; 
 RND <= RNC ; 
 RNL <= RNK ; 
 RMR <=  RMQ & QRA  ; 
 RMF <=  RME & QRA  |  RNP  ; 
 RMQ <= RMP ; 
 RMS <= RMR ; 
 RMT <= RMS ; 
 RMU <= RMT ; 
 RMB <=  RMQ & qra  |  RMA  ; 
 LBC <=  LBC & jlc & tla  |  lbc & JLC  |  LAC & TLA  ; 
 AGH <= AEH ; 
 AGI <= AEI ; 
 AGJ <= AEJ ; 
 AGK <= AEK ; 
 ack <= wck & QKR |  aqk & qkr ; 
 adc <= wdc & QKR |  arc & qkr ; 
 adk <= wdk & QKR |  ark & qkr ; 
 AGL <= AEL ; 
 AGM <= AEM ; 
 AGN <= AEN ; 
 AGO <= AEO ; 
 CEA <=  BID  |  ZZI & BIB  |  BIA  |  ZZO & ZZI  |  BIC  ; 
 AGP <= AEP ; 
 AHA <= AFA ; 
 AHB <= AFB ; 
 AHC <= AFC ; 
 CEB <=  BIH  |  BIE  |  BIF  |  ZZO & ZZI  |  BIG  ; 
 AHD <= AFD ; 
 AHE <= AFE ; 
 AHF <= AFF ; 
 AHG <= AFG ; 
 AHH <= AFH ; 
 AHI <= AFI ; 
 AHJ <= AFJ ; 
 AHK <= AFK ; 
 gac <= fac & TGA |  jac & tga ; 
 gck <= eac & TGA |  gck & tga ; 
 GAE <= FAB & TGA |  GAE & tga ; 
 AHL <= AFL ; 
 AHM <= AFM ; 
 AHN <= AFN ; 
 AHO <= AFO ; 
 gag <=  eag & TGF  |  ZZO & TGF  |  gag & tgf  ; 
 gch <=  faa & TGF  |  fba & TGF  |  gch & tgf  ; 
 gal <=  TGB & fad  |  fap & TGD  |  gal & tgb  ; 
 gan <=  TGB & fad  |  fbe & TGD  |  gan & tgb  ; 
 gbc <=  faa & TGF  |  fal & TGF  |  gbc & tgf  ; 
 gbd <=  faa & TGF  |  fbc & TGF  |  gbd & tgf  ; 
 gbg <=  fag & TGC  |  fbe & TGE  |  gbg & tgc  ; 
 gba <=  faa & TGC  |  fak & TGE  |  gba & tgc  ; 
 gbk <=  faf & TGF  |  fal & TGF  |  gbk & tgf  ; 
 gbf <=  faf & TGF  |  FBE & TGF  |  gbf & tgf  ; 
 QKB <=  QKB & jaq  |  JCI & QAA  ; 
 HFM <= HEH & HEA ; 
 HFN <= HEH & HEB ; 
 QKA <=  QKA & qkk  |  GAL & QAA  ; 
 MAA <= MAA & tld |  GAG & TLD ; 
 MAB <= MAB & tld |  GAH & TLD ; 
 MAC <= MAC & tld |  GAI & TLD ; 
 AAC <=  IAC & TAA  |  DAC & TBA  |  IEC & TCA  |  WAC & TDA  |  TMA  ; 
 OHA <=  IAC & TAA  |  DAC & TBA  |  IEC & TCA  |  WAC & TDA  |  TMA  ; 
 OAC <=  DAC & TEA  |  EAC & TEC  |  NAC & TEE  ; 
 OAK <=  DAK & TEA  |  ECK & TEC  |  WCM & TEE  ; 
 ASK <=  IAK & TAB  |  DAK & TBB  |  IEK & TCB  |  WAK & TDB  |  TMB  ; 
 AAK <=  IAK & TAB  |  DAK & TBB  |  IEK & TCB  |  WAK & TDB  |  TMB  ; 
 ATC <=  IBC & TAC  |  DBC & TBC  |  EAC & TCC  |  WBC & TDC  |  TMC  ; 
 ABC <=  IBC & TAC  |  DBC & TBC  |  EAC & TCC  |  WBC & TDC  |  TMC  ; 
 DAC <= ICC ; 
 DAK <= ICK ; 
 DBC <= IDC ; 
 DBK <= IDK ; 
 orc <= gck ; 
 EDC <= EAC ; 
 QZF <= QZE ; 
 ATK <=  IBK & TAD  |  DBK & TBD  |  ECK & TCD  |  WBK & TDD  |  TMD  ; 
 ABK <=  IBK & TAD  |  DBK & TBD  |  ECK & TCD  |  WBK & TDD  |  TMD  ; 
 OBC <=  DBC & TEB  |  EDC & TED  |  WDE & TEF  ; 
 OBK <=  DBK & TEB  |  EDK & TED  |  WDM & TEF  ; 
 ebk <= iek ; 
 eak <= iek ; 
 eac <= iec ; 
 eck <= iek ; 
 NAC <=  NAC & jsc & tha  |  nac & JSC  |  WCE & THA  ; 
 NBC <=  NAC & jsc & tha  |  nac & JSC  |  WCE & THA  ; 
 occ <= pcc ; 
 ock <= pck ; 
 odc <= pdc ; 
 odk <= pdk ; 
 QGB <=  ife  |  ifff   |  ifg  |  ifh  ; 
 QKC <=  JAA  |  QKC & jaq  ; 
 QFA <= IMG ; 
 rmv <= rmh ; 
 RAG <= JBG ; 
 OKA <=  IKA & jbc  |  IKA & qkk  |  JBC & QKB  ; 
 OEC <= KAC ; 
 EDK <= ECK ; 
 KAC <=  KAC & tlc  |  MAA & QMG  |  JNC  ; 
 KAE <=  KAE & tlc  |  MAC & QMG  |  JNE  ; 
 QKD <=  IKA & JBC  |  IKB & JBD  ; 
 QKE <=  QKB & JBC  |  QKB & JBD  ; 
 OKB <=  IKB & jbd  |  IKB & qkk  |  JBD & QKB  ; 
 LAC <=  IPC & tlb & jcr  |  IQC & TLB  ; 
 PAD <=  PAD & jgd & tpa  |  pad & JGD  |  AAD & TPA  ; 
 PCD <=  PAD & jgd & tpa  |  pad & JGD  |  AAD & TPA  ; 
 PED <=  PAD & jgd & tpa  |  pad & JGD  |  AAD & TPA  ; 
 PAL <=  PAL & jgl & tpb  |  pal & JGL  |  AAL & TPB  ; 
 PCL <=  PAL & jgl & tpb  |  pal & JGL  |  AAL & TPB  ; 
 PEL <=  PAL & jgl & tpb  |  pal & JGL  |  AAL & TPB  ; 
 BAL <=  BAL & jdl & tfb  |  bal & JDL  |  AAL & TFB  ; 
 BEL <=  BAL & jdl & tfb  |  bal & JDL  |  AAL & TFB  ; 
 QWB <= QWA ; 
 QWC <= QWB ; 
 qwi <= jdf ; 
 qwd <= jda ; 
 PBD <=  PBD & jhd & tpc  |  pbd & JHD  |  ABD & TPC  ; 
 PDD <=  PBD & jhd & tpc  |  pbd & JHD  |  ABD & TPC  ; 
 PFD <=  PBD & jhd & tpc  |  pbd & JHD  |  ABD & TPC  ; 
 BBD <=  BBD & jed & tfc  |  bbd & JED  |  ABD & TFC  ; 
 BFD <=  BBD & jed & tfc  |  bbd & JED  |  ABD & TFC  ; 
 QWA <=  QKJ  ; 
 QWJ <=  QKJ  |  QZF  ; 
 PBL <=  PBL & jhl & tpd  |  pbl & JHL  |  ABL & TPD  ; 
 PDL <=  PBL & jhl & tpd  |  pbl & JHL  |  ABL & TPD  ; 
 PFL <=  PBL & jhl & tpd  |  pbl & JHL  |  ABL & TPD  ; 
 BBL <=  BBL & jel & tfd  |  bbl & JEL  |  ABL & TFD  ; 
 BFL <=  BBL & jel & tfd  |  bbl & JEL  |  ABL & TFD  ; 
 QLL <=  QLL & qlm  |  RKD & rmg  ; 
 RKB <= RKA ; 
 RKC <= RKB ; 
 RKD <= RKC ; 
 RLB <= RLA ; 
 RLD <=  ZZO & qqh  |  ZZO & QAC  |  RLC  ; 
 RLA <=  QLD & qlk  |  JFX & QAC  |  JJH & qrc  ; 
 QLM <=  QLL & jic & jid  ; 
 QLA <= JRC ; 
 QLB <= QLA ; 
 QLC <= QLB ; 
 RLC <= RLB ; 
 QLF <=  QLF & jjg  |  JCK & QAC  |  RSA  ; 
 QLG <=  QLG & jjg  |  ZZO & QAC  |  RKA  ; 
 QLD <=  JKA & qrb & qlo  |  QLC  ; 
 QLN <=  RML & rha  |  QLF & QLK  |  QTP  ; 
 QLO <=  RML & rha  |  QLF & QLK  |  QTP  ; 
 QLI <=  QLI & jjg  |  ZZO & QLD  |  QLJ  ; 
 QLK <=  QLK & jjg  |  JLG & QLD  ; 
 LBD <=  LBD & jld & tla  |  lbd & JLD  |  LAD & TLA  ; 
 AIH <= AGH ; 
 AII <= AGI ; 
 AIJ <= AGJ ; 
 AIK <= AGK ; 
 acl <= wcl & QKR |  aql & qkr ; 
 add <= wdd & QKR |  ard & qkr ; 
 adl <= wdl & QKR |  arl & qkr ; 
 AIL <= AGL ; 
 AIM <= AGM ; 
 AIN <= AGN ; 
 AIO <= AGO ; 
 CFA <=  BJD  |  ZZI & BJB  |  BJA  |  ZZO & ZZI  |  BJC  ; 
 AIP <= AGP ; 
 AJA <= AHA ; 
 AJB <= AHB ; 
 AJC <= AHC ; 
 CFB <=  BJH  |  BJE  |  BJF  |  ZZO & ZZI  |  BJG  ; 
 AJD <= AHD ; 
 AJE <= AHE ; 
 AJF <= AHF ; 
 AJG <= AHG ; 
 AJH <= AHH ; 
 AJI <= AHI ; 
 AJJ <= AHJ ; 
 AJK <= AHK ; 
 gcl <= ead & TGA |  gcl & tga ; 
 gah <= eah & TGA |  gah & tga ; 
 gaf <= fag & TGA |  jfx & tga ; 
 AJL <= AHL ; 
 AJM <= AHM ; 
 AJN <= AHN ; 
 AJO <= AHO ; 
 gca <=  TGB & fag  |  fba & TGD  |  gca & tgb  ; 
 gcb <=  TGB & fag  |  fbb & TGD  |  gcb & tgb  ; 
 QLP <=  QLP & jqa  |  JCL & QAC  |  JXB  |  JQB & JCQ  ; 
 QLQ <=  QLP & jqa  |  JCL & QAC  |  JXB  |  JQB & JCQ  ; 
 gcc <=  TGC & fag  |  fbc & TGE  |  gcc & tgc  ; 
 gcd <=  TGC & fag  |  fbd & TGE  |  gcd & tgc  ; 
 RKA <= QAC & GBO ; 
 QLJ <= QAC & GBP ; 
 QRB <= QRA ; 
 QRC <= QRB ; 
 QRD <= QRC ; 
 QRE <= QRD ; 
 qna <=  qac  |  jfx  ; 
 qne <=  qac  |  jfx  |  GAA  ; 
 AAD <=  IAD & TAA  |  DAD & TBA  |  IED & TCA  |  WAD & TDA  |  TMA  ; 
 OHB <=  IAD & TAA  |  DAD & TBA  |  IED & TCA  |  WAD & TDA  |  TMA  ; 
 OAD <=  DAD & TEA  |  EAD & TEC  |  NAD & TEE  ; 
 OAL <=  DAL & TEA  |  ECL & TEC  |  WCN & TEE  ; 
 ASL <=  IAL & TAB  |  DAL & TBB  |  IEL & TCB  |  WAL & TDB  |  TMB  ; 
 AAL <=  IAL & TAB  |  DAL & TBB  |  IEL & TCB  |  WAL & TDB  |  TMB  ; 
 ATD <=  IBD & TAC  |  DBD & TBC  |  EAD & TCC  |  WBD & TDC  |  TMC  ; 
 ABD <=  IBD & TAC  |  DBD & TBC  |  EAD & TCC  |  WBD & TDC  |  TMC  ; 
 DAD <= ICD ; 
 DAL <= ICL ; 
 DBD <= IDD ; 
 DBL <= IDL ; 
 ord <= gcl ; 
 EDD <= EAD ; 
 EDL <= ECL ; 
 RJL <= JJC ; 
 ATL <=  IBL & TAD  |  DBL & TBD  |  ECL & TCD  |  WBL & TDD  |  TMD  ; 
 ABL <=  IBL & TAD  |  DBL & TBD  |  ECL & TCD  |  WBL & TDD  |  TMD  ; 
 OBD <=  DBD & TEB  |  EDD & TED  |  WDF & TEF  ; 
 OBL <=  DBL & TEB  |  EDL & TED  |  WDN & TEF  ; 
 ebl <= iel ; 
 eal <= iel ; 
 ead <= ied ; 
 ecl <= iel ; 
 NAD <=  NAD & jsd & tha  |  nad & JSD  |  WCF & THA  ; 
 NBD <=  NAD & jsd & tha  |  nad & JSD  |  WCF & THA  ; 
 QFB <=  QFB & QLS  |  QFA & qls  ; 
 OLF <=  QFB & QLS  |  QFA & qls  ; 
 ocd <= pcd ; 
 ocl <= pcl ; 
 odd <= pdd ; 
 odl <= pdl ; 
 QNI <= JAG & GCA ; 
 QNM <= JAG & GCB ; 
 QNQ <= JAG & GCC ; 
 QNU <= JAG & GCD ; 
 QRA <=  RIX  |  JRA  |  QHF  |  IJD  ; 
 OJC <=  JRF  |  JRA  |  IHB & jcd  |  JRE  |  IJD  ; 
 OMA <=  QLG & jrc  |  JRB  |  JRD  |  IJD  ; 
 OMB <=  QLG & jrc  |  JRB  |  JRD  |  IJD  ; 
 QLR <= QLQ ; 
 QLS <= QLR ; 
 RJC <= RJB ; 
 RIX <= JRB ; 
 OJD <=  JCA  |  JJB  |  JCN  |  QQC  ; 
 OED <=  KAD  ; 
 oei <=  qfc  |  QSG  ; 
 KAD <=  KAD & tlc  |  MAB & QMG  |  JND  |  RSC & QSB  ; 
 qib <= qia ; 
 qic <= qib ; 
 qid <= qic ; 
 OTC <= QLQ ; 
 qia <=  ijd & qhf  |  ijd & QRA  ; 
 LAD <=  IPD & tlb & jcr  |  IQD & TLB  ; 
 PAE <=  PAE & jge & tpa  |  pae & JGE  |  AAE & TPA  ; 
 PCE <=  PAE & jge & tpa  |  pae & JGE  |  AAE & TPA  ; 
 PEE <=  PAE & jge & tpa  |  pae & JGE  |  AAE & TPA  ; 
 PAM <=  PAM & jgm & tpb  |  pam & JGM  |  AAM & TPB  ; 
 PCM <=  PAM & jgm & tpb  |  pam & JGM  |  AAM & TPB  ; 
 PEM <=  PAM & jgm & tpb  |  pam & JGM  |  AAM & TPB  ; 
 qvc <=  quf  |  jfa  ; 
 qvd <=  quf  |  jfa  |  jfb  ; 
 BAM <=  BAM & jdm & tfb  |  bam & JDM  |  AAM & TFB  ; 
 BCM <=  BAM & jdm & tfb  |  bam & JDM  |  AAM & TFB  ; 
 BEM <=  BAM & jdm & tfb  |  bam & JDM  |  AAM & TFB  ; 
 qwh <=  jda  |  jdb  |  jdc  |  jdd  |  jde  ; 
 PBE <=  PBE & jhe & tpc  |  pbe & JHE  |  ABE & TPC  ; 
 PDE <=  PBE & jhe & tpc  |  pbe & JHE  |  ABE & TPC  ; 
 PFE <=  PBE & jhe & tpc  |  pbe & JHE  |  ABE & TPC  ; 
 BBE <=  BBE & jee & tfc  |  bbe & JEE  |  ABE & TFC  ; 
 BDE <=  BBE & jee & tfc  |  bbe & JEE  |  ABE & TFC  ; 
 BFE <=  BBE & jee & tfc  |  bbe & JEE  |  ABE & TFC  ; 
 PBM <=  PBM & jhm & tpd  |  pbm & JHM  |  ABM & TPD  ; 
 PDM <=  PBM & jhm & tpd  |  pbm & JHM  |  ABM & TPD  ; 
 BBM <=  BBM & jem & tfd  |  bbm & JEM  |  ABM & TFD  ; 
 BDM <=  BBM & jem & tfd  |  bbm & JEM  |  ABM & TFD  ; 
 RBX <=  RBX & jcx & jcc  |  RBB  ; 
 qnj <= qni ; 
 qnn <= qnm ; 
 qnr <= qnq ; 
 qnv <= qnu ; 
 QMK <=  QMK & qln  |  QMJ  ; 
 QML <=  QMK & qln  |  QMJ  ; 
 LBE <=  LBE & jle & tla  |  lbe & JLE  |  LAE & TLA  ; 
 AKH <= AIH ; 
 AKI <= AII ; 
 AKJ <= AIJ ; 
 AKK <= AIK ; 
 acm <= wcm & QKR |  aqm & qkr ; 
 ade <= wde & QKR |  are & qkr ; 
 adm <= wdm & QKR |  arm & qkr ; 
 AKL <= AIL ; 
 AKM <= AIM ; 
 AKN <= AIN ; 
 AKO <= AIO ; 
 CGA <=  BKD  |  ZZI & BKB  |  BKA  |  ZZO & ZZI  |  BKC  ; 
 AKP <= AIP ; 
 ALA <= AJA ; 
 ALB <= AJB ; 
 ALC <= AJC ; 
 CGB <=  BKH  |  BKE  |  BKF  |  ZZO & ZZI  |  BKG  ; 
 ALD <= AJD ; 
 ALE <= AJE ; 
 ALF <= AJF ; 
 ALG <= AJG ; 
 ALH <= AJH ; 
 ALI <= AJI ; 
 ALJ <= AJJ ; 
 ALK <= AJK ; 
 gcm <= eae & TGA |  gcm & tga ; 
 gcj <= eab & TGA |  gcj & tga ; 
 gcn <= eaf & TGA |  gcn & tga ; 
 ALL <= AJL ; 
 ALM <= AJM ; 
 ALN <= AJN ; 
 ALO <= AJO ; 
 RBB <= jcd & RBA ; 
 RBC <= jcd & RBB ; 
 RBD <= jcd & RBC ; 
 RBE <= jcd & JOX ; 
 gbn <=  TGB & fah  |  faj & TGD  |  gbn & tgb  ; 
 gbm <=  TGB & fah  |  fai & TGD  |  gbm & tgb  ; 
 gap <=  fab & TGC  |  fbe & TGE  |  gap & tgc  ; 
 gbo <=  fah & TGC  |  fak & TGE  |  gbo & tgc  ; 
 QLE <=  JJE & RLB  |  JKA & qrb  |  QLC  ; 
 RAF <=  ZZO & RLB  |  ZZO & qrb  |  JCM  ; 
 QKO <=  GAP & gab & JAG  |  QKO & raf  ; 
 QKS <=  GAP & gab & JAG  |  QKO & raf  ; 
 RAB <= RAA ; 
 RAC <= RAB ; 
 RAD <= RAC ; 
 RAE <= RAD ; 
 QCX <=  QCY & jco & rat  |  QCD & qck  |  QCH  ; 
 QCZ <=  QCY & jco & rat  |  QCD & qck  |  QCH  ; 
 QCY <=  QCY & jco & rat  |  QCD & qck  |  QCH  ; 
 AAE <=  IAE & TAA  |  DAE & TBA  |  IEE & TCA  |  WAE & TDA  |  TMA  ; 
 OHC <=  IAE & TAA  |  DAE & TBA  |  IEE & TCA  |  WAE & TDA  |  TMA  ; 
 OAE <=  DAE & TEA  |  EAE & TEC  |  NAE & TEE  ; 
 OAM <=  DAM & TEA  |  ECM & TEC  |  WCO & TEE  ; 
 ASM <=  IAM & TAB  |  DAM & TBB  |  IEM & TCB  |  WAM & TDB  |  TMB  ; 
 AAM <=  IAM & TAB  |  DAM & TBB  |  IEM & TCB  |  WAM & TDB  |  TMB  ; 
 QXA <=  REC  |  RAA  |  QZE  |  JCF  ; 
 QXB <=  REC  |  RAA  |  QZE  |  JCF  ; 
 ATE <=  IBE & TAC  |  DBE & TBC  |  EAE & TCC  |  WBE & TDC  |  TMC  ; 
 ABE <=  IBE & TAC  |  DBE & TBC  |  EAE & TCC  |  WBE & TDC  |  TMC  ; 
 DAE <= ICE ; 
 DAM <= ICM ; 
 DBE <= IDE ; 
 DBM <= IDM ; 
 ore <= gcm ; 
 EDE <= EAE ; 
 EDM <= ECM ; 
 oig <= qxe ; 
 ATM <=  IBM & TAD  |  DBM & TBD  |  ECM & TCD  |  WBM & TDD  |  TMD  ; 
 ABM <=  IBM & TAD  |  DBM & TBD  |  ECM & TCD  |  WBM & TDD  |  TMD  ; 
 OBE <=  DBE & TEB  |  EDE & TED  |  WDG & TEF  ; 
 OBM <=  DBM & TEB  |  EDM & TED  |  WDO & TEF  ; 
 eae <= iee ; 
 eam <= iem ; 
 ecm <= iem ; 
 eao <= ieo ; 
 REC <=  JCA  |  JCG  |  JCB  |  JCM  ; 
 OIA <=  JCA  |  JCG  |  JCB  |  JCM  ; 
 oce <= pce ; 
 ocm <= pcm ; 
 ode <= pde ; 
 odm <= pdm ; 
 OIC <=  JBB & QCY  |  ifi & JAO  |  IFI & JAP  |  JAM  |  JAN  ; 
 QQZ <=  JBB & QCY  |  ifi & JAO  |  IFI & JAP  |  JAM  |  JAN  ; 
 OID <= QQQ & QCI ; 
 QQO <= QQQ & QQH ; 
 QCI <= QQQ & QQH ; 
 QKW <= QQQ & QCI ; 
 OIE <=  jbb & JCW  |  jbe & RAF  |  IFI & HEO  |  ifi & HEP  ; 
 QKY <=  jbb & JCW  |  jbe & RAF  |  IFI & HEO  |  ifi & HEP  ; 
 OEE <= KAE ; 
 QRF <= QRE ; 
 OLC <= QTX ; 
 OTA <= QTX ; 
 qmb <= qma ; 
 qmc <= qmb ; 
 qmf <= qme ; 
 qmg <= qmf ; 
 otd <= qrf ; 
 qmj <= qmi ; 
 oib <= rab ; 
 qck <= qcj ; 
 LAE <=  IPE & tlb & jcr  |  IQE & TLB  ; 
 PAF <=  PAF & jgf & tpa  |  paf & JGF  |  AAF & TPA  ; 
 PCF <=  PAF & jgf & tpa  |  paf & JGF  |  AAF & TPA  ; 
 PEF <=  PAF & jgf & tpa  |  paf & JGF  |  AAF & TPA  ; 
 PAN <=  PAN & jgn & tpb  |  pan & JGN  |  AAN & TPB  ; 
 PCN <=  PAN & jgn & tpb  |  pan & JGN  |  AAN & TPB  ; 
 PEN <=  PAN & jgn & tpb  |  pan & JGN  |  AAN & TPB  ; 
 BAN <=  BAN & jdn & tfb  |  ban & JDN  |  AAN & TFB  ; 
 BCN <=  BAN & jdn & tfb  |  ban & JDN  |  AAN & TFB  ; 
 BEN <=  BAN & jdn & tfb  |  ban & JDN  |  AAN & TFB  ; 
 qwf <=  jda  |  jdb  |  jdc  ; 
 qwe <=  jda  |  jdb  ; 
 PBF <=  PBF & jhf & tpc  |  pbf & JHF  |  ABF & TPC  ; 
 PDF <=  PBF & jhf & tpc  |  pbf & JHF  |  ABF & TPC  ; 
 PFF <=  PBF & jhf & tpc  |  pbf & JHF  |  ABF & TPC  ; 
 BBF <=  BBF & jef & tfc  |  bbf & JEF  |  ABF & TFC  ; 
 BDF <=  BBF & jef & tfc  |  bbf & JEF  |  ABF & TFC  ; 
 BFF <=  BBF & jef & tfc  |  bbf & JEF  |  ABF & TFC  ; 
 PBN <=  PBN & jhn & tpd  |  pbn & JHN  |  ABN & TPD  ; 
 PDN <=  PBN & jhn & tpd  |  pbn & JHN  |  ABN & TPD  ; 
 BBN <=  BBN & jen & tfd  |  bbn & JEN  |  ABN & TFD  ; 
 BDN <=  BBN & jen & tfd  |  bbn & JEN  |  ABN & TFD  ; 
 HIA <= GDA ; 
 HIB <= GDB ; 
 HIC <= GDC ; 
 HKA <= HJA ; 
 HKB <= HJB ; 
 HKC <= HJC ; 
 QQC <=  QQC & qqr & jjp  |  JQC & JQE  ; 
 QQP <=  QQC & qqr & jjp  |  JQC & JQE  ; 
 QQQ <=  QQC & qqr & jjp  |  JQC & JQE  ; 
 HJA <= HIA ; 
 HJB <= HIB ; 
 HJC <= HIC ; 
 HLA <= HKA ; 
 HLB <= HKB ; 
 HLC <= HKC ; 
 HMA <= HLA ; 
 HMB <= HLB ; 
 HMC <= HLC ; 
 GDY <= GDX ; 
 LBF <=  LBF & jlf & tla  |  lbf & JLF  |  LAF & TLA  ; 
 AMH <= AKH ; 
 AMI <= AKI ; 
 AMJ <= AKJ ; 
 AMK <= AKK ; 
 acn <= wcn & QKR |  aqn & qkr ; 
 adf <= wdf & QKR |  arf & qkr ; 
 adn <= wdn & QKR |  arn & qkr ; 
 AML <= AKL ; 
 AMM <= AKM ; 
 AMN <= AKN ; 
 AMO <= AKO ; 
 CHA <=  BLD  |  ZZI & BLB  |  BLA  |  ZZO & ZZI  |  BLC  ; 
 AMP <= AKP ; 
 ANA <= ALA ; 
 ANB <= ALB ; 
 ANC <= ALC ; 
 CHB <=  BLH  |  BLE  |  BLF  |  ZZO & ZZI  |  BLG  ; 
 ANDD  <= ALD ; 
 ANE <= ALE ; 
 ANF <= ALF ; 
 ANG <= ALG ; 
 ANH <= ALH ; 
 ANI <= ALI ; 
 ANJ <= ALJ ; 
 ANK <= ALK ; 
 ANL <= ALL ; 
 ANM <= ALM ; 
 ANN <= ALN ; 
 ANO <= ALO ; 
 QQB <=  JQF & jjp & ihc  |  JQC & JQE  ; 
 QQW <=  JQF & jjp & ihc  |  JQC & JQE  ; 
 QQD <= QQC ; 
 QQE <= QQD ; 
 QQF <= JJE ; 
 QQG <= QQF ; 
 QHE <= QHD ; 
 QHF <= QHE ; 
 qtq <= qtp ; 
 qtr <= qtp ; 
 RLX <=  RLX & jfy  |  GAF & QAA  |  IHB  ; 
 AAF <=  IAF & TAA  |  DAF & TBA  |  IEF & TCA  |  WAF & TDA  |  TMA  ; 
 OHD <=  IAF & TAA  |  DAF & TBA  |  IEF & TCA  |  WAF & TDA  |  TMA  ; 
 OAF <=  DAF & TEA  |  EAF & TEC  |  WCH & TEE  ; 
 OAN <=  DAN & TEA  |  ECN & TEC  |  WCP & TEE  ; 
 ASN <=  IAN & TAB  |  DAN & TBB  |  IEN & TCB  |  WAN & TDB  |  TMB  ; 
 AAN <=  IAN & TAB  |  DAN & TBB  |  IEN & TCB  |  WAN & TDB  |  TMB  ; 
 QXC <=  REC  |  RAA  |  QZE  |  JCF  ; 
 QXD <=  REC  |  RAA  |  QZE  |  JCF  ; 
 ATF <=  IBF & TAC  |  DBF & TBC  |  EAF & TCC  |  WBF & TDC  |  TMC  ; 
 ABF <=  IBF & TAC  |  DBF & TBC  |  EAF & TCC  |  WBF & TDC  |  TMC  ; 
 DAF <= ICF ; 
 DAN <= ICN ; 
 DBF <= IDF ; 
 DBN <= IDN ; 
 orf <= gcn ; 
 EDF <= EAF ; 
 EDN <= ECN ; 
 ATN <=  IBN & TAD  |  DBN & TBD  |  ECN & TCD  |  WBN & TDD  |  TMD  ; 
 ABN <=  IBN & TAD  |  DBN & TBD  |  ECN & TCD  |  WBN & TDD  |  TMD  ; 
 OBF <=  DBF & TEB  |  EDF & TED  |  WDH & TEF  ; 
 OBN <=  DBN & TEB  |  EDN & TED  |  WDP & TEF  ; 
 eaf <= ief ; 
 QBA <= IJC ; 
 ean <= ien ; 
 ecn <= ien ; 
 NAE <=  NAE & jse & tha  |  nae & JSE  |  WCG & THA  ; 
 rba <=  ihb  |  JCB  |  JCD  |  JCH  ; 
 ocf <= pcf ; 
 ocn <= pcn ; 
 odf <= pdf ; 
 odn <= pdn ; 
 OGA <=  HIA & JOA  |  HJA & JOB  |  HKA & JOC  |  HLA & JOD  |  GDJ  ; 
 OGB <=  HIB & JOA  |  HJB & JOB  |  HKB & JOC  |  HLB & JOD  |  GDK  ; 
 QHC <=  IOA  |  IOB  |  IOC  |  IOD  ; 
 QHD <=  IOA & RMV  |  IOB & RMV  |  IOC & RMV  |  IOD & RMV  |  RMN  ; 
 OEJ <=  IOA & RMV  |  IOB & RMV  |  IOC & RMV  |  IOD & RMV  |  RMN  ; 
 OGC <=  HIC & JOA  |  HJC & JOB  |  HKC & JOC  |  HLC & JOD  |  GDL  ; 
 OGD <=  JOA & JOJ  |  JOB & JOJ  |  JOC & JOJ  |  JOD & JOJ  |  QCJ  ; 
 QCD <=  JOA & JOJ  |  JOB & JOJ  |  JOC & JOJ  |  JOD & JOJ  |  QCJ  ; 
 OEM <=  QML  |  QNN  |  QNR  |  QSE  ; 
 OEF <= KAF ; 
 ote <= qqf ; 
 QQY <= QQT ; 
 GDX <= IHC ; 
 OGI <=  JOA & JOO  |  JOB & JOO  |  JOC & JOO  |  JOD & JOO  |  QCJ  ; 
 QQT <=  IHB & jce  |  JOX & jjh  |  QQA & jjl  |  JIA  ; 
 QQA <=  IHB & jce  |  JOX & jjh  |  QQA & jjl  |  JIA  ; 
 OEP <=  QMK  |  QNB  |  QSE  |  JCS  ; 
 LAF <=  IPF & tlb & jcr  |  IQF & TLB  |  JCR  ; 
 PAG <=  PAG & jgg & tpa  |  pag & JGG  |  AAG & TPA  ; 
 PCG <=  PAG & jgg & tpa  |  pag & JGG  |  AAG & TPA  ; 
 PEG <=  PAG & jgg & tpa  |  pag & JGG  |  AAG & TPA  ; 
 PAO <=  PAO & jgo & tpb  |  pao & JGO  |  AAO & TPB  ; 
 PCO <=  PAO & jgo & tpb  |  pao & JGO  |  AAO & TPB  ; 
 PEO <=  PAO & jgo & tpb  |  pao & JGO  |  AAO & TPB  ; 
 qve <=  quf  |  jfa  |  jfb  |  jfc  ; 
 BAO <=  BAO & jdo & tfb  |  bao & JDO  |  AAO & TFB  ; 
 BCO <=  BAO & jdo & tfb  |  bao & JDO  |  AAO & TFB  ; 
 BEO <=  BAO & jdo & tfb  |  bao & JDO  |  AAO & TFB  ; 
 qwg <=  jda  |  jdb  |  jdc  |  jdd  ; 
 PBG <=  PBG & jhg & tpc  |  pbg & JHG  |  ABG & TPC  ; 
 PDG <=  PBG & jhg & tpc  |  pbg & JHG  |  ABG & TPC  ; 
 PFG <=  PBG & jhg & tpc  |  pbg & JHG  |  ABG & TPC  ; 
 BBG <=  BBG & jeg & tfc  |  bbg & JEG  |  ABG & TFC  ; 
 BDG <=  BBG & jeg & tfc  |  bbg & JEG  |  ABG & TFC  ; 
 BFG <=  BBG & jeg & tfc  |  bbg & JEG  |  ABG & TFC  ; 
 PBO <=  PBO & jho & tpd  |  pbo & JHO  |  ABO & TPD  ; 
 PDO <=  PBO & jho & tpd  |  pbo & JHO  |  ABO & TPD  ; 
 BBO <=  BBO & jeo & tfd  |  bbo & JEO  |  ABO & TFD  ; 
 BDO <=  BBO & jeo & tfd  |  bbo & JEO  |  ABO & TFD  ; 
 GDA <=  gda & gda  |  TME  ; 
 GDB <=  GDB & gda  |  TME  |  gdb & GDA  ; 
 GDD <=  GDD & tme & jva  |  JVA & gdd  ; 
 GDG <=  GDD & tme & jva  |  JVA & gdd  ; 
 GDE <=  GDE & tme & jvb  |  JVB & gde  ; 
 GDH <=  GDE & tme & jvb  |  JVB & gde  ; 
 GDC <=  GDC & jua  |  gdc & JUA  |  TME  ; 
 GDF <=  GDF & tme & jvc  |  JVC & gdf  ; 
 GDI <=  GDF & tme & jvc  |  JVC & gdf  ; 
 QKP <=  jvd & QKP  |  QQO  ; 
 QKQ <=  JVD & QKP  ; 
 QTF <= QTE ; 
 QTG <= QTF ; 
 QTH <= QTG ; 
 QTI <= QTH ; 
 AOH <= AMH ; 
 AOI <= AMI ; 
 AOJ <= AMJ ; 
 AOK <= AMK ; 
 aco <= wco & QKR |  aqo & qkr ; 
 ado <= wdo & QKR |  aro & qkr ; 
 adg <= wdg & QKR |  arg & qkr ; 
 AOL <= AML ; 
 AOM <= AMM ; 
 AON <= AMN ; 
 AOO <= AMO ; 
 CIA <=  BMD  |  ZZI & BMB  |  BMA  |  ZZO & ZZI  |  BMC  ; 
 AOP <= AMP ; 
 APA <= ANA ; 
 APB <= ANB ; 
 APC <= ANC ; 
 CIB <=  BMH  |  BME  |  BMF  |  ZZO & ZZI  |  BMG  ; 
 APD <= ANDD  ; 
 APE <= ANE ; 
 APF <= ANF ; 
 APG <= ANG ; 
 APH <= ANH ; 
 API <= ANI ; 
 APJ <= ANJ ; 
 APK <= ANK ; 
 APL <= ANL ; 
 APM <= ANM ; 
 APN <= ANN ; 
 APO <= ANO ; 
 RAX <=  RAX & jcu  |  RAA  |  RJA  ; 
 raa <= jia & ZZI ; 
 rat <= jia & ZZI ; 
 qtb <= qta ; 
 QTC <= QTB ; 
 QTD <= QTC ; 
 QTE <= QTD ; 
 QKR <=  QKQ  |  TME  ; 
 qnb <= qna ; 
 qnc <= qnb ; 
 qnf <= qne ; 
 qng <= qnf ; 
 QMA <= QAC & JCL ; 
 QME <= QAC & JCJ ; 
 QMI <= QAC & JFH ; 
 RQB <= RQA ; 
 rqc <= rqb ; 
 AAG <=  IAG & TAA  |  DAG & TBA  |  IEG & TCA  |  WAG & TDA  |  TMA  ; 
 OHE <=  IAG & TAA  |  DAG & TBA  |  IEG & TCA  |  WAG & TDA  |  TMA  ; 
 OAG <=  DAG & TEA  |  EAG & TEC  |  WCI & TEE  ; 
 OAO <=  DAO & TEA  |  ECO & TEC  |  WDA & TEE  ; 
 ASO <=  IAO & TAB  |  DAO & TBB  |  IEO & TCB  |  WAO & TDB  |  TMB  ; 
 AAO <=  IAO & TAB  |  DAO & TBB  |  IEO & TCB  |  WAO & TDB  |  TMB  ; 
 ATG <=  IBG & TAC  |  DBG & TBC  |  EAG & TCC  |  WBG & TDC  |  TMC  ; 
 ABG <=  IBG & TAC  |  DBG & TBC  |  EAG & TCC  |  WBG & TDC  |  TMC  ; 
 DAG <= ICG ; 
 DAO <= ICO ; 
 DBG <= IDG ; 
 DBO <= IDO ; 
 qsi <= iqi ; 
 qqx <= qqd ; 
 QTO <= QTM ; 
 QTN <= QTM ; 
 ATO <=  IBO & TAD  |  DBO & TBD  |  ECO & TCD  |  WBO & TDD  |  TMD  ; 
 ABO <=  IBO & TAD  |  DBO & TBD  |  ECO & TCD  |  WBO & TDD  |  TMD  ; 
 OBG <=  DBG & TEB  |  EDG & TED  |  WDI & TEF  ; 
 OBO <=  DBO & TEB  |  EDO & TED  ; 
 EDG <= EAG ; 
 EDO <= ECO ; 
 eag <= ieg ; 
 eco <= ieo ; 
 QAA <= IJB & IJA ; 
 QAB <= IJB & IJA ; 
 QAC <= IJB & IJA ; 
 QAD <= IJB & IJA ; 
 QEA <=  QYB  |  QYC  ; 
 QEB <=  QNQ  |  QNU  ; 
 ocg <= pcg ; 
 oco <= pco ; 
 odg <= pdg ; 
 odo <= pdo ; 
 QSA <=  QSA & jxa & qtp  |  IQG  ; 
 OES <=  JJK & QML  |  JKE  |  QQE  ; 
 old <=  ZZO & QML  |  qab  |  gch  ; 
 OFC <= QRD ; 
 OQB <= JXA ; 
 OLB <= QKK ; 
 otf <= qsd ; 
 GDJ <= QCI & GDG ; 
 GDK <= QCI & GDH ; 
 GDL <= QCI & GDI ; 
 QCJ <= QCI & QCI ; 
 QSB <=  QSB & jxa & qtp  |  IQH  ; 
 OET <=  JKC  |  QMJ  |  QNA  |  RQB  ; 
 OEH <= QRF ; 
 oeq <= qqf ; 
 oer <= rsa ; 
 QTJ <= QTI ; 
 KAF <=  KAF & tlc  |  ZZI & QMG  ; 
 QTX <=  QTX & rji  |  QTJ & JTB  |  ZZI & QTN  ; 
 QTP <=  ZZO & rji  |  ZZO & JTB  |  qtm & QTN  ; 
 OFA <= QNB & RLB ; 
 ofb <=  rlb  |  qsh  |  QSB  ; 
 oqa <=  rla  |  qsh  |  QSB  ; 
 PAH <=  PAH & jgh & tpa  |  pah & JGH  |  AAH & TPA  ; 
 PCH <=  PAH & jgh & tpa  |  pah & JGH  |  AAH & TPA  ; 
 PEH <=  PAH & jgh & tpa  |  pah & JGH  |  AAH & TPA  ; 
 BAH <=  BAH & jdh & tfa  |  bah & JDH  |  AAH & TFA  ; 
 BEH <=  BAH & jdh & tfa  |  bah & JDH  |  AAH & TFA  ; 
 PAP <=  PAP & jgp & tpb  |  pap & JGP  |  AAP & TPB  ; 
 PCP <=  PAP & jgp & tpb  |  pap & JGP  |  AAP & TPB  ; 
 PEP <=  PAP & jgp & tpb  |  pap & JGP  |  AAP & TPB  ; 
 qvf <=  quf  |  jfa  |  jfb  |  jfc  |  jfd  ; 
 qvg <=  quf  |  jfa  |  jfb  |  jfc  |  jfd  ; 
 BAP <=  BAP & jdp & tfb  |  bap & JDP  |  AAP & TFB  ; 
 BEP <=  BAP & jdp & tfb  |  bap & JDP  |  AAP & TFB  ; 
 OLA <= QKE & qkd ; 
 PBH <=  PBH & jhh & tpc  |  pbh & JHH  |  ABH & TPC  ; 
 PDH <=  PBH & jhh & tpc  |  pbh & JHH  |  ABH & TPC  ; 
 PFH <=  PBH & jhh & tpc  |  pbh & JHH  |  ABH & TPC  ; 
 BBH <=  BBH & jeh & tfc  |  bbh & JEH  |  ABH & TFC  ; 
 BFH <=  BBH & jeh & tfc  |  bbh & JEH  |  ABH & TFC  ; 
 PBP <=  PBP & jhp & tpd  |  pbp & JHP  |  ABP & TPD  ; 
 PDP <=  PBP & jhp & tpd  |  pbp & JHP  |  ABP & TPD  ; 
 BBP <=  BBP & jep & tfd  |  bbp & JEP  |  ABP & TFD  ; 
 HNA <= HMA ; 
 HNB <= HMB ; 
 HNC <= HMC ; 
 QSC <=  QSC & jxb  |  ZZO & qln  |  RRF  ; 
 QSD <=  ZZO & jxb  |  QSD & qln  |  RRH  ; 
 HPA <= HOA ; 
 HPB <= HOB ; 
 HPC <= HOC ; 
 QSF <= QSE ; 
 RSB <= RSA ; 
 QSG <= QSF ; 
 QQK <=  JJE & RLC & JLG  ; 
 QQR <=  JJE & RLC & JLG  ; 
 HOA <= HNA ; 
 HOB <= HNB ; 
 HOC <= HNC ; 
 RRE <= RRD ; 
 RRF <= RRE ; 
 rrg <= jxb ; 
 RRH <= RRG ; 
 RRB <= RRA ; 
 RSC <= RSB ; 
 RRC <= RRB ; 
 RRD <= RRC ; 
 AQH <= AOH ; 
 AQI <= AOI ; 
 AQJ <= AOJ ; 
 AQK <= AOK ; 
 ach <= wch & QKR |  aqh & qkr ; 
 acp <= wcp & QKR |  aqp & qkr ; 
 adh <= wdh & QKR |  arh & qkr ; 
 AQL <= AOL ; 
 AQM <= AOM ; 
 AQN <= AON ; 
 AQO <= AOO ; 
 CJA <=  BND  |  ZZI & BNB  |  BNA  |  ZZO & ZZI  |  BNC  ; 
 AQP <= AOP ; 
 ARA <= APA ; 
 ARB <= APB ; 
 ARC <= APC ; 
 CJB <=  BNH  |  BNE  |  BNF  |  ZZO & ZZI  |  BNG  ; 
 ARD <= APD ; 
 ARE <= APE ; 
 ARF <= APF ; 
 ARG <= APG ; 
 ARH <= APH ; 
 ARI <= API ; 
 ARJ <= APJ ; 
 ARK <= APK ; 
 ARL <= APL ; 
 ARM <= APM ; 
 ARN <= APN ; 
 ARO <= APO ; 
 QQJ <=  JQJ & qtq  |  JCP & qcx  |  JQH & qcx  ; 
 QQH <=  JQI & qtq  |  JCP & qcx  |  JQH & qcx  ; 
 RBF <= qqj & RBE ; 
 RBG <= qqj & RBF ; 
 RBH <= qqj & RBG ; 
 RBI <= qqj & RBH ; 
 QSH <= QSD & QSF ; 
 QSE <= QSD & QSD ; 
 QQN <=  ZZI & QQL  ; 
 QQM <=  JCV & QQL  ; 
 QQL <=  QCX & qqj & JOL  |  QKY  ; 
 QQS <=  QCX & qqj & JOL  |  QKY  ; 
 rqa <=  jqb  |  jcq  ; 
 ASH <=  IAH & TAA  |  DAH & TBA  |  IEH & TCA  |  WAH & TDA  |  TMA  ; 
 AAH <=  IAH & TAA  |  DAH & TBA  |  IEH & TCA  |  WAH & TDA  |  TMA  ; 
 OAH <=  DAH & TEA  |  EAH & TEC  |  WCJ & TEE  ; 
 OAP <=  DAP & TEA  |  EAP & TEC  |  WDB & TEE  ; 
 ASP <=  IAP & TAB  |  DAP & TBB  |  IEP & TCB  |  WAP & TDB  |  TMB  ; 
 AAP <=  IAP & TAB  |  DAP & TBB  |  IEP & TCB  |  WAP & TDB  |  TMB  ; 
 ATH <=  IBH & TAC  |  DBH & TBC  |  EAH & TCC  |  WBH & TDC  |  TMC  ; 
 ABH <=  IBH & TAC  |  DBH & TBC  |  EAH & TCC  |  WBH & TDC  |  TMC  ; 
 DAH <= ICH ; 
 DAP <= ICP ; 
 DBH <= IDH ; 
 DBP <= IDP ; 
 ABP <=  IBP & TAD  |  DBP & TBD  |  EAP & TCD  |  WBP & TDD  |  TMD  ; 
 ATP <=  IBP & TAD  |  DBP & TBD  |  EAP & TCD  |  WBP & TDD  |  TMD  ; 
 OBH <=  DBH & TEB  |  EDH & TED  |  WDJ & TEF  ; 
 OBP <=  DBP & TEB  |  EDP & TED  ; 
 eah <= ieh ; 
 eap <= iep ; 
 ebp <= iep ; 
 OGJ <=  JOE & JOP  |  JOF & JOP  |  JOG & JOP  |  JOH & JOP  ; 
 EDH <= EAH ; 
 EDP <= EAP ; 
 QKT <= JCY ; 
 och <= pch ; 
 ocp <= pcp ; 
 odh <= pdh ; 
 odp <= pdp ; 
 OGE <=  HMA & JOE  |  HNA & JOF  |  HOA & JOG  |  HPA & JOH  ; 
 OGF <=  HMB & JOE  |  HNB & JOF  |  HOB & JOG  |  HPB & JOH  ; 
 OEG <=  RLD & qqg  |  RLD & QQJ  |  JCY & JIE  ; 
 QFC <=  RLD & qqg  |  RLD & QQJ  |  JCY & JIE  ; 
 OGG <=  HMC & JOE  |  HNC & JOF  |  HOC & JOG  |  HPC & JOH  ; 
 OGH <=  JOE & JOK  |  JOF & JOK  |  JOG & JOK  |  JOH & JOK  ; 
 QCH <=  JOE & JOK  |  JOF & JOK  |  JOG & JOK  |  JOH & JOK  ; 
 OEV <=  QNQ  |  QNU  |  QQD  ; 
 OEL <=  RKA  |  QLJ  |  JKD  ; 
 OEN <= JKC ; 
 OEO <= JKC ; 
 OEX <= QYB ; 
 OEY <= QYC ; 
 RRA <= IQG ; 
 RSA <= RRH ; 
 qlx <= qlp ; 
 OEK <=  JJK & QSG  ; 
 OEU <=  QMI  |  QNI  ; 
 OEW <=  QMK  |  QMJ  ; 
end
endmodule;
