module ga( IZZ,
 IAA, 
 IAB, 
 IAC, 
 IAD, 
 IAE, 
 IAF, 
 IAG, 
 IAH, 
 IAI, 
 IAJ, 
 IAK, 
 IAL, 
 IAM, 
 IAN, 
 IAO, 
 IAP, 
 IBA, 
 IBB, 
 IBC, 
 IBD, 
 IBE, 
 IBF, 
 IBG, 
 IBH, 
 IBI, 
 IBJ, 
 IBK, 
 IBL, 
 IBM, 
 IBN, 
 IBO, 
 IBP, 
 ICA, 
 ICB, 
 ICC, 
 ICD, 
 ICE, 
 ICF, 
 ICG, 
 ICH, 
 ICI, 
 ICJ, 
 ICK, 
 ICL, 
 ICM, 
 ICN, 
 ICO, 
 ICP, 
 IDA, 
 IDB, 
 IDC, 
 IDD, 
 IDE, 
 IDF, 
 IDG, 
 IDH, 
 IDI, 
 IDJ, 
 IDK, 
 IDL, 
 IDM, 
 IDN, 
 IDO, 
 IDP, 
 IGA, 
 IPB, 
 IPC, 
 IPD, 
 OAA, 
 OAB, 
 OAC, 
 OAD, 
 OAE, 
 OAF, 
 OAG, 
 OAH, 
 OAI, 
 OAJ, 
 OAK, 
 OAL, 
 OAM, 
 OAN, 
 OAO, 
 OAP, 
 OBA, 
 OBB, 
 OBC, 
 OBD, 
 OBE, 
 OBF, 
 OBG, 
 OBH, 
 OBI, 
 OBJ, 
 OBK, 
 OBL, 
 OBM, 
 OBN, 
 OBO, 
 OBP, 
 OCA, 
 OCB, 
 OCC, 
 OCD, 
 OCE, 
 OCF, 
 OCG, 
 OCH, 
 OCI, 
 OCJ, 
 OCK, 
 OCL, 
 OCM, 
 OCN, 
 OCO, 
 OCP, 
 ODA, 
 ODB, 
 ODC, 
 ODD, 
 ODE, 
 ODF, 
 ODG, 
 ODH, 
 ODI, 
 ODJ, 
 ODK, 
 ODL, 
 ODM, 
 ODN, 
 ODO, 
ODP ); 
    
 input IZZ; 
 input IAA; 
 input IAB; 
 input IAC; 
 input IAD; 
 input IAE; 
 input IAF; 
 input IAG; 
 input IAH; 
 input IAI; 
 input IAJ; 
 input IAK; 
 input IAL; 
 input IAM; 
 input IAN; 
 input IAO; 
 input IAP; 
 input IBA; 
 input IBB; 
 input IBC; 
 input IBD; 
 input IBE; 
 input IBF; 
 input IBG; 
 input IBH; 
 input IBI; 
 input IBJ; 
 input IBK; 
 input IBL; 
 input IBM; 
 input IBN; 
 input IBO; 
 input IBP; 
 input ICA; 
 input ICB; 
 input ICC; 
 input ICD; 
 input ICE; 
 input ICF; 
 input ICG; 
 input ICH; 
 input ICI; 
 input ICJ; 
 input ICK; 
 input ICL; 
 input ICM; 
 input ICN; 
 input ICO; 
 input ICP; 
 input IDA; 
 input IDB; 
 input IDC; 
 input IDD; 
 input IDE; 
 input IDF; 
 input IDG; 
 input IDH; 
 input IDI; 
 input IDJ; 
 input IDK; 
 input IDL; 
 input IDM; 
 input IDN; 
 input IDO; 
 input IDP; 
 input IGA; 
 input IPB; 
 input IPC; 
 input IPD; 
 output OAA; 
 output OAB; 
 output OAC; 
 output OAD; 
 output OAE; 
 output OAF; 
 output OAG; 
 output OAH; 
 output OAI; 
 output OAJ; 
 output OAK; 
 output OAL; 
 output OAM; 
 output OAN; 
 output OAO; 
 output OAP; 
 output OBA; 
 output OBB; 
 output OBC; 
 output OBD; 
 output OBE; 
 output OBF; 
 output OBG; 
 output OBH; 
 output OBI; 
 output OBJ; 
 output OBK; 
 output OBL; 
 output OBM; 
 output OBN; 
 output OBO; 
 output OBP; 
 output OCA; 
 output OCB; 
 output OCC; 
 output OCD; 
 output OCE; 
 output OCF; 
 output OCG; 
 output OCH; 
 output OCI; 
 output OCJ; 
 output OCK; 
 output OCL; 
 output OCM; 
 output OCN; 
 output OCO; 
 output OCP; 
 output ODA; 
 output ODB; 
 output ODC; 
 output ODD; 
 output ODE; 
 output ODF; 
 output ODG; 
 output ODH; 
 output ODI; 
 output ODJ; 
 output ODK; 
 output ODL; 
 output ODM; 
 output ODN; 
 output ODO; 
 output ODP; 
  
  
reg  aaa ;
reg  aab ;
reg  aac ;
reg  aad ;
reg  aba ;
reg  abb ;
reg  abc ;
reg  abd ;
reg  aca ;
reg  acb ;
reg  acc ;
reg  acd ;
reg  ada ;
reg  adb ;
reg  adc ;
reg  add ;
reg  aea ;
reg  aeb ;
reg  aec ;
reg  aed ;
reg  afa ;
reg  afb ;
reg  afc ;
reg  afd ;
reg  aga ;
reg  agb ;
reg  agc ;
reg  agd ;
reg  aha ;
reg  ahb ;
reg  ahc ;
reg  ahd ;
reg  aia ;
reg  aib ;
reg  aic ;
reg  aid ;
reg  aja ;
reg  ajb ;
reg  ajc ;
reg  ajd ;
reg  aka ;
reg  akb ;
reg  akc ;
reg  akd ;
reg  ala ;
reg  alb ;
reg  alc ;
reg  ald ;
reg  ama ;
reg  amb ;
reg  amc ;
reg  amd ;
reg  ana ;
reg  anb ;
reg  anc ;
reg  andd  ;
reg  aoa ;
reg  aob ;
reg  aoc ;
reg  aod ;
reg  apa ;
reg  apb ;
reg  apc ;
reg  apd ;
reg  BAA ;
reg  BAB ;
reg  BAC ;
reg  BAD ;
reg  BBA ;
reg  BBB ;
reg  BBC ;
reg  BBD ;
reg  BBF ;
reg  BBG ;
reg  BCA ;
reg  BCB ;
reg  BCC ;
reg  BCD ;
reg  BCF ;
reg  BCG ;
reg  BDA ;
reg  BDB ;
reg  BDC ;
reg  BDD ;
reg  BDF ;
reg  BDG ;
reg  BEA ;
reg  BEB ;
reg  BEC ;
reg  BED ;
reg  BEF ;
reg  BEG ;
reg  BFA ;
reg  BFB ;
reg  BFC ;
reg  BFD ;
reg  BFF ;
reg  BFG ;
reg  BGA ;
reg  BGB ;
reg  BGC ;
reg  BGD ;
reg  BGF ;
reg  BGG ;
reg  BHA ;
reg  BHB ;
reg  BHC ;
reg  BHD ;
reg  BHF ;
reg  BHG ;
reg  BIA ;
reg  BIB ;
reg  BIC ;
reg  BID ;
reg  BIF ;
reg  BIG ;
reg  BJA ;
reg  BJB ;
reg  BJC ;
reg  BJD ;
reg  BJF ;
reg  BJG ;
reg  BKA ;
reg  BKB ;
reg  BKC ;
reg  BKD ;
reg  BKF ;
reg  BKG ;
reg  BLA ;
reg  BLB ;
reg  BLC ;
reg  BLD ;
reg  BLF ;
reg  BLG ;
reg  BMA ;
reg  BMB ;
reg  BMC ;
reg  BMD ;
reg  BMF ;
reg  BMG ;
reg  BNA ;
reg  BNB ;
reg  BNC ;
reg  BND ;
reg  BNF ;
reg  BNG ;
reg  BOA ;
reg  BOB ;
reg  BOC ;
reg  BOD ;
reg  BOF ;
reg  BOG ;
reg  BPA ;
reg  BPB ;
reg  BPC ;
reg  BPD ;
reg  gaa ;
reg  gab ;
reg  gac ;
reg  gad ;
reg  gba ;
reg  gbb ;
reg  gbc ;
reg  gbd ;
reg  gca ;
reg  gcb ;
reg  gcc ;
reg  gcd ;
reg  gda ;
reg  gdb ;
reg  gdc ;
reg  gdd ;
reg  gea ;
reg  geb ;
reg  gec ;
reg  ged ;
reg  gfa ;
reg  gfb ;
reg  gfc ;
reg  gfd ;
reg  gga ;
reg  ggb ;
reg  ggc ;
reg  ggd ;
reg  gha ;
reg  ghb ;
reg  ghc ;
reg  ghd ;
reg  gia ;
reg  gib ;
reg  gic ;
reg  gid ;
reg  gja ;
reg  gjb ;
reg  gjc ;
reg  gjd ;
reg  gka ;
reg  gkb ;
reg  gkc ;
reg  gkd ;
reg  gla ;
reg  glb ;
reg  glc ;
reg  gld ;
reg  gma ;
reg  gmb ;
reg  gmc ;
reg  gmd ;
reg  gna ;
reg  gnb ;
reg  gnc ;
reg  gnd ;
reg  goa ;
reg  gob ;
reg  goc ;
reg  god ;
reg  gpa ;
reg  gpb ;
reg  gpc ;
reg  gpd ;
reg  hba ;
reg  hbb ;
reg  hbc ;
reg  hbd ;
reg  hca ;
reg  hcb ;
reg  hcc ;
reg  hcd ;
reg  hda ;
reg  hdb ;
reg  hdc ;
reg  hdd ;
reg  hea ;
reg  heb ;
reg  hec ;
reg  hed ;
reg  hfa ;
reg  hfb ;
reg  hfc ;
reg  hfd ;
reg  hga ;
reg  hgb ;
reg  hgc ;
reg  hgd ;
reg  hha ;
reg  hhb ;
reg  hhc ;
reg  hhd ;
reg  hia ;
reg  hib ;
reg  hic ;
reg  hid ;
reg  hja ;
reg  hjb ;
reg  hjc ;
reg  hjd ;
reg  hka ;
reg  hkb ;
reg  hkc ;
reg  hkd ;
reg  hla ;
reg  hlb ;
reg  hlc ;
reg  hld ;
reg  hma ;
reg  hmb ;
reg  hmc ;
reg  hmd ;
reg  hna ;
reg  hnb ;
reg  hnc ;
reg  hnd ;
reg  hoa ;
reg  hob ;
reg  hoc ;
reg  hod ;
reg  hpa ;
reg  hpb ;
reg  hpc ;
reg  hpd ;
reg  KAB ;
reg  KAC ;
reg  KAD ;
reg  KBC ;
reg  KBD ;
reg  KCD ;
reg  lbc ;
reg  lbd ;
reg  lcd ;
reg  maa ;
reg  mab ;
reg  mac ;
reg  mba ;
reg  mbb ;
reg  mbc ;
reg  mca ;
reg  mcb ;
reg  mcc ;
reg  mda ;
reg  mdb ;
reg  mdc ;
reg  nba ;
reg  nbb ;
reg  nbc ;
reg  nca ;
reg  ncb ;
reg  ncc ;
reg  nda ;
reg  ndb ;
reg  ndc ;
reg  OAA ;
reg  OAB ;
reg  OAC ;
reg  OAD ;
reg  OAE ;
reg  OAF ;
reg  OAG ;
reg  OAH ;
reg  OAI ;
reg  OAJ ;
reg  OAK ;
reg  OAL ;
reg  OAM ;
reg  OAN ;
reg  OAO ;
reg  OAP ;
reg  OBA ;
reg  OBB ;
reg  OBC ;
reg  OBD ;
reg  OBE ;
reg  OBF ;
reg  OBG ;
reg  OBH ;
reg  OBI ;
reg  OBJ ;
reg  OBK ;
reg  OBL ;
reg  OBM ;
reg  OBN ;
reg  OBO ;
reg  OBP ;
reg  OCA ;
reg  OCB ;
reg  OCC ;
reg  OCD ;
reg  OCE ;
reg  OCF ;
reg  OCG ;
reg  OCH ;
reg  OCI ;
reg  OCJ ;
reg  OCK ;
reg  OCL ;
reg  OCM ;
reg  OCN ;
reg  OCO ;
reg  OCP ;
reg  ODA ;
reg  ODB ;
reg  ODC ;
reg  ODD ;
reg  ODE ;
reg  ODF ;
reg  ODG ;
reg  ODH ;
reg  ODI ;
reg  ODJ ;
reg  ODK ;
reg  ODL ;
reg  ODM ;
reg  ODN ;
reg  ODO ;
reg  ODP ;
reg  qaa ;
reg  QAB ;
reg  QAC ;
reg  QAD ;
reg  qba ;
reg  qbb ;
reg  qbc ;
reg  qbd ;
reg  qbe ;
reg  QCA ;
reg  qcb ;
reg  qcc ;
reg  qcd ;
reg  qce ;
reg  QDA ;
reg  QDB ;
reg  QDC ;
reg  QDD ;
reg  QDE ;
reg  qdf ;
reg  QEA ;
reg  QEC ;
reg  QED ;
reg  QEE ;
reg  QEF ;
reg  qeg ;
reg  QFC ;
reg  QFE ;
reg  RAA ;
reg  RAB ;
reg  RAC ;
reg  RAD ;
reg  RAE ;
reg  raf ;
reg  RBA ;
reg  RBB ;
reg  RBC ;
reg  RBD ;
reg  RBE ;
reg  rbf ;
reg  RCA ;
reg  RCB ;
reg  RCC ;
reg  RCD ;
reg  RCE ;
reg  rcf ;
reg  RDA ;
reg  RDB ;
reg  RDC ;
reg  RDD ;
reg  RDE ;
reg  rdf ;
reg  rea ;
reg  reb ;
reg  rec ;
reg  red ;
reg  ree ;
reg  rfa ;
reg  rfb ;
reg  rfc ;
reg  rfd ;
reg  rfe ;
reg  rga ;
reg  rgb ;
reg  rgc ;
reg  rgd ;
reg  rge ;
reg  rha ;
reg  rhb ;
reg  rhc ;
reg  rhd ;
reg  rhe ;
reg  RMA ;
reg  RMB ;
reg  RMC ;
reg  RMD ;
reg  rme ;
reg  rmf ;
reg  RMG ;
reg  SAA ;
reg  SAB ;
reg  SAC ;
reg  sba ;
reg  sbb ;
reg  sbc ;
reg  SBD ;
reg  SBE ;
reg  SBF ;
reg  SBG ;
reg  SBH ;
reg  SBI ;
reg  SBJ ;
reg  SBK ;
reg  sca ;
reg  scb ;
reg  scc ;
reg  scd ;
reg  sce ;
reg  scf ;
reg  SCG ;
reg  SCH ;
reg  sda ;
reg  swa ;
reg  swb ;
reg  swc ;
reg  swd ;
reg  swe ;
reg  swf ;
reg  swg ;
reg  swh ;
reg  swi ;
reg  swj ;
reg  swk ;
reg  swl ;
reg  swm ;
reg  swn ;
reg  swo ;
reg  swp ;
reg  sxa ;
reg  sxb ;
reg  sxc ;
reg  sxd ;
reg  sxe ;
reg  sxf ;
reg  sxg ;
reg  sxh ;
reg  sxi ;
reg  sxj ;
reg  sxk ;
reg  sxl ;
reg  sxm ;
reg  sxn ;
reg  sxo ;
reg  sxp ;
reg  sya ;
reg  syb ;
reg  syc ;
reg  syd ;
reg  sye ;
reg  syf ;
reg  syg ;
reg  syh ;
reg  syi ;
reg  syj ;
reg  syk ;
reg  syl ;
reg  sym ;
reg  syn ;
reg  syo ;
reg  syp ;
reg  sza ;
reg  szb ;
reg  szc ;
reg  szd ;
reg  sze ;
reg  szf ;
reg  szg ;
reg  szh ;
reg  szi ;
reg  szj ;
reg  szk ;
reg  szl ;
reg  szm ;
reg  szn ;
reg  szo ;
reg  szp ;
reg  TAA ;
reg  TAB ;
reg  TAC ;
reg  TAD ;
reg  TAE ;
reg  TAF ;
reg  TAG ;
reg  TAH ;
reg  tba ;
reg  tbb ;
reg  tbc ;
reg  tbd ;
reg  tbe ;
reg  tbf ;
reg  tbg ;
reg  tbh ;
reg  TCA ;
reg  TCB ;
reg  TCC ;
reg  TCD ;
reg  TCE ;
reg  TCF ;
reg  TCG ;
reg  TCH ;
reg  TCI ;
reg  TCJ ;
reg  TCK ;
reg  TCL ;
reg  TCM ;
reg  TCN ;
reg  TCO ;
reg  TCP ;
reg  TDA ;
reg  TDB ;
reg  TDC ;
reg  TDD ;
reg  TDE ;
reg  TDF ;
reg  TDG ;
reg  TDH ;
reg  TEA ;
reg  TEB ;
reg  TEC ;
reg  TFA ;
reg  TFB ;
reg  VAA ;
reg  VBA ;
reg  VBB ;
reg  vca ;
reg  vcb ;
reg  VCC ;
reg  VCD ;
reg  vda ;
reg  vdb ;
reg  VDC ;
reg  vea ;
reg  VEB ;
reg  vma ;
reg  vmb ;
reg  vmc ;
reg  vmd ;
reg  vna ;
reg  vnb ;
reg  vnc ;
reg  vnd ;
reg  voa ;
reg  vob ;
reg  voc ;
reg  vod ;
reg  vpa ;
reg  vpb ;
reg  vpc ;
reg  vpd ;
reg  vqa ;
reg  vqb ;
reg  vqc ;
reg  vqd ;
reg  vra ;
reg  vrb ;
reg  vrc ;
reg  vrd ;
reg  vsa ;
reg  vsb ;
reg  vsc ;
reg  vsd ;
reg  vta ;
reg  vtb ;
reg  vtc ;
reg  vtd ;
reg  vua ;
reg  vub ;
reg  vuc ;
reg  vud ;
reg  vva ;
reg  vvb ;
reg  vvc ;
reg  vvd ;
reg  vwa ;
reg  vwb ;
reg  vwc ;
reg  vwd ;
reg  vxa ;
reg  vxb ;
reg  vxc ;
reg  vxd ;
reg  XAB ;
reg  XAC ;
reg  XAD ;
reg  XAE ;
reg  xba ;
reg  xbb ;
reg  xbc ;
reg  xbd ;
reg  xbe ;
reg  xbf ;
reg  XMA ;
reg  XMB ;
reg  xmc ;
reg  xmd ;
reg  xme ;
reg  XPA ;
reg  XPB ;
reg  xpc ;
reg  xpd ;
reg  xpe ;
reg  XSA ;
reg  XSB ;
reg  xsc ;
reg  xsd ;
reg  xse ;
reg  xsf ;
reg  XVA ;
reg  XVB ;
reg  xvc ;
reg  xvd ;
reg  xve ;
reg  xvf ;
wire  AAA ;
wire  AAB ;
wire  AAC ;
wire  AAD ;
wire  ABA ;
wire  ABB ;
wire  ABC ;
wire  ABD ;
wire  ACA ;
wire  ACB ;
wire  ACC ;
wire  ACD ;
wire  ADA ;
wire  ADB ;
wire  ADC ;
wire  ADD ;
wire  AEA ;
wire  AEB ;
wire  AEC ;
wire  AED ;
wire  AFA ;
wire  AFB ;
wire  AFC ;
wire  AFD ;
wire  AGA ;
wire  AGB ;
wire  AGC ;
wire  AGD ;
wire  AHA ;
wire  AHB ;
wire  AHC ;
wire  AHD ;
wire  AIA ;
wire  AIB ;
wire  AIC ;
wire  AID ;
wire  AJA ;
wire  AJB ;
wire  AJC ;
wire  AJD ;
wire  AKA ;
wire  AKB ;
wire  AKC ;
wire  AKD ;
wire  ALA ;
wire  ALB ;
wire  ALC ;
wire  ALD ;
wire  AMA ;
wire  AMB ;
wire  AMC ;
wire  AMD ;
wire  ANA ;
wire  ANB ;
wire  ANC ;
wire  ANDD  ;
wire  AOA ;
wire  AOB ;
wire  AOC ;
wire  AOD ;
wire  APA ;
wire  APB ;
wire  APC ;
wire  APD ;
wire  baa ;
wire  bab ;
wire  bac ;
wire  bad ;
wire  bba ;
wire  bbb ;
wire  bbc ;
wire  bbd ;
wire  bbf ;
wire  bbg ;
wire  bca ;
wire  bcb ;
wire  bcc ;
wire  bcd ;
wire  bcf ;
wire  bcg ;
wire  bda ;
wire  bdb ;
wire  bdc ;
wire  bdd ;
wire  bdf ;
wire  bdg ;
wire  bea ;
wire  beb ;
wire  bec ;
wire  bed ;
wire  bef ;
wire  beg ;
wire  bfa ;
wire  bfb ;
wire  bfc ;
wire  bfd ;
wire  bff ;
wire  bfg ;
wire  bga ;
wire  bgb ;
wire  bgc ;
wire  bgd ;
wire  bgf ;
wire  bgg ;
wire  bha ;
wire  bhb ;
wire  bhc ;
wire  bhd ;
wire  bhf ;
wire  bhg ;
wire  bia ;
wire  bib ;
wire  bic ;
wire  bid ;
wire  bif ;
wire  big ;
wire  bja ;
wire  bjb ;
wire  bjc ;
wire  bjd ;
wire  bjf ;
wire  bjg ;
wire  bka ;
wire  bkb ;
wire  bkc ;
wire  bkd ;
wire  bkf ;
wire  bkg ;
wire  bla ;
wire  blb ;
wire  blc ;
wire  bld ;
wire  blf ;
wire  blg ;
wire  bma ;
wire  bmb ;
wire  bmc ;
wire  bmd ;
wire  bmf ;
wire  bmg ;
wire  bna ;
wire  bnb ;
wire  bnc ;
wire  bnd ;
wire  bnf ;
wire  bng ;
wire  boa ;
wire  bob ;
wire  boc ;
wire  bod ;
wire  bof ;
wire  bog ;
wire  bpa ;
wire  bpb ;
wire  bpc ;
wire  bpd ;
wire  cab ;
wire  CAB ;
wire  cac ;
wire  CAC ;
wire  cad ;
wire  CAD ;
wire  cae ;
wire  CAE ;
wire  cbb ;
wire  CBB ;
wire  cbc ;
wire  CBC ;
wire  cbd ;
wire  CBD ;
wire  cbe ;
wire  CBE ;
wire  ccb ;
wire  CCB ;
wire  ccc ;
wire  CCC ;
wire  ccd ;
wire  CCD ;
wire  cce ;
wire  CCE ;
wire  cdb ;
wire  CDB ;
wire  cdc ;
wire  CDC ;
wire  cdd ;
wire  CDD ;
wire  cde ;
wire  CDE ;
wire  ceb ;
wire  CEB ;
wire  cec ;
wire  CEC ;
wire  ced ;
wire  CED ;
wire  cee ;
wire  CEE ;
wire  cfb ;
wire  CFB ;
wire  cfc ;
wire  CFC ;
wire  cfd ;
wire  CFD ;
wire  cfe ;
wire  CFE ;
wire  cgb ;
wire  CGB ;
wire  cgc ;
wire  CGC ;
wire  cgd ;
wire  CGD ;
wire  cge ;
wire  CGE ;
wire  chb ;
wire  CHB ;
wire  chc ;
wire  CHC ;
wire  chd ;
wire  CHD ;
wire  che ;
wire  CHE ;
wire  cib ;
wire  CIB ;
wire  cic ;
wire  CIC ;
wire  cid ;
wire  CID ;
wire  cie ;
wire  CIE ;
wire  cjb ;
wire  CJB ;
wire  cjc ;
wire  CJC ;
wire  cjd ;
wire  CJD ;
wire  cje ;
wire  CJE ;
wire  ckb ;
wire  CKB ;
wire  ckc ;
wire  CKC ;
wire  ckd ;
wire  CKD ;
wire  cke ;
wire  CKE ;
wire  clb ;
wire  CLB ;
wire  clc ;
wire  CLC ;
wire  cld ;
wire  CLD ;
wire  cle ;
wire  CLE ;
wire  cmb ;
wire  CMB ;
wire  cmc ;
wire  CMC ;
wire  cmd ;
wire  CMD ;
wire  cme ;
wire  CME ;
wire  cnb ;
wire  CNB ;
wire  cnc ;
wire  CNC ;
wire  cnd ;
wire  CND ;
wire  cne ;
wire  CNE ;
wire  cob ;
wire  COB ;
wire  coc ;
wire  COC ;
wire  cod ;
wire  COD ;
wire  coe ;
wire  COE ;
wire  cpb ;
wire  CPB ;
wire  cpc ;
wire  CPC ;
wire  cpd ;
wire  CPD ;
wire  dbb ;
wire  DBB ;
wire  dbc ;
wire  DBC ;
wire  dbd ;
wire  DBD ;
wire  dcb ;
wire  DCB ;
wire  dcc ;
wire  DCC ;
wire  dcd ;
wire  DCD ;
wire  ddb ;
wire  DDB ;
wire  ddc ;
wire  DDC ;
wire  ddd ;
wire  DDD ;
wire  deb ;
wire  DEB ;
wire  dec ;
wire  DEC ;
wire  ded ;
wire  DED ;
wire  dfb ;
wire  DFB ;
wire  dfc ;
wire  DFC ;
wire  dfd ;
wire  DFD ;
wire  dgb ;
wire  DGB ;
wire  dgc ;
wire  DGC ;
wire  dgd ;
wire  DGD ;
wire  dhb ;
wire  DHB ;
wire  dhc ;
wire  DHC ;
wire  dhd ;
wire  DHD ;
wire  dib ;
wire  DIB ;
wire  dic ;
wire  DIC ;
wire  did ;
wire  DID ;
wire  djb ;
wire  DJB ;
wire  djc ;
wire  DJC ;
wire  djd ;
wire  DJD ;
wire  dkb ;
wire  DKB ;
wire  dkc ;
wire  DKC ;
wire  dkd ;
wire  DKD ;
wire  dlb ;
wire  DLB ;
wire  dlc ;
wire  DLC ;
wire  dld ;
wire  DLD ;
wire  dmb ;
wire  DMB ;
wire  dmc ;
wire  DMC ;
wire  dmd ;
wire  DMD ;
wire  dnb ;
wire  DNB ;
wire  dnc ;
wire  DNC ;
wire  dnd ;
wire  DND ;
wire  dob ;
wire  DOB ;
wire  doc ;
wire  DOC ;
wire  dod ;
wire  DOD ;
wire  dpb ;
wire  DPB ;
wire  dpc ;
wire  DPC ;
wire  dpd ;
wire  DPD ;
wire  eaa ;
wire  EAA ;
wire  eab ;
wire  EAB ;
wire  eac ;
wire  EAC ;
wire  ead ;
wire  EAD ;
wire  eba ;
wire  EBA ;
wire  ebb ;
wire  EBB ;
wire  ebc ;
wire  EBC ;
wire  ebd ;
wire  EBD ;
wire  eca ;
wire  ECA ;
wire  ecb ;
wire  ECB ;
wire  ecc ;
wire  ECC ;
wire  ecd ;
wire  ECD ;
wire  eda ;
wire  EDA ;
wire  edb ;
wire  EDB ;
wire  edc ;
wire  EDC ;
wire  edd ;
wire  EDD ;
wire  eea ;
wire  EEA ;
wire  eeb ;
wire  EEB ;
wire  eec ;
wire  EEC ;
wire  eed ;
wire  EED ;
wire  efa ;
wire  EFA ;
wire  efb ;
wire  EFB ;
wire  efc ;
wire  EFC ;
wire  efd ;
wire  EFD ;
wire  ega ;
wire  EGA ;
wire  egb ;
wire  EGB ;
wire  egc ;
wire  EGC ;
wire  egd ;
wire  EGD ;
wire  eha ;
wire  EHA ;
wire  ehb ;
wire  EHB ;
wire  ehc ;
wire  EHC ;
wire  ehd ;
wire  EHD ;
wire  eia ;
wire  EIA ;
wire  eib ;
wire  EIB ;
wire  eic ;
wire  EIC ;
wire  eid ;
wire  EID ;
wire  eja ;
wire  EJA ;
wire  ejb ;
wire  EJB ;
wire  ejc ;
wire  EJC ;
wire  ejd ;
wire  EJD ;
wire  eka ;
wire  EKA ;
wire  ekb ;
wire  EKB ;
wire  ekc ;
wire  EKC ;
wire  ekd ;
wire  EKD ;
wire  ela ;
wire  ELA ;
wire  elb ;
wire  ELB ;
wire  elc ;
wire  ELC ;
wire  eld ;
wire  ELD ;
wire  ema ;
wire  EMA ;
wire  emb ;
wire  EMB ;
wire  emc ;
wire  EMC ;
wire  emd ;
wire  EMD ;
wire  ena ;
wire  ENA ;
wire  enb ;
wire  ENB ;
wire  enc ;
wire  ENC ;
wire  endd ;
wire  ENDD ;
wire  eoa ;
wire  EOA ;
wire  eob ;
wire  EOB ;
wire  eoc ;
wire  EOC ;
wire  eod ;
wire  EOD ;
wire  epa ;
wire  EPA ;
wire  epb ;
wire  EPB ;
wire  epc ;
wire  EPC ;
wire  epd ;
wire  EPD ;
wire  fab ;
wire  FAB ;
wire  fac ;
wire  FAC ;
wire  fad ;
wire  FAD ;
wire  fae ;
wire  FAE ;
wire  faf ;
wire  FAF ;
wire  fag ;
wire  FAG ;
wire  fah ;
wire  FAH ;
wire  fai ;
wire  FAI ;
wire  faj ;
wire  FAJ ;
wire  fak ;
wire  FAK ;
wire  fal ;
wire  FAL ;
wire  fam ;
wire  FAM ;
wire  fan ;
wire  FAN ;
wire  fao ;
wire  FAO ;
wire  fbf ;
wire  FBF ;
wire  fbg ;
wire  FBG ;
wire  fbj ;
wire  FBJ ;
wire  fbk ;
wire  FBK ;
wire  fbn ;
wire  FBN ;
wire  fbo ;
wire  FBO ;
wire  GAA ;
wire  GAB ;
wire  GAC ;
wire  GAD ;
wire  GBA ;
wire  GBB ;
wire  GBC ;
wire  GBD ;
wire  GCA ;
wire  GCB ;
wire  GCC ;
wire  GCD ;
wire  GDA ;
wire  GDB ;
wire  GDC ;
wire  GDD ;
wire  GEA ;
wire  GEB ;
wire  GEC ;
wire  GED ;
wire  GFA ;
wire  GFB ;
wire  GFC ;
wire  GFD ;
wire  GGA ;
wire  GGB ;
wire  GGC ;
wire  GGD ;
wire  GHA ;
wire  GHB ;
wire  GHC ;
wire  GHD ;
wire  GIA ;
wire  GIB ;
wire  GIC ;
wire  GID ;
wire  GJA ;
wire  GJB ;
wire  GJC ;
wire  GJD ;
wire  GKA ;
wire  GKB ;
wire  GKC ;
wire  GKD ;
wire  GLA ;
wire  GLB ;
wire  GLC ;
wire  GLD ;
wire  GMA ;
wire  GMB ;
wire  GMC ;
wire  GMD ;
wire  GNA ;
wire  GNB ;
wire  GNC ;
wire  GND ;
wire  GOA ;
wire  GOB ;
wire  GOC ;
wire  GOD ;
wire  GPA ;
wire  GPB ;
wire  GPC ;
wire  GPD ;
wire  HBA ;
wire  HBB ;
wire  HBC ;
wire  HBD ;
wire  HCA ;
wire  HCB ;
wire  HCC ;
wire  HCD ;
wire  HDA ;
wire  HDB ;
wire  HDC ;
wire  HDD ;
wire  HEA ;
wire  HEB ;
wire  HEC ;
wire  HED ;
wire  HFA ;
wire  HFB ;
wire  HFC ;
wire  HFD ;
wire  HGA ;
wire  HGB ;
wire  HGC ;
wire  HGD ;
wire  HHA ;
wire  HHB ;
wire  HHC ;
wire  HHD ;
wire  HIA ;
wire  HIB ;
wire  HIC ;
wire  HID ;
wire  HJA ;
wire  HJB ;
wire  HJC ;
wire  HJD ;
wire  HKA ;
wire  HKB ;
wire  HKC ;
wire  HKD ;
wire  HLA ;
wire  HLB ;
wire  HLC ;
wire  HLD ;
wire  HMA ;
wire  HMB ;
wire  HMC ;
wire  HMD ;
wire  HNA ;
wire  HNB ;
wire  HNC ;
wire  HND ;
wire  HOA ;
wire  HOB ;
wire  HOC ;
wire  HOD ;
wire  HPA ;
wire  HPB ;
wire  HPC ;
wire  HPD ;
wire  iaa ;
wire  iab ;
wire  iac ;
wire  iad ;
wire  iae ;
wire  iaf ;
wire  iag ;
wire  iah ;
wire  iai ;
wire  iaj ;
wire  iak ;
wire  ial ;
wire  iam ;
wire  ian ;
wire  iao ;
wire  iap ;
wire  iba ;
wire  ibb ;
wire  ibc ;
wire  ibd ;
wire  ibe ;
wire  ibf ;
wire  ibg ;
wire  ibh ;
wire  ibi ;
wire  ibj ;
wire  ibk ;
wire  ibl ;
wire  ibm ;
wire  ibn ;
wire  ibo ;
wire  ibp ;
wire  ica ;
wire  icb ;
wire  icc ;
wire  icd ;
wire  ice ;
wire  icf ;
wire  icg ;
wire  ich ;
wire  ici ;
wire  icj ;
wire  ick ;
wire  icl ;
wire  icm ;
wire  icn ;
wire  ico ;
wire  icp ;
wire  ida ;
wire  idb ;
wire  idc ;
wire  idd ;
wire  ide ;
wire  idf ;
wire  idg ;
wire  idh ;
wire  idi ;
wire  idj ;
wire  idk ;
wire  idl ;
wire  idm ;
wire  idn ;
wire  ido ;
wire  idp ;
wire  iga ;
wire  ipb ;
wire  ipc ;
wire  ipd ;
wire  jaa ;
wire  JAA ;
wire  jab ;
wire  JAB ;
wire  jac ;
wire  JAC ;
wire  jad ;
wire  JAD ;
wire  jae ;
wire  JAE ;
wire  jaf ;
wire  JAF ;
wire  jag ;
wire  JAG ;
wire  jah ;
wire  JAH ;
wire  jba ;
wire  JBA ;
wire  jbb ;
wire  JBB ;
wire  jbc ;
wire  JBC ;
wire  jbd ;
wire  JBD ;
wire  jbe ;
wire  JBE ;
wire  jbf ;
wire  JBF ;
wire  jbg ;
wire  JBG ;
wire  jbh ;
wire  JBH ;
wire  jbi ;
wire  JBI ;
wire  jbj ;
wire  JBJ ;
wire  jbk ;
wire  JBK ;
wire  jbl ;
wire  JBL ;
wire  jca ;
wire  JCA ;
wire  jcb ;
wire  JCB ;
wire  jcc ;
wire  JCC ;
wire  jcd ;
wire  JCD ;
wire  kab ;
wire  kac ;
wire  kad ;
wire  kbc ;
wire  kbd ;
wire  kcd ;
wire  LBC ;
wire  LBD ;
wire  LCD ;
wire  MAA ;
wire  MAB ;
wire  MAC ;
wire  MBA ;
wire  MBB ;
wire  MBC ;
wire  MCA ;
wire  MCB ;
wire  MCC ;
wire  MDA ;
wire  MDB ;
wire  MDC ;
wire  NBA ;
wire  NBB ;
wire  NBC ;
wire  NCA ;
wire  NCB ;
wire  NCC ;
wire  NDA ;
wire  NDB ;
wire  NDC ;
wire  oaa ;
wire  oab ;
wire  oac ;
wire  oad ;
wire  oae ;
wire  oaf ;
wire  oag ;
wire  oah ;
wire  oai ;
wire  oaj ;
wire  oak ;
wire  oal ;
wire  oam ;
wire  oan ;
wire  oao ;
wire  oap ;
wire  oba ;
wire  obb ;
wire  obc ;
wire  obd ;
wire  obe ;
wire  obf ;
wire  obg ;
wire  obh ;
wire  obi ;
wire  obj ;
wire  obk ;
wire  obl ;
wire  obm ;
wire  obn ;
wire  obo ;
wire  obp ;
wire  oca ;
wire  ocb ;
wire  occ ;
wire  ocd ;
wire  oce ;
wire  ocf ;
wire  ocg ;
wire  och ;
wire  oci ;
wire  ocj ;
wire  ock ;
wire  ocl ;
wire  ocm ;
wire  ocn ;
wire  oco ;
wire  ocp ;
wire  oda ;
wire  odb ;
wire  odc ;
wire  odd ;
wire  ode ;
wire  odf ;
wire  odg ;
wire  odh ;
wire  odi ;
wire  odj ;
wire  odk ;
wire  odl ;
wire  odm ;
wire  odn ;
wire  odo ;
wire  odp ;
wire  pab ;
wire  PAB ;
wire  pac ;
wire  PAC ;
wire  pad ;
wire  PAD ;
wire  pba ;
wire  PBA ;
wire  pbb ;
wire  PBB ;
wire  pbc ;
wire  PBC ;
wire  pbd ;
wire  PBD ;
wire  pca ;
wire  PCA ;
wire  pcb ;
wire  PCB ;
wire  pcc ;
wire  PCC ;
wire  pcd ;
wire  PCD ;
wire  pda ;
wire  PDA ;
wire  pdb ;
wire  PDB ;
wire  pdc ;
wire  PDC ;
wire  pdd ;
wire  PDD ;
wire  QAA ;
wire  qab ;
wire  qac ;
wire  qad ;
wire  QBA ;
wire  QBB ;
wire  QBC ;
wire  QBD ;
wire  QBE ;
wire  qca ;
wire  QCB ;
wire  QCC ;
wire  QCD ;
wire  QCE ;
wire  qda ;
wire  qdb ;
wire  qdc ;
wire  qdd ;
wire  qde ;
wire  QDF ;
wire  qea ;
wire  qec ;
wire  qed ;
wire  qee ;
wire  qef ;
wire  QEG ;
wire  qfc ;
wire  qfe ;
wire  raa ;
wire  rab ;
wire  rac ;
wire  rad ;
wire  rae ;
wire  RAF ;
wire  rba ;
wire  rbb ;
wire  rbc ;
wire  rbd ;
wire  rbe ;
wire  RBF ;
wire  rca ;
wire  rcb ;
wire  rcc ;
wire  rcd ;
wire  rce ;
wire  RCF ;
wire  rda ;
wire  rdb ;
wire  rdc ;
wire  rdd ;
wire  rde ;
wire  RDF ;
wire  REA ;
wire  REB ;
wire  REC ;
wire  RED ;
wire  REE ;
wire  RFA ;
wire  RFB ;
wire  RFC ;
wire  RFD ;
wire  RFE ;
wire  RGA ;
wire  RGB ;
wire  RGC ;
wire  RGD ;
wire  RGE ;
wire  RHA ;
wire  RHB ;
wire  RHC ;
wire  RHD ;
wire  RHE ;
wire  rma ;
wire  rmb ;
wire  rmc ;
wire  rmd ;
wire  RME ;
wire  RMF ;
wire  rmg ;
wire  saa ;
wire  sab ;
wire  sac ;
wire  SBA ;
wire  SBB ;
wire  SBC ;
wire  sbd ;
wire  sbe ;
wire  sbf ;
wire  sbg ;
wire  sbh ;
wire  sbi ;
wire  sbj ;
wire  sbk ;
wire  SCA ;
wire  SCB ;
wire  SCC ;
wire  SCD ;
wire  SCE ;
wire  SCF ;
wire  scg ;
wire  sch ;
wire  SDA ;
wire  SWA ;
wire  SWB ;
wire  SWC ;
wire  SWD ;
wire  SWE ;
wire  SWF ;
wire  SWG ;
wire  SWH ;
wire  SWI ;
wire  SWJ ;
wire  SWK ;
wire  SWL ;
wire  SWM ;
wire  SWN ;
wire  SWO ;
wire  SWP ;
wire  SXA ;
wire  SXB ;
wire  SXC ;
wire  SXD ;
wire  SXE ;
wire  SXF ;
wire  SXG ;
wire  SXH ;
wire  SXI ;
wire  SXJ ;
wire  SXK ;
wire  SXL ;
wire  SXM ;
wire  SXN ;
wire  SXO ;
wire  SXP ;
wire  SYA ;
wire  SYB ;
wire  SYC ;
wire  SYD ;
wire  SYE ;
wire  SYF ;
wire  SYG ;
wire  SYH ;
wire  SYI ;
wire  SYJ ;
wire  SYK ;
wire  SYL ;
wire  SYM ;
wire  SYN ;
wire  SYO ;
wire  SYP ;
wire  SZA ;
wire  SZB ;
wire  SZC ;
wire  SZD ;
wire  SZE ;
wire  SZF ;
wire  SZG ;
wire  SZH ;
wire  SZI ;
wire  SZJ ;
wire  SZK ;
wire  SZL ;
wire  SZM ;
wire  SZN ;
wire  SZO ;
wire  SZP ;
wire  taa ;
wire  tab ;
wire  tac ;
wire  tad ;
wire  tae ;
wire  taf ;
wire  tag ;
wire  tah ;
wire  TBA ;
wire  TBB ;
wire  TBC ;
wire  TBD ;
wire  TBE ;
wire  TBF ;
wire  TBG ;
wire  TBH ;
wire  tca ;
wire  tcb ;
wire  tcc ;
wire  tcd ;
wire  tce ;
wire  tcf ;
wire  tcg ;
wire  tch ;
wire  tci ;
wire  tcj ;
wire  tck ;
wire  tcl ;
wire  tcm ;
wire  tcn ;
wire  tco ;
wire  tcp ;
wire  tda ;
wire  tdb ;
wire  tdc ;
wire  tdd ;
wire  tde ;
wire  tdf ;
wire  tdg ;
wire  tdh ;
wire  tea ;
wire  teb ;
wire  tec ;
wire  tfa ;
wire  tfb ;
wire  uaa ;
wire  UAA ;
wire  uba ;
wire  UBA ;
wire  ubb ;
wire  UBB ;
wire  ubc ;
wire  UBC ;
wire  ubd ;
wire  UBD ;
wire  uca ;
wire  UCA ;
wire  ucb ;
wire  UCB ;
wire  ucc ;
wire  UCC ;
wire  ucd ;
wire  UCD ;
wire  uce ;
wire  UCE ;
wire  ucf ;
wire  UCF ;
wire  uda ;
wire  UDA ;
wire  udb ;
wire  UDB ;
wire  udc ;
wire  UDC ;
wire  uea ;
wire  UEA ;
wire  vaa ;
wire  vba ;
wire  vbb ;
wire  VCA ;
wire  VCB ;
wire  vcc ;
wire  vcd ;
wire  VDA ;
wire  VDB ;
wire  vdc ;
wire  VEA ;
wire  veb ;
wire  VMA ;
wire  VMB ;
wire  VMC ;
wire  VMD ;
wire  VNA ;
wire  VNB ;
wire  VNC ;
wire  VND ;
wire  VOA ;
wire  VOB ;
wire  VOC ;
wire  VOD ;
wire  VPA ;
wire  VPB ;
wire  VPC ;
wire  VPD ;
wire  VQA ;
wire  VQB ;
wire  VQC ;
wire  VQD ;
wire  VRA ;
wire  VRB ;
wire  VRC ;
wire  VRD ;
wire  VSA ;
wire  VSB ;
wire  VSC ;
wire  VSD ;
wire  VTA ;
wire  VTB ;
wire  VTC ;
wire  VTD ;
wire  VUA ;
wire  VUB ;
wire  VUC ;
wire  VUD ;
wire  VVA ;
wire  VVB ;
wire  VVC ;
wire  VVD ;
wire  VWA ;
wire  VWB ;
wire  VWC ;
wire  VWD ;
wire  VXA ;
wire  VXB ;
wire  VXC ;
wire  VXD ;
wire  wca ;
wire  WCA ;
wire  wda ;
wire  WDA ;
wire  wdb ;
wire  WDB ;
wire  wea ;
wire  WEA ;
wire  web ;
wire  WEB ;
wire  wfa ;
wire  WFA ;
wire  wma ;
wire  WMA ;
wire  wmb ;
wire  WMB ;
wire  wmc ;
wire  WMC ;
wire  wpa ;
wire  WPA ;
wire  wpb ;
wire  WPB ;
wire  wpc ;
wire  WPC ;
wire  wsa ;
wire  WSA ;
wire  wsb ;
wire  WSB ;
wire  wsc ;
wire  WSC ;
wire  wva ;
wire  WVA ;
wire  wvb ;
wire  WVB ;
wire  wvc ;
wire  WVC ;
wire  xab ;
wire  xac ;
wire  xad ;
wire  xae ;
wire  XBA ;
wire  XBB ;
wire  XBC ;
wire  XBD ;
wire  XBE ;
wire  XBF ;
wire  xma ;
wire  xmb ;
wire  XMC ;
wire  XMD ;
wire  XME ;
wire  xpa ;
wire  xpb ;
wire  XPC ;
wire  XPD ;
wire  XPE ;
wire  xsa ;
wire  xsb ;
wire  XSC ;
wire  XSD ;
wire  XSE ;
wire  XSF ;
wire  xva ;
wire  xvb ;
wire  XVC ;
wire  XVD ;
wire  XVE ;
wire  XVF ;
wire  yac ;
wire  YAC ;
wire  yad ;
wire  YAD ;
wire  yae ;
wire  YAE ;
wire  yaf ;
wire  YAF ;
wire  yma ;
wire  YMA ;
wire  ymb ;
wire  YMB ;
wire  ymc ;
wire  YMC ;
wire  ymd ;
wire  YMD ;
wire  yme ;
wire  YME ;
wire  ZZI ;
wire  ZZO ;
assign ZZI = 1'b1;
assign ZZO = 1'b0;
assign rma = ~RMA;  //complement 
assign GAA = ~gaa;  //complement 
assign rmb = ~RMB;  //complement 
assign GAB = ~gab;  //complement 
assign VMA = ~vma;  //complement 
assign rmc = ~RMC;  //complement 
assign GAC = ~gac;  //complement 
assign VNA = ~vna;  //complement 
assign VOA = ~voa;  //complement 
assign rmd = ~RMD;  //complement 
assign GAD = ~gad;  //complement 
assign GIA = ~gia;  //complement 
assign HIA = ~hia;  //complement 
assign GIB = ~gib;  //complement 
assign HIB = ~hib;  //complement 
assign dib =  bia  ; 
assign DIB = ~dib;  //complement 
assign dic =  aib & bia  |  bib  ; 
assign DIC = ~dic;  //complement 
assign VSA = ~vsa;  //complement 
assign GIC = ~gic;  //complement 
assign HIC = ~hic;  //complement 
assign did =  bia & aib & aic  |  bib & aic  |  bic  ; 
assign DID = ~did; //complement 
assign VUA = ~vua;  //complement 
assign VTA = ~vta;  //complement 
assign GID = ~gid;  //complement 
assign HID = ~hid;  //complement 
assign tca = ~TCA;  //complement 
assign tda = ~TDA;  //complement 
assign taa = ~TAA;  //complement 
assign TBA = ~tba;  //complement 
assign EAA = TCA & ~AAA & ~BAA  |  ZZO & ~AAA & BAA  |  tca & AAA & ~BAA  |  TCA & AAA & BAA; 
assign eaa = ~EAA;  //complement 
assign EAB = TCA & ~AAB & ~BAB  |         ZZO & ~AAB & BAB  |  tca & AAB & ~BAB  |  TCA & AAB & BAB ; 
assign eab = ~EAB;  //complement 
assign CAB =  AAA  ; 
assign cab = ~CAB;  //complement 
assign CAC =  BAB & AAA  |  AAB  ; 
assign cac = ~CAC;  //complement 
assign EAC = TCA & ~AAC & ~BAC  |  ZZO & ~AAC & BAC  |  tca & AAC & ~BAC  |  TCA & AAC & BAC; 
assign eac = ~EAC;  //complement 
assign EAD = TCA & ~AAD & ~BAD  |         ZZO & ~AAD & BAD  |  tca & AAD & ~BAD  |  TCA & AAD & BAD ; 
assign ead = ~EAD;  //complement 
assign CAD =  AAA & BAB & BAC  |  AAB & BAC  |  AAC  ; 
assign cad = ~CAD; //complement 
assign CAE =  AAA & BAB & BAC & BAD  |  AAB & BAC & BAD  |  AAC & BAD  |  AAD  ; 
assign cae = ~CAE;  //complement 
assign FAI =  BIA & BIF & BIG & BID  ; 
assign fai = ~FAI;  //complement  
assign kab = ~KAB;  //complement 
assign PCA =  KAC & LBC  |  KBC  ; 
assign pca = ~PCA; //complement 
assign EIA = TCI & ~AIA & ~BIA  |  ZZO & ~AIA & BIA  |  tci & AIA & ~BIA  |  TCI & AIA & BIA; 
assign eia = ~EIA;  //complement 
assign EIB = TCI & ~AIB & ~BIB  |         ZZO & ~AIB & BIB  |  tci & AIB & ~BIB  |  TCI & AIB & BIB ; 
assign eib = ~EIB;  //complement 
assign CIB =  AIA  ; 
assign cib = ~CIB;  //complement 
assign CIC =  BIB & AIA  |  AIB  ; 
assign cic = ~CIC;  //complement 
assign bib = ~BIB;  //complement 
assign bif = ~BIF;  //complement 
assign EIC = TCI & ~AIC & ~BIC  |  ZZO & ~AIC & BIC  |  tci & AIC & ~BIC  |  TCI & AIC & BIC; 
assign eic = ~EIC;  //complement 
assign EID = TCI & ~AID & ~BID  |         ZZO & ~AID & BID  |  tci & AID & ~BID  |  TCI & AID & BID ; 
assign eid = ~EID;  //complement 
assign CID =  AIA & BIB & BIC  |  AIB & BIC  |  AIC  ; 
assign cid = ~CID; //complement 
assign bic = ~BIC;  //complement 
assign big = ~BIG;  //complement 
assign tci = ~TCI;  //complement 
assign CIE =  AIA & BIB & BIC & BID  |  AIB & BIC & BID  |  AIC & BID  |  AID  ; 
assign cie = ~CIE;  //complement 
assign AAA = ~aaa;  //complement 
assign baa = ~BAA;  //complement 
assign AAB = ~aab;  //complement 
assign bab = ~BAB;  //complement 
assign oaa = ~OAA;  //complement 
assign YAC =  TEB & XAB & XAB  ; 
assign yac = ~YAC;  //complement 
assign YAD =  XBC & TEB & XAB  |  TEB & XAC  ; 
assign yad = ~YAD;  //complement 
assign JAA =  RAA & rab & rae  |  raa & RAB & rae  |  raa & rab & RAE  |  RAA & RAB & RAE  ; 
assign jaa = ~JAA; //complement 
assign jba =  RAA & rab & rae  |  raa & RAB & rae  |  raa & rab & RAE  |  raa & rab & rae  ; 
assign JBA = ~jba;  //complement 
assign AAC = ~aac;  //complement 
assign bac = ~BAC;  //complement 
assign oac = ~OAC;  //complement 
assign SWB = ~swb;  //complement 
assign SWC = ~swc;  //complement 
assign SWD = ~swd;  //complement 
assign raa = ~RAA;  //complement 
assign REA = ~rea;  //complement 
assign AAD = ~aad;  //complement 
assign bad = ~BAD;  //complement 
assign oad = ~OAD;  //complement 
assign saa = ~SAA;  //complement 
assign SBA = ~sba;  //complement 
assign AIA = ~aia;  //complement 
assign bia = ~BIA;  //complement 
assign AIB = ~aib;  //complement 
assign oca = ~OCA;  //complement 
assign ocb = ~OCB;  //complement 
assign JAE =  RCA & rcb & rce  |  rca & RCB & rce  |  rca & rcb & RCE  |  RCA & RCB & RCE  ; 
assign jae = ~JAE; //complement 
assign jbe =  RCA & rcb & rce  |  rca & RCB & rce  |  rca & rcb & RCE  |  rca & rcb & rce  ; 
assign JBE = ~jbe;  //complement 
assign AIC = ~aic;  //complement 
assign SYB = ~syb;  //complement 
assign SYC = ~syc;  //complement 
assign SYD = ~syd;  //complement 
assign rca = ~RCA;  //complement 
assign RGA = ~rga;  //complement 
assign AID = ~aid;  //complement 
assign bid = ~BID;  //complement 
assign occ = ~OCC;  //complement 
assign ocd = ~OCD;  //complement 
assign oab = ~OAB;  //complement 
assign XMC = ~xmc;  //complement 
assign RME = ~rme;  //complement 
assign RMF = ~rmf;  //complement 
assign GBA = ~gba;  //complement 
assign HBA = ~hba;  //complement 
assign XMD = ~xmd;  //complement 
assign XME = ~xme;  //complement 
assign GBB = ~gbb;  //complement 
assign HBB = ~hbb;  //complement 
assign dbb =  bba  ; 
assign DBB = ~dbb;  //complement 
assign dbc =  abb & bba  |  bbb  ; 
assign DBC = ~dbc;  //complement 
assign VMB = ~vmb;  //complement 
assign rmg = ~RMG;  //complement 
assign GBC = ~gbc;  //complement 
assign HBC = ~hbc;  //complement 
assign dbd =  bba & abb & abc  |  bbb & abc  |  bbc  ; 
assign DBD = ~dbd; //complement 
assign VOB = ~vob;  //complement 
assign YMB =  XVE & XSE & xpe  ; 
assign ymb = ~YMB;  //complement 
assign YMC =  XVE & xse  ; 
assign ymc = ~YMC;  //complement 
assign YMD =  xve & TFB  ; 
assign ymd = ~YMD;  //complement 
assign GBD = ~gbd;  //complement 
assign HBD = ~hbd;  //complement 
assign VNB = ~vnb;  //complement 
assign XSC = ~xsc;  //complement 
assign YMA =  XVF & XSF & XPE & xme  ; 
assign yma = ~YMA;  //complement  
assign YME =  XVF & XSF & XPE & XME  ; 
assign yme = ~YME;  //complement 
assign GJA = ~gja;  //complement 
assign HJA = ~hja;  //complement 
assign XSD = ~xsd;  //complement 
assign XSF = ~xsf;  //complement 
assign XSE = ~xse;  //complement 
assign GJB = ~gjb;  //complement 
assign HJB = ~hjb;  //complement 
assign djb =  bja  ; 
assign DJB = ~djb;  //complement 
assign djc =  ajb & bja  |  bjb  ; 
assign DJC = ~djc;  //complement 
assign VSB = ~vsb;  //complement 
assign VTB = ~vtb;  //complement 
assign GJC = ~gjc;  //complement 
assign HJC = ~hjc;  //complement 
assign djd =  bja & ajb & ajc  |  bjb & ajc  |  bjc  ; 
assign DJD = ~djd; //complement 
assign VUB = ~vub;  //complement 
assign GJD = ~gjd;  //complement 
assign HJD = ~hjd;  //complement 
assign tcb = ~TCB;  //complement 
assign tdb = ~TDB;  //complement 
assign tab = ~TAB;  //complement 
assign TBB = ~tbb;  //complement 
assign MAA = ~maa;  //complement 
assign EBA = TCB & ~ABA & ~BBA  |  ZZO & ~ABA & BBA  |  tcb & ABA & ~BBA  |  TCB & ABA & BBA; 
assign eba = ~EBA;  //complement 
assign EBB = TCB & ~ABB & ~BBB  |         ZZO & ~ABB & BBB  |  tcb & ABB & ~BBB  |  TCB & ABB & BBB ; 
assign ebb = ~EBB;  //complement 
assign CBB =  ABA  ; 
assign cbb = ~CBB;  //complement 
assign CBC =  BBB & ABA  |  ABB  ; 
assign cbc = ~CBC;  //complement 
assign bbb = ~BBB;  //complement 
assign bbf = ~BBF;  //complement 
assign EBC = TCB & ~ABC & ~BBC  |  ZZO & ~ABC & BBC  |  tcb & ABC & ~BBC  |  TCB & ABC & BBC; 
assign ebc = ~EBC;  //complement 
assign EBD = TCB & ~ABD & ~BBD  |         ZZO & ~ABD & BBD  |  tcb & ABD & ~BBD  |  TCB & ABD & BBD ; 
assign ebd = ~EBD;  //complement 
assign CBD =  ABA & BBB & BBC  |  ABB & BBC  |  ABC  ; 
assign cbd = ~CBD; //complement 
assign bbc = ~BBC;  //complement 
assign bbg = ~BBG;  //complement 
assign FAB =  BBA & BBF & BBG & BBD  ; 
assign fab = ~FAB;  //complement  
assign CBE =  ABA & BBB & BBC & BBD  |  ABB & BBC & BBD  |  ABC & BBD  |  ABD  ; 
assign cbe = ~CBE;  //complement 
assign PAB =  MAA  ; 
assign pab = ~PAB;  //complement 
assign NCA = ~nca;  //complement 
assign FAJ =  BJA & BJF & BJG & BJD  ; 
assign faj = ~FAJ;  //complement  
assign FBJ =  BJA & BJF & BJG & BJD  ; 
assign fbj = ~FBJ;  //complement 
assign kac = ~KAC;  //complement 
assign PCB =  KAC & LBC & NCA  |  KBC & NCA  |  MCA  ; 
assign pcb = ~PCB; //complement 
assign EJA = TCJ & ~AJA & ~BJA  |  ZZO & ~AJA & BJA  |  tcj & AJA & ~BJA  |  TCJ & AJA & BJA; 
assign eja = ~EJA;  //complement 
assign EJB = TCJ & ~AJB & ~BJB  |         ZZO & ~AJB & BJB  |  tcj & AJB & ~BJB  |  TCJ & AJB & BJB ; 
assign ejb = ~EJB;  //complement 
assign CJB =  AJA  ; 
assign cjb = ~CJB;  //complement 
assign CJC =  BJB & AJA  |  AJB  ; 
assign cjc = ~CJC;  //complement 
assign bjb = ~BJB;  //complement 
assign bjf = ~BJF;  //complement 
assign EJC = TCJ & ~AJC & ~BJC  |  ZZO & ~AJC & BJC  |  tcj & AJC & ~BJC  |  TCJ & AJC & BJC; 
assign ejc = ~EJC;  //complement 
assign EJD = TCJ & ~AJD & ~BJD  |         ZZO & ~AJD & BJD  |  tcj & AJD & ~BJD  |  TCJ & AJD & BJD ; 
assign ejd = ~EJD;  //complement 
assign CJD =  AJA & BJB & BJC  |  AJB & BJC  |  AJC  ; 
assign cjd = ~CJD; //complement 
assign bjc = ~BJC;  //complement 
assign bjg = ~BJG;  //complement 
assign tcj = ~TCJ;  //complement 
assign CJE =  AJA & BJB & BJC & BJD  |  AJB & BJC & BJD  |  AJC & BJD  |  AJD  ; 
assign cje = ~CJE;  //complement 
assign MCA = ~mca;  //complement 
assign ABA = ~aba;  //complement 
assign bba = ~BBA;  //complement 
assign oae = ~OAE;  //complement 
assign SWA = ~swa;  //complement 
assign SWE = ~swe;  //complement 
assign SWI = ~swi;  //complement 
assign rae = ~RAE;  //complement 
assign REE = ~ree;  //complement 
assign ABB = ~abb;  //complement 
assign oaf = ~OAF;  //complement 
assign YAE =  XAB & XBC & XBD & TEB  |  XAC & XBD & TEB  |  XAD & TEB  ; 
assign yae = ~YAE;  //complement 
assign sbd = ~SBD;  //complement 
assign SCA = ~sca;  //complement 
assign ABC = ~abc;  //complement 
assign oag = ~OAG;  //complement 
assign SWF = ~swf;  //complement 
assign SWG = ~swg;  //complement 
assign SWH = ~swh;  //complement 
assign rab = ~RAB;  //complement 
assign REB = ~reb;  //complement 
assign ABD = ~abd;  //complement 
assign bbd = ~BBD;  //complement 
assign oah = ~OAH;  //complement 
assign UBB =  SBA & sbd & sbg  |  sba & SBD & sbg  |  sba & sbd & SBG  |  SBA & SBD & SBG  ; 
assign ubb = ~UBB; //complement 
assign uca =  SBA & sbd & sbg  |  sba & SBD & sbg  |  sba & sbd & SBG  |  sba & sbd & sbg  ; 
assign UCA = ~uca;  //complement 
assign UCF =  sca & SCD & SCD  |  SCA & scd  ; 
assign ucf = ~UCF;  //complement 
assign UEA =  SCA & SDA & SCD  ; 
assign uea = ~UEA;  //complement 
assign AJA = ~aja;  //complement 
assign bja = ~BJA;  //complement 
assign SYA = ~sya;  //complement 
assign SYE = ~sye;  //complement 
assign SYI = ~syi;  //complement 
assign rce = ~RCE;  //complement 
assign RGE = ~rge;  //complement 
assign AJB = ~ajb;  //complement 
assign oce = ~OCE;  //complement 
assign ocf = ~OCF;  //complement 
assign vcc = ~VCC;  //complement 
assign VDA = ~vda;  //complement 
assign sbg = ~SBG;  //complement 
assign SCD = ~scd;  //complement 
assign AJC = ~ajc;  //complement 
assign SYF = ~syf;  //complement 
assign SYG = ~syg;  //complement 
assign SYH = ~syh;  //complement 
assign rcb = ~RCB;  //complement 
assign RGB = ~rgb;  //complement 
assign AJD = ~ajd;  //complement 
assign bjd = ~BJD;  //complement 
assign ocg = ~OCG;  //complement 
assign och = ~OCH;  //complement 
assign GCA = ~gca;  //complement 
assign HCA = ~hca;  //complement 
assign xma = ~XMA;  //complement 
assign xmb = ~XMB;  //complement 
assign GCB = ~gcb;  //complement 
assign HCB = ~hcb;  //complement 
assign dcb =  bca  ; 
assign DCB = ~dcb;  //complement 
assign dcc =  acb & bca  |  bcb  ; 
assign DCC = ~dcc;  //complement 
assign VMC = ~vmc;  //complement 
assign WMA =  VMB & VMC & VMD  ; 
assign wma = ~WMA;  //complement 
assign WMB =  vmb & VMC & VMD  ; 
assign wmb = ~WMB;  //complement 
assign WMC =  vmc & VMD & VMD  ; 
assign wmc = ~WMC;  //complement 
assign GCC = ~gcc;  //complement 
assign HCC = ~hcc;  //complement 
assign dcd =  bca & acb & acc  |  bcb & acc  |  bcc  ; 
assign DCD = ~dcd; //complement 
assign VOC = ~voc;  //complement 
assign GCD = ~gcd;  //complement 
assign HCD = ~hcd;  //complement 
assign VNC = ~vnc;  //complement 
assign GKA = ~gka;  //complement 
assign HKA = ~hka;  //complement 
assign xsa = ~XSA;  //complement 
assign xsb = ~XSB;  //complement 
assign GKB = ~gkb;  //complement 
assign HKB = ~hkb;  //complement 
assign dkb =  bka  ; 
assign DKB = ~dkb;  //complement 
assign dkc =  akb & bka  |  bkb  ; 
assign DKC = ~dkc;  //complement 
assign VSC = ~vsc;  //complement 
assign WSA =  VSB & VSC & VSD  ; 
assign wsa = ~WSA;  //complement 
assign WSB =  vsb & VSC & VSD  ; 
assign wsb = ~WSB;  //complement 
assign WSC =  vsc & VSD & VSD  ; 
assign wsc = ~WSC;  //complement 
assign GKC = ~gkc;  //complement 
assign HKC = ~hkc;  //complement 
assign dkd =  bka & akb & akc  |  bkb & akc  |  bkc  ; 
assign DKD = ~dkd; //complement 
assign VUC = ~vuc;  //complement 
assign VTC = ~vtc;  //complement 
assign GKD = ~gkd;  //complement 
assign HKD = ~hkd;  //complement 
assign tcc = ~TCC;  //complement 
assign tdc = ~TDC;  //complement 
assign tac = ~TAC;  //complement 
assign TBC = ~tbc;  //complement 
assign MAB = ~mab;  //complement 
assign ECA = TCC & ~ACA & ~BCA  |  ZZO & ~ACA & BCA  |  tcc & ACA & ~BCA  |  TCC & ACA & BCA; 
assign eca = ~ECA;  //complement 
assign ECB = TCC & ~ACB & ~BCB  |         ZZO & ~ACB & BCB  |  tcc & ACB & ~BCB  |  TCC & ACB & BCB ; 
assign ecb = ~ECB;  //complement 
assign CCB =  ACA  ; 
assign ccb = ~CCB;  //complement 
assign CCC =  BCB & ACA  |  ACB  ; 
assign ccc = ~CCC;  //complement 
assign bcb = ~BCB;  //complement 
assign bcf = ~BCF;  //complement 
assign ECC = TCC & ~ACC & ~BCC  |  ZZO & ~ACC & BCC  |  tcc & ACC & ~BCC  |  TCC & ACC & BCC; 
assign ecc = ~ECC;  //complement 
assign ECD = TCC & ~ACD & ~BCD  |         ZZO & ~ACD & BCD  |  tcc & ACD & ~BCD  |  TCC & ACD & BCD ; 
assign ecd = ~ECD;  //complement 
assign CCD =  ACA & BCB & BCC  |  ACB & BCC  |  ACC  ; 
assign ccd = ~CCD; //complement 
assign bcc = ~BCC;  //complement 
assign bcg = ~BCG;  //complement 
assign FAC =  BCA & BCF & BCG & BCD  ; 
assign fac = ~FAC;  //complement  
assign CCE =  ACA & BCB & BCC & BCD  |  ACB & BCC & BCD  |  ACC & BCD  |  ACD  ; 
assign cce = ~CCE;  //complement 
assign PAC =  MAB  ; 
assign pac = ~PAC;  //complement 
assign NCB = ~ncb;  //complement 
assign FAK =  BKA & BKF & BKG & BKD  ; 
assign fak = ~FAK;  //complement  
assign FBK =  BKA & BKF & BKG & BKD  ; 
assign fbk = ~FBK;  //complement 
assign kad = ~KAD;  //complement 
assign PCC =  KAC & LBC & NCB  |  KBC & NCB  |  MCB  ; 
assign pcc = ~PCC; //complement 
assign EKA = TCK & ~AKA & ~BKA  |  ZZO & ~AKA & BKA  |  tck & AKA & ~BKA  |  TCK & AKA & BKA; 
assign eka = ~EKA;  //complement 
assign EKB = TCK & ~AKB & ~BKB  |         ZZO & ~AKB & BKB  |  tck & AKB & ~BKB  |  TCK & AKB & BKB ; 
assign ekb = ~EKB;  //complement 
assign CKB =  AKA  ; 
assign ckb = ~CKB;  //complement 
assign CKC =  BKB & AKA  |  AKB  ; 
assign ckc = ~CKC;  //complement 
assign bkb = ~BKB;  //complement 
assign bkf = ~BKF;  //complement 
assign EKC = TCK & ~AKC & ~BKC  |  ZZO & ~AKC & BKC  |  tck & AKC & ~BKC  |  TCK & AKC & BKC; 
assign ekc = ~EKC;  //complement 
assign EKD = TCK & ~AKD & ~BKD  |         ZZO & ~AKD & BKD  |  tck & AKD & ~BKD  |  TCK & AKD & BKD ; 
assign ekd = ~EKD;  //complement 
assign CKD =  AKA & BKB & BKC  |  AKB & BKC  |  AKC  ; 
assign ckd = ~CKD; //complement 
assign bkc = ~BKC;  //complement 
assign bkg = ~BKG;  //complement 
assign tck = ~TCK;  //complement 
assign CKE =  AKA & BKB & BKC & BKD  |  AKB & BKC & BKD  |  AKC & BKD  |  AKD  ; 
assign cke = ~CKE;  //complement 
assign MCB = ~mcb;  //complement 
assign ACA = ~aca;  //complement 
assign bca = ~BCA;  //complement 
assign ACB = ~acb;  //complement 
assign oai = ~OAI;  //complement 
assign oaj = ~OAJ;  //complement 
assign YAF =  XAB & XBC & XBD & XBE & TEB  |  XAC & XBD & XBE & TEB  |  XAD & XBE & TEB  |  XAE & TEB  ; 
assign yaf = ~YAF;  //complement 
assign JAB =  RAC & rad & raf  |  rac & RAD & raf  |  rac & rad & RAF  |  RAC & RAD & RAF  ; 
assign jab = ~JAB; //complement 
assign jbb =  RAC & rad & raf  |  rac & RAD & raf  |  rac & rad & RAF  |  rac & rad & raf  ; 
assign JBB = ~jbb;  //complement 
assign ACC = ~acc;  //complement 
assign SWJ = ~swj;  //complement 
assign SWK = ~swk;  //complement 
assign SWL = ~swl;  //complement 
assign rac = ~RAC;  //complement 
assign REC = ~rec;  //complement 
assign sbj = ~SBJ;  //complement 
assign ACD = ~acd;  //complement 
assign bcd = ~BCD;  //complement 
assign oak = ~OAK;  //complement 
assign oal = ~OAL;  //complement 
assign WEB =  VEA & veb  |  VEB & vea  ; 
assign web = ~WEB;  //complement 
assign wfa =  veb  |  vea  ; 
assign WFA = ~wfa;  //complement 
assign UDC =  SCA & SCD & sda  |  sca & SDA  |  scd & SDA  ; 
assign udc = ~UDC; //complement 
assign AKA = ~aka;  //complement 
assign bka = ~BKA;  //complement 
assign vba = ~VBA;  //complement 
assign VCA = ~vca;  //complement 
assign AKB = ~akb;  //complement 
assign oci = ~OCI;  //complement 
assign ocj = ~OCJ;  //complement 
assign vdc = ~VDC;  //complement 
assign VEA = ~vea;  //complement 
assign veb = ~VEB;  //complement 
assign JAF =  RCC & rcd & rcf  |  rcc & RCD & rcf  |  rcc & rcd & RCF  |  RCC & RCD & RCF  ; 
assign jaf = ~JAF; //complement 
assign jbf =  RCC & rcd & rcf  |  rcc & RCD & rcf  |  rcc & rcd & RCF  |  rcc & rcd & rcf  ; 
assign JBF = ~jbf;  //complement 
assign AKC = ~akc;  //complement 
assign SYJ = ~syj;  //complement 
assign SYK = ~syk;  //complement 
assign SYL = ~syl;  //complement 
assign rcc = ~RCC;  //complement 
assign RGC = ~rgc;  //complement 
assign sbk = ~SBK;  //complement 
assign AKD = ~akd;  //complement 
assign bkd = ~BKD;  //complement 
assign ock = ~OCK;  //complement 
assign ocl = ~OCL;  //complement 
assign GDA = ~gda;  //complement 
assign HDA = ~hda;  //complement 
assign GDB = ~gdb;  //complement 
assign HDB = ~hdb;  //complement 
assign ddb =  bda  ; 
assign DDB = ~ddb;  //complement 
assign ddc =  adb & bda  |  bdb  ; 
assign DDC = ~ddc;  //complement 
assign VMD = ~vmd;  //complement 
assign GDC = ~gdc;  //complement 
assign HDC = ~hdc;  //complement 
assign ddd =  bda & adb & adc  |  bdb & adc  |  bdc  ; 
assign DDD = ~ddd; //complement 
assign VOD = ~vod;  //complement 
assign GDD = ~gdd;  //complement 
assign HDD = ~hdd;  //complement 
assign VND = ~vnd;  //complement 
assign GLA = ~gla;  //complement 
assign HLA = ~hla;  //complement 
assign GLB = ~glb;  //complement 
assign HLB = ~hlb;  //complement 
assign dlb =  bla  ; 
assign DLB = ~dlb;  //complement 
assign dlc =  alb & bla  |  blb  ; 
assign DLC = ~dlc;  //complement 
assign VSD = ~vsd;  //complement 
assign GLC = ~glc;  //complement 
assign HLC = ~hlc;  //complement 
assign dld =  bla & alb & alc  |  blb & alc  |  blc  ; 
assign DLD = ~dld; //complement 
assign VUD = ~vud;  //complement 
assign VTD = ~vtd;  //complement 
assign GLD = ~gld;  //complement 
assign HLD = ~hld;  //complement 
assign tcd = ~TCD;  //complement 
assign tdd = ~TDD;  //complement 
assign tad = ~TAD;  //complement 
assign TBD = ~tbd;  //complement 
assign MAC = ~mac;  //complement 
assign EDA = TCD & ~ADA & ~BDA  |  ZZO & ~ADA & BDA  |  tcd & ADA & ~BDA  |  TCD & ADA & BDA; 
assign eda = ~EDA;  //complement 
assign EDB = TCD & ~ADB & ~BDB  |         ZZO & ~ADB & BDB  |  tcd & ADB & ~BDB  |  TCD & ADB & BDB ; 
assign edb = ~EDB;  //complement 
assign CDB =  ADA  ; 
assign cdb = ~CDB;  //complement 
assign CDC =  BDB & ADA  |  ADB  ; 
assign cdc = ~CDC;  //complement 
assign bdb = ~BDB;  //complement 
assign bdf = ~BDF;  //complement 
assign EDC = TCD & ~ADC & ~BDC  |  ZZO & ~ADC & BDC  |  tcd & ADC & ~BDC  |  TCD & ADC & BDC; 
assign edc = ~EDC;  //complement 
assign EDD = TCD & ~ADD & ~BDD  |         ZZO & ~ADD & BDD  |  tcd & ADD & ~BDD  |  TCD & ADD & BDD ; 
assign edd = ~EDD;  //complement 
assign CDD =  ADA & BDB & BDC  |  ADB & BDC  |  ADC  ; 
assign cdd = ~CDD; //complement 
assign bdc = ~BDC;  //complement 
assign bdg = ~BDG;  //complement 
assign FAD =  BDA & BDF & BDG & BDD  ; 
assign fad = ~FAD;  //complement  
assign CDE =  ADA & BDB & BDC & BDD  |  ADB & BDC & BDD  |  ADC & BDD  |  ADD  ; 
assign cde = ~CDE;  //complement 
assign PAD =  MAC  ; 
assign pad = ~PAD;  //complement 
assign NCC = ~ncc;  //complement 
assign FAL =  BLA & BLF & BLG & BLD  ; 
assign fal = ~FAL;  //complement  
assign kbc = ~KBC;  //complement 
assign PCD =  KAC & LBC & NCC  |  KBC & NCC  |  MCC  ; 
assign pcd = ~PCD; //complement 
assign ELA = TCL & ~ALA & ~BLA  |  ZZO & ~ALA & BLA  |  tcl & ALA & ~BLA  |  TCL & ALA & BLA; 
assign ela = ~ELA;  //complement 
assign ELB = TCL & ~ALB & ~BLB  |         ZZO & ~ALB & BLB  |  tcl & ALB & ~BLB  |  TCL & ALB & BLB ; 
assign elb = ~ELB;  //complement 
assign CLB =  ALA  ; 
assign clb = ~CLB;  //complement 
assign CLC =  BLB & ALA  |  ALB  ; 
assign clc = ~CLC;  //complement 
assign blb = ~BLB;  //complement 
assign blf = ~BLF;  //complement 
assign ELC = TCL & ~ALC & ~BLC  |  ZZO & ~ALC & BLC  |  tcl & ALC & ~BLC  |  TCL & ALC & BLC; 
assign elc = ~ELC;  //complement 
assign ELD = TCL & ~ALD & ~BLD  |         ZZO & ~ALD & BLD  |  tcl & ALD & ~BLD  |  TCL & ALD & BLD ; 
assign eld = ~ELD;  //complement 
assign CLD =  ALA & BLB & BLC  |  ALB & BLC  |  ALC  ; 
assign cld = ~CLD; //complement 
assign blc = ~BLC;  //complement 
assign blg = ~BLG;  //complement 
assign tcl = ~TCL;  //complement 
assign CLE =  ALA & BLB & BLC & BLD  |  ALB & BLC & BLD  |  ALC & BLD  |  ALD  ; 
assign cle = ~CLE;  //complement 
assign MCC = ~mcc;  //complement 
assign ADA = ~ada;  //complement 
assign bda = ~BDA;  //complement 
assign XBF = ~xbf;  //complement 
assign XBB = ~xbb;  //complement 
assign RAF = ~raf;  //complement 
assign SWM = ~swm;  //complement 
assign ADB = ~adb;  //complement 
assign oam = ~OAM;  //complement 
assign oan = ~OAN;  //complement 
assign XBC = ~xbc;  //complement 
assign sbe = ~SBE;  //complement 
assign SCB = ~scb;  //complement 
assign ADC = ~adc;  //complement 
assign xab = ~XAB;  //complement 
assign SWN = ~swn;  //complement 
assign SWO = ~swo;  //complement 
assign SWP = ~swp;  //complement 
assign rad = ~RAD;  //complement 
assign RED = ~red;  //complement 
assign ADD = ~add;  //complement 
assign bdd = ~BDD;  //complement 
assign oao = ~OAO;  //complement 
assign oap = ~OAP;  //complement 
assign WCA =  VCA & vcb & vcc  |  vca & VCB & vcc  |  vca & vcb & VCC  |  VCA & VCB & VCC  ; 
assign wca = ~WCA; //complement 
assign wda =  VCA & vcb & vcc  |  vca & VCB & vcc  |  vca & vcb & VCC  |  vca & vcb & vcc  ; 
assign WDA = ~wda;  //complement 
assign JBI =  REB & rec & red  |  reb & REC & red  |  reb & rec & RED  |  REB & REC & RED  ; 
assign jbi = ~JBI; //complement 
assign jca =  REB & rec & red  |  reb & REC & red  |  reb & rec & RED  |  reb & rec & red  ; 
assign JCA = ~jca;  //complement 
assign ALA = ~ala;  //complement 
assign bla = ~BLA;  //complement 
assign xac = ~XAC;  //complement 
assign RCF = ~rcf;  //complement 
assign SYM = ~sym;  //complement 
assign XBA = ~xba;  //complement 
assign ALB = ~alb;  //complement 
assign ocm = ~OCM;  //complement 
assign ocn = ~OCN;  //complement 
assign UCD =  SCB & sce & scg  |  scb & SCE & scg  |  scb & sce & SCG  |  SCB & SCE & SCG  ; 
assign ucd = ~UCD; //complement 
assign uda =  SCB & sce & scg  |  scb & SCE & scg  |  scb & sce & SCG  |  scb & sce & scg  ; 
assign UDA = ~uda;  //complement 
assign scg = ~SCG;  //complement 
assign SDA = ~sda;  //complement 
assign ALC = ~alc;  //complement 
assign SYN = ~syn;  //complement 
assign SYO = ~syo;  //complement 
assign SYP = ~syp;  //complement 
assign rcd = ~RCD;  //complement 
assign RGD = ~rgd;  //complement 
assign ALD = ~ald;  //complement 
assign bld = ~BLD;  //complement 
assign oco = ~OCO;  //complement 
assign ocp = ~OCP;  //complement 
assign JBK =  RGB & rgc & rgd  |  rgb & RGC & rgd  |  rgb & rgc & RGD  |  RGB & RGC & RGD  ; 
assign jbk = ~JBK; //complement 
assign jcc =  RGB & rgc & rgd  |  rgb & RGC & rgd  |  rgb & rgc & RGD  |  rgb & rgc & rgd  ; 
assign JCC = ~jcc;  //complement 
assign GEA = ~gea;  //complement 
assign HEA = ~hea;  //complement 
assign GEB = ~geb;  //complement 
assign HEB = ~heb;  //complement 
assign deb =  bea  ; 
assign DEB = ~deb;  //complement 
assign dec =  aeb & bea  |  beb  ; 
assign DEC = ~dec;  //complement 
assign VPA = ~vpa;  //complement 
assign GEC = ~gec;  //complement 
assign HEC = ~hec;  //complement 
assign ded =  bea & aeb & aec  |  beb & aec  |  bec  ; 
assign DED = ~ded; //complement 
assign VRA = ~vra;  //complement 
assign GED = ~ged;  //complement 
assign HED = ~hed;  //complement 
assign VQA = ~vqa;  //complement 
assign GMA = ~gma;  //complement 
assign HMA = ~hma;  //complement 
assign GMB = ~gmb;  //complement 
assign HMB = ~hmb;  //complement 
assign dmb =  bma  ; 
assign DMB = ~dmb;  //complement 
assign dmc =  amb & bma  |  bmb  ; 
assign DMC = ~dmc;  //complement 
assign VVA = ~vva;  //complement 
assign GMC = ~gmc;  //complement 
assign HMC = ~hmc;  //complement 
assign dmd =  bma & amb & amc  |  bmb & amc  |  bmc  ; 
assign DMD = ~dmd; //complement 
assign VXA = ~vxa;  //complement 
assign VWA = ~vwa;  //complement 
assign GMD = ~gmd;  //complement 
assign HMD = ~hmd;  //complement 
assign tce = ~TCE;  //complement 
assign tde = ~TDE;  //complement 
assign tae = ~TAE;  //complement 
assign TBE = ~tbe;  //complement 
assign EEA = TCE & ~AEA & ~BEA  |  ZZO & ~AEA & BEA  |  tce & AEA & ~BEA  |  TCE & AEA & BEA; 
assign eea = ~EEA;  //complement 
assign EEB = TCE & ~AEB & ~BEB  |         ZZO & ~AEB & BEB  |  tce & AEB & ~BEB  |  TCE & AEB & BEB ; 
assign eeb = ~EEB;  //complement 
assign CEB =  AEA  ; 
assign ceb = ~CEB;  //complement 
assign CEC =  BEB & AEA  |  AEB  ; 
assign cec = ~CEC;  //complement 
assign beb = ~BEB;  //complement 
assign bef = ~BEF;  //complement 
assign EEC = TCE & ~AEC & ~BEC  |  ZZO & ~AEC & BEC  |  tce & AEC & ~BEC  |  TCE & AEC & BEC; 
assign eec = ~EEC;  //complement 
assign EED = TCE & ~AED & ~BED  |         ZZO & ~AED & BED  |  tce & AED & ~BED  |  TCE & AED & BED ; 
assign eed = ~EED;  //complement 
assign CED =  AEA & BEB & BEC  |  AEB & BEC  |  AEC  ; 
assign ced = ~CED; //complement 
assign bec = ~BEC;  //complement 
assign beg = ~BEG;  //complement 
assign FAE =  BEA & BEF & BEG & BED  ; 
assign fae = ~FAE;  //complement  
assign CEE =  AEA & BEB & BEC & BED  |  AEB & BEC & BED  |  AEC & BED  |  AED  ; 
assign cee = ~CEE;  //complement 
assign pba =  kab  ; 
assign PBA = ~pba;  //complement 
assign FAM =  BMA & BMF & BMG & BMD  ; 
assign fam = ~FAM;  //complement  
assign kbd = ~KBD;  //complement 
assign PDA =  KAD & LBD & LCD  |  KBD & LCD  |  KCD  ; 
assign pda = ~PDA;  //complement 
assign EMA = TCM & ~AMA & ~BMA  |  ZZO & ~AMA & BMA  |  tcm & AMA & ~BMA  |  TCM & AMA & BMA; 
assign ema = ~EMA;  //complement 
assign EMB = TCM & ~AMB & ~BMB  |         ZZO & ~AMB & BMB  |  tcm & AMB & ~BMB  |  TCM & AMB & BMB ; 
assign emb = ~EMB;  //complement 
assign CMB =  AMA  ; 
assign cmb = ~CMB;  //complement 
assign CMC =  BMB & AMA  |  AMB  ; 
assign cmc = ~CMC;  //complement 
assign bmb = ~BMB;  //complement 
assign bmf = ~BMF;  //complement 
assign EMC = TCM & ~AMC & ~BMC  |  ZZO & ~AMC & BMC  |  tcm & AMC & ~BMC  |  TCM & AMC & BMC; 
assign emc = ~EMC;  //complement 
assign EMD = TCM & ~AMD & ~BMD  |         ZZO & ~AMD & BMD  |  tcm & AMD & ~BMD  |  TCM & AMD & BMD ; 
assign emd = ~EMD;  //complement 
assign CMD =  AMA & BMB & BMC  |  AMB & BMC  |  AMC  ; 
assign cmd = ~CMD; //complement 
assign bmc = ~BMC;  //complement 
assign bmg = ~BMG;  //complement 
assign tcm = ~TCM;  //complement 
assign CME =  AMA & BMB & BMC & BMD  |  AMB & BMC & BMD  |  AMC & BMD  |  AMD  ; 
assign cme = ~CME;  //complement 
assign AEA = ~aea;  //complement 
assign bea = ~BEA;  //complement 
assign XBE = ~xbe;  //complement 
assign xad = ~XAD;  //complement 
assign AEB = ~aeb;  //complement 
assign oba = ~OBA;  //complement 
assign obb = ~OBB;  //complement 
assign XBD = ~xbd;  //complement 
assign JAC =  RBA & rbb & rbe  |  rba & RBB & rbe  |  rba & rbb & RBE  |  RBA & RBB & RBE  ; 
assign jac = ~JAC; //complement 
assign jbc =  RBA & rbb & rbe  |  rba & RBB & rbe  |  rba & rbb & RBE  |  rba & rbb & rbe  ; 
assign JBC = ~jbc;  //complement 
assign AEC = ~aec;  //complement 
assign xae = ~XAE;  //complement 
assign SXB = ~sxb;  //complement 
assign SXC = ~sxc;  //complement 
assign SXD = ~sxd;  //complement 
assign rba = ~RBA;  //complement 
assign RFA = ~rfa;  //complement 
assign AED = ~aed;  //complement 
assign bed = ~BED;  //complement 
assign obc = ~OBC;  //complement 
assign obd = ~OBD;  //complement 
assign UAA =  SAA & sab & sac  |  saa & SAB & sac  |  saa & sab & SAC  |  SAA & SAB & SAC  ; 
assign uaa = ~UAA; //complement 
assign uba =  SAA & sab & sac  |  saa & SAB & sac  |  saa & sab & SAC  |  saa & sab & sac  ; 
assign UBA = ~uba;  //complement 
assign sab = ~SAB;  //complement 
assign SBB = ~sbb;  //complement 
assign vaa = ~VAA;  //complement 
assign AMA = ~ama;  //complement 
assign bma = ~BMA;  //complement 
assign UBC =  SBB & sbe & sbh  |  sbb & SBE & sbh  |  sbb & sbe & SBH  |  SBB & SBE & SBH  ; 
assign ubc = ~UBC; //complement 
assign ucb =  SBB & sbe & sbh  |  sbb & SBE & sbh  |  sbb & sbe & SBH  |  sbb & sbe & sbh  ; 
assign UCB = ~ucb;  //complement 
assign AMB = ~amb;  //complement 
assign oda = ~ODA;  //complement 
assign odb = ~ODB;  //complement 
assign vbb = ~VBB;  //complement 
assign VCB = ~vcb;  //complement 
assign JAG =  RDA & rdb & rde  |  rda & RDB & rde  |  rda & rdb & RDE  |  RDA & RDB & RDE  ; 
assign jag = ~JAG; //complement 
assign jbg =  RDA & rdb & rde  |  rda & RDB & rde  |  rda & rdb & RDE  |  rda & rdb & rde  ; 
assign JBG = ~jbg;  //complement 
assign AMC = ~amc;  //complement 
assign SZB = ~szb;  //complement 
assign SZC = ~szc;  //complement 
assign SZD = ~szd;  //complement 
assign rda = ~RDA;  //complement 
assign RHA = ~rha;  //complement 
assign AMD = ~amd;  //complement 
assign bmd = ~BMD;  //complement 
assign odc = ~ODC;  //complement 
assign odd = ~ODD;  //complement 
assign sbh = ~SBH;  //complement 
assign SCE = ~sce;  //complement 
assign XPC = ~xpc;  //complement 
assign GFA = ~gfa;  //complement 
assign HFA = ~hfa;  //complement 
assign XPD = ~xpd;  //complement 
assign XPE = ~xpe;  //complement 
assign GFB = ~gfb;  //complement 
assign HFB = ~hfb;  //complement 
assign dfb =  bfa  ; 
assign DFB = ~dfb;  //complement 
assign dfc =  afb & bfa  |  bfb  ; 
assign DFC = ~dfc;  //complement 
assign VPB = ~vpb;  //complement 
assign GFC = ~gfc;  //complement 
assign HFC = ~hfc;  //complement 
assign dfd =  bfa & afb & afc  |  bfb & afc  |  bfc  ; 
assign DFD = ~dfd; //complement 
assign VRB = ~vrb;  //complement 
assign XVC = ~xvc;  //complement 
assign GFD = ~gfd;  //complement 
assign HFD = ~hfd;  //complement 
assign VQB = ~vqb;  //complement 
assign GNA = ~gna;  //complement 
assign HNA = ~hna;  //complement 
assign XVD = ~xvd;  //complement 
assign XVE = ~xve;  //complement 
assign XVF = ~xvf;  //complement 
assign GNB = ~gnb;  //complement 
assign HNB = ~hnb;  //complement 
assign dnb =  bna  ; 
assign DNB = ~dnb;  //complement 
assign dnc =  anb & bna  |  bnb  ; 
assign DNC = ~dnc;  //complement 
assign VVB = ~vvb;  //complement 
assign GNC = ~gnc;  //complement 
assign HNC = ~hnc;  //complement 
assign dnd =  bna & anb & anc  |  bnb & anc  |  bnc  ; 
assign DND = ~dnd; //complement 
assign VXB = ~vxb;  //complement 
assign VWB = ~vwb;  //complement 
assign GND = ~gnd;  //complement 
assign HND = ~hnd;  //complement 
assign tcf = ~TCF;  //complement 
assign tdf = ~TDF;  //complement 
assign taf = ~TAF;  //complement 
assign TBF = ~tbf;  //complement 
assign MBA = ~mba;  //complement 
assign EFA = TCF & ~AFA & ~BFA  |  ZZO & ~AFA & BFA  |  tcf & AFA & ~BFA  |  TCF & AFA & BFA; 
assign efa = ~EFA;  //complement 
assign EFB = TCF & ~AFB & ~BFB  |         ZZO & ~AFB & BFB  |  tcf & AFB & ~BFB  |  TCF & AFB & BFB ; 
assign efb = ~EFB;  //complement 
assign CFB =  AFA  ; 
assign cfb = ~CFB;  //complement 
assign CFC =  BFB & AFA  |  AFB  ; 
assign cfc = ~CFC;  //complement 
assign bfb = ~BFB;  //complement 
assign bff = ~BFF;  //complement 
assign EFC = TCF & ~AFC & ~BFC  |  ZZO & ~AFC & BFC  |  tcf & AFC & ~BFC  |  TCF & AFC & BFC; 
assign efc = ~EFC;  //complement 
assign EFD = TCF & ~AFD & ~BFD  |         ZZO & ~AFD & BFD  |  tcf & AFD & ~BFD  |  TCF & AFD & BFD ; 
assign efd = ~EFD;  //complement 
assign CFD =  AFA & BFB & BFC  |  AFB & BFC  |  AFC  ; 
assign cfd = ~CFD; //complement 
assign bfc = ~BFC;  //complement 
assign bfg = ~BFG;  //complement 
assign NBA = ~nba;  //complement 
assign FAF =  BFA & BFF & BFG & BFD  ; 
assign faf = ~FAF;  //complement  
assign FBF =  BFA & BFF & BFG & BFD  ; 
assign fbf = ~FBF;  //complement 
assign CFE =  AFA & BFB & BFC & BFD  |  AFB & BFC & BFD  |  AFC & BFD  |  AFD  ; 
assign cfe = ~CFE;  //complement 
assign PBB =  KAB & NBA  |  MBA  ; 
assign pbb = ~PBB; //complement 
assign NDA = ~nda;  //complement 
assign FAN =  BNA & BNF & BNG & BND  ; 
assign fan = ~FAN;  //complement  
assign FBN =  BNA & BNF & BNG & BND  ; 
assign fbn = ~FBN;  //complement 
assign kcd = ~KCD;  //complement 
assign PDB =  KAD & LBD & LCD & NDA  |  KBD & LCD & NDA  |  KCD & NDA  |  MDA  ; 
assign pdb = ~PDB;  //complement 
assign ENA = TCN & ~ANA & ~BNA  |  ZZO & ~ANA & BNA  |  tcn & ANA & ~BNA  |  TCN & ANA & BNA; 
assign ena = ~ENA;  //complement 
assign ENB = TCN & ~ANB & ~BNB  |         ZZO & ~ANB & BNB  |  tcn & ANB & ~BNB  |  TCN & ANB & BNB ; 
assign enb = ~ENB;  //complement 
assign CNB =  ANA  ; 
assign cnb = ~CNB;  //complement 
assign CNC =  BNB & ANA  |  ANB  ; 
assign cnc = ~CNC;  //complement 
assign bnb = ~BNB;  //complement 
assign bnf = ~BNF;  //complement 
assign ENC = TCN & ~ANC & ~BNC  |  ZZO & ~ANC & BNC  |  tcn & ANC & ~BNC  |  TCN & ANC & BNC; 
assign enc = ~ENC;  //complement 
assign ENDD = TCN & ~ANDD  & ~BND  |         ZZO & ~ANDD  & BND  |  tcn & ANDD  & ~BND  |  TCN & ANDD  & BND ; 
assign endd = ~ENDD;  //complement 
assign CND =  ANA & BNB & BNC  |  ANB & BNC  |  ANC  ; 
assign cnd = ~CND; //complement 
assign bnc = ~BNC;  //complement 
assign bng = ~BNG;  //complement 
assign tcn = ~TCN;  //complement 
assign CNE =  ANA & BNB & BNC & BND  |  ANB & BNC & BND  |  ANC & BND  |  ANDD   ; 
assign cne = ~CNE;  //complement 
assign MDA = ~mda;  //complement 
assign AFA = ~afa;  //complement 
assign bfa = ~BFA;  //complement 
assign SXA = ~sxa;  //complement 
assign SXE = ~sxe;  //complement 
assign SXI = ~sxi;  //complement 
assign rbe = ~RBE;  //complement 
assign RFE = ~rfe;  //complement 
assign AFB = ~afb;  //complement 
assign obe = ~OBE;  //complement 
assign obf = ~OBF;  //complement 
assign AFC = ~afc;  //complement 
assign SXF = ~sxf;  //complement 
assign SXG = ~sxg;  //complement 
assign SXH = ~sxh;  //complement 
assign rbb = ~RBB;  //complement 
assign RFB = ~rfb;  //complement 
assign AFD = ~afd;  //complement 
assign bfd = ~BFD;  //complement 
assign obg = ~OBG;  //complement 
assign obh = ~OBH;  //complement 
assign WDB =  VDA & vdb & vdc  |  vda & VDB & vdc  |  vda & vdb & VDC  |  VDA & VDB & VDC  ; 
assign wdb = ~WDB; //complement 
assign wea =  VDA & vdb & vdc  |  vda & VDB & vdc  |  vda & vdb & VDC  |  vda & vdb & vdc  ; 
assign WEA = ~wea;  //complement 
assign ANA = ~ana;  //complement 
assign bna = ~BNA;  //complement 
assign SZA = ~sza;  //complement 
assign SZE = ~sze;  //complement 
assign SZI = ~szi;  //complement 
assign rde = ~RDE;  //complement 
assign RHE = ~rhe;  //complement 
assign ANB = ~anb;  //complement 
assign ode = ~ODE;  //complement 
assign odf = ~ODF;  //complement 
assign ANC = ~anc;  //complement 
assign SZF = ~szf;  //complement 
assign SZG = ~szg;  //complement 
assign SZH = ~szh;  //complement 
assign rdb = ~RDB;  //complement 
assign RHB = ~rhb;  //complement 
assign ANDD  = ~andd ;  //complement 
assign bnd = ~BND;  //complement 
assign odg = ~ODG;  //complement 
assign odh = ~ODH;  //complement 
assign GGA = ~gga;  //complement 
assign HGA = ~hga;  //complement 
assign xpa = ~XPA;  //complement 
assign xpb = ~XPB;  //complement 
assign GGB = ~ggb;  //complement 
assign HGB = ~hgb;  //complement 
assign dgb =  bga  ; 
assign DGB = ~dgb;  //complement 
assign dgc =  agb & bga  |  bgb  ; 
assign DGC = ~dgc;  //complement 
assign VPC = ~vpc;  //complement 
assign WPA =  VPB & VPC & VPD  ; 
assign wpa = ~WPA;  //complement 
assign WPB =  vpb & VPC & VPD  ; 
assign wpb = ~WPB;  //complement 
assign WPC =  vpc & VPD & VPD  ; 
assign wpc = ~WPC;  //complement 
assign GGC = ~ggc;  //complement 
assign HGC = ~hgc;  //complement 
assign dgd =  bga & agb & agc  |  bgb & agc  |  bgc  ; 
assign DGD = ~dgd; //complement 
assign VRC = ~vrc;  //complement 
assign GGD = ~ggd;  //complement 
assign HGD = ~hgd;  //complement 
assign VQC = ~vqc;  //complement 
assign GOA = ~goa;  //complement 
assign HOA = ~hoa;  //complement 
assign xva = ~XVA;  //complement 
assign xvb = ~XVB;  //complement 
assign GOB = ~gob;  //complement 
assign HOB = ~hob;  //complement 
assign dob =  boa  ; 
assign DOB = ~dob;  //complement 
assign doc =  aob & boa  |  bob  ; 
assign DOC = ~doc;  //complement 
assign VVC = ~vvc;  //complement 
assign WVA =  VVB & VVC & VVD  ; 
assign wva = ~WVA;  //complement 
assign WVB =  vvb & VVC & VVD  ; 
assign wvb = ~WVB;  //complement 
assign WVC =  vvc & VVD & VVD  ; 
assign wvc = ~WVC;  //complement 
assign GOC = ~goc;  //complement 
assign HOC = ~hoc;  //complement 
assign dod =  boa & aob & aoc  |  bob & aoc  |  boc  ; 
assign DOD = ~dod; //complement 
assign VXC = ~vxc;  //complement 
assign VWC = ~vwc;  //complement 
assign GOD = ~god;  //complement 
assign HOD = ~hod;  //complement 
assign tcg = ~TCG;  //complement 
assign tdg = ~TDG;  //complement 
assign tag = ~TAG;  //complement 
assign TBG = ~tbg;  //complement 
assign MBB = ~mbb;  //complement 
assign EGA = TCG & ~AGA & ~BGA  |  ZZO & ~AGA & BGA  |  tcg & AGA & ~BGA  |  TCG & AGA & BGA; 
assign ega = ~EGA;  //complement 
assign EGB = TCG & ~AGB & ~BGB  |         ZZO & ~AGB & BGB  |  tcg & AGB & ~BGB  |  TCG & AGB & BGB ; 
assign egb = ~EGB;  //complement 
assign CGB =  AGA  ; 
assign cgb = ~CGB;  //complement 
assign CGC =  BGB & AGA  |  AGB  ; 
assign cgc = ~CGC;  //complement 
assign bgb = ~BGB;  //complement 
assign bgf = ~BGF;  //complement 
assign EGC = TCG & ~AGC & ~BGC  |  ZZO & ~AGC & BGC  |  tcg & AGC & ~BGC  |  TCG & AGC & BGC; 
assign egc = ~EGC;  //complement 
assign EGD = TCG & ~AGD & ~BGD  |         ZZO & ~AGD & BGD  |  tcg & AGD & ~BGD  |  TCG & AGD & BGD ; 
assign egd = ~EGD;  //complement 
assign CGD =  AGA & BGB & BGC  |  AGB & BGC  |  AGC  ; 
assign cgd = ~CGD; //complement 
assign bgc = ~BGC;  //complement 
assign bgg = ~BGG;  //complement 
assign NBB = ~nbb;  //complement 
assign FAG =  BGA & BGF & BGG & BGD  ; 
assign fag = ~FAG;  //complement  
assign FBG =  BGA & BGF & BGG & BGD  ; 
assign fbg = ~FBG;  //complement 
assign CGE =  AGA & BGB & BGC & BGD  |  AGB & BGC & BGD  |  AGC & BGD  |  AGD  ; 
assign cge = ~CGE;  //complement 
assign PBC =  KAB & NBB  |  MBB  ; 
assign pbc = ~PBC; //complement 
assign NDB = ~ndb;  //complement 
assign FAO =  BOA & BOF & BOG & BOD  ; 
assign fao = ~FAO;  //complement  
assign FBO =  BOA & BOF & BOG & BOD  ; 
assign fbo = ~FBO;  //complement 
assign LCD = ~lcd;  //complement 
assign PDC =  KAD & LBD & LCD & NDB  |  KBD & LCD & NDB  |  KCD & NDB  |  MDB  ; 
assign pdc = ~PDC;  //complement 
assign EOA = TCO & ~AOA & ~BOA  |  ZZO & ~AOA & BOA  |  tco & AOA & ~BOA  |  TCO & AOA & BOA; 
assign eoa = ~EOA;  //complement 
assign EOB = TCO & ~AOB & ~BOB  |         ZZO & ~AOB & BOB  |  tco & AOB & ~BOB  |  TCO & AOB & BOB ; 
assign eob = ~EOB;  //complement 
assign COB =  AOA  ; 
assign cob = ~COB;  //complement 
assign COC =  BOB & AOA  |  AOB  ; 
assign coc = ~COC;  //complement 
assign bob = ~BOB;  //complement 
assign bof = ~BOF;  //complement 
assign EOC = TCO & ~AOC & ~BOC  |  ZZO & ~AOC & BOC  |  tco & AOC & ~BOC  |  TCO & AOC & BOC; 
assign eoc = ~EOC;  //complement 
assign EOD = TCO & ~AOD & ~BOD  |         ZZO & ~AOD & BOD  |  tco & AOD & ~BOD  |  TCO & AOD & BOD ; 
assign eod = ~EOD;  //complement 
assign COD =  AOA & BOB & BOC  |  AOB & BOC  |  AOC  ; 
assign cod = ~COD; //complement 
assign boc = ~BOC;  //complement 
assign bog = ~BOG;  //complement 
assign tco = ~TCO;  //complement 
assign COE =  AOA & BOB & BOC & BOD  |  AOB & BOC & BOD  |  AOC & BOD  |  AOD  ; 
assign coe = ~COE;  //complement 
assign MDB = ~mdb;  //complement 
assign AGA = ~aga;  //complement 
assign bga = ~BGA;  //complement 
assign AGB = ~agb;  //complement 
assign obi = ~OBI;  //complement 
assign obj = ~OBJ;  //complement 
assign sbf = ~SBF;  //complement 
assign SCC = ~scc;  //complement 
assign JAD =  RBC & rbd & rbf  |  rbc & RBD & rbf  |  rbc & rbd & RBF  |  RBC & RBD & RBF  ; 
assign jad = ~JAD; //complement 
assign jbd =  RBC & rbd & rbf  |  rbc & RBD & rbf  |  rbc & rbd & RBF  |  rbc & rbd & rbf  ; 
assign JBD = ~jbd;  //complement 
assign AGC = ~agc;  //complement 
assign SXJ = ~sxj;  //complement 
assign SXK = ~sxk;  //complement 
assign SXL = ~sxl;  //complement 
assign rbc = ~RBC;  //complement 
assign RFC = ~rfc;  //complement 
assign AGD = ~agd;  //complement 
assign bgd = ~BGD;  //complement 
assign obk = ~OBK;  //complement 
assign obl = ~OBL;  //complement 
assign vcd = ~VCD;  //complement 
assign VDB = ~vdb;  //complement 
assign sac = ~SAC;  //complement 
assign SBC = ~sbc;  //complement 
assign AOA = ~aoa;  //complement 
assign boa = ~BOA;  //complement 
assign UCE =  SCC & scf & sch  |  scc & SCF & sch  |  scc & scf & SCH  |  SCC & SCF & SCH  ; 
assign uce = ~UCE; //complement 
assign udb =  SCC & scf & sch  |  scc & SCF & sch  |  scc & scf & SCH  |  scc & scf & sch  ; 
assign UDB = ~udb;  //complement 
assign QAA = ~qaa;  //complement 
assign qab = ~QAB;  //complement 
assign qac = ~QAC;  //complement 
assign qad = ~QAD;  //complement 
assign AOB = ~aob;  //complement 
assign odi = ~ODI;  //complement 
assign odj = ~ODJ;  //complement 
assign UBD =  SBC & sbf & sbi  |  sbc & SBF & sbi  |  sbc & sbf & SBI  |  SBC & SBF & SBI  ; 
assign ubd = ~UBD; //complement 
assign ucc =  SBC & sbf & sbi  |  sbc & SBF & sbi  |  sbc & sbf & SBI  |  sbc & sbf & sbi  ; 
assign UCC = ~ucc;  //complement 
assign JAH =  RDC & rdd & rdf  |  rdc & RDD & rdf  |  rdc & rdd & RDF  |  RDC & RDD & RDF  ; 
assign jah = ~JAH; //complement 
assign jbh =  RDC & rdd & rdf  |  rdc & RDD & rdf  |  rdc & rdd & RDF  |  rdc & rdd & rdf  ; 
assign JBH = ~jbh;  //complement 
assign AOC = ~aoc;  //complement 
assign SZJ = ~szj;  //complement 
assign SZK = ~szk;  //complement 
assign SZL = ~szl;  //complement 
assign rdc = ~RDC;  //complement 
assign RHC = ~rhc;  //complement 
assign AOD = ~aod;  //complement 
assign bod = ~BOD;  //complement 
assign odk = ~ODK;  //complement 
assign odl = ~ODL;  //complement 
assign sbi = ~SBI;  //complement 
assign SCF = ~scf;  //complement 
assign GHA = ~gha;  //complement 
assign HHA = ~hha;  //complement 
assign GHB = ~ghb;  //complement 
assign HHB = ~hhb;  //complement 
assign dhb =  bha  ; 
assign DHB = ~dhb;  //complement 
assign dhc =  ahb & bha  |  bhb  ; 
assign DHC = ~dhc;  //complement 
assign VPD = ~vpd;  //complement 
assign GHC = ~ghc;  //complement 
assign HHC = ~hhc;  //complement 
assign dhd =  bha & ahb & ahc  |  bhb & ahc  |  bhc  ; 
assign DHD = ~dhd; //complement 
assign VRD = ~vrd;  //complement 
assign GHD = ~ghd;  //complement 
assign HHD = ~hhd;  //complement 
assign VQD = ~vqd;  //complement 
assign qdd = ~QDD;  //complement 
assign qed = ~QED;  //complement 
assign tfa = ~TFA;  //complement 
assign tfb = ~TFB;  //complement 
assign GPA = ~gpa;  //complement 
assign HPA = ~hpa;  //complement 
assign GPB = ~gpb;  //complement 
assign HPB = ~hpb;  //complement 
assign dpb =  bpa  ; 
assign DPB = ~dpb;  //complement 
assign dpc =  apb & bpa  |  bpb  ; 
assign DPC = ~dpc;  //complement 
assign VVD = ~vvd;  //complement 
assign GPC = ~gpc;  //complement 
assign HPC = ~hpc;  //complement 
assign dpd =  bpa & apb & apc  |  bpb & apc  |  bpc  ; 
assign DPD = ~dpd; //complement 
assign VXD = ~vxd;  //complement 
assign VWD = ~vwd;  //complement 
assign GPD = ~gpd;  //complement 
assign HPD = ~hpd;  //complement 
assign qea = ~QEA;  //complement 
assign qef = ~QEF;  //complement 
assign tch = ~TCH;  //complement 
assign tdh = ~TDH;  //complement 
assign qdb = ~QDB;  //complement 
assign tah = ~TAH;  //complement 
assign TBH = ~tbh;  //complement 
assign MBC = ~mbc;  //complement 
assign EHA = TCH & ~AHA & ~BHA  |  ZZO & ~AHA & BHA  |  tch & AHA & ~BHA  |  TCH & AHA & BHA; 
assign eha = ~EHA;  //complement 
assign EHB = TCH & ~AHB & ~BHB  |         ZZO & ~AHB & BHB  |  tch & AHB & ~BHB  |  TCH & AHB & BHB ; 
assign ehb = ~EHB;  //complement 
assign CHB =  AHA  ; 
assign chb = ~CHB;  //complement 
assign CHC =  BHB & AHA  |  AHB  ; 
assign chc = ~CHC;  //complement 
assign bhb = ~BHB;  //complement 
assign bhf = ~BHF;  //complement 
assign EHC = TCH & ~AHC & ~BHC  |  ZZO & ~AHC & BHC  |  tch & AHC & ~BHC  |  TCH & AHC & BHC; 
assign ehc = ~EHC;  //complement 
assign EHD = TCH & ~AHD & ~BHD  |         ZZO & ~AHD & BHD  |  tch & AHD & ~BHD  |  TCH & AHD & BHD ; 
assign ehd = ~EHD;  //complement 
assign CHD =  AHA & BHB & BHC  |  AHB & BHC  |  AHC  ; 
assign chd = ~CHD; //complement 
assign bhc = ~BHC;  //complement 
assign bhg = ~BHG;  //complement 
assign NBC = ~nbc;  //complement 
assign FAH =  BHA & BHF & BHG & BHD  ; 
assign fah = ~FAH;  //complement  
assign CHE =  AHA & BHB & BHC & BHD  |  AHB & BHC & BHD  |  AHC & BHD  |  AHD  ; 
assign che = ~CHE;  //complement 
assign PBD =  KAB & NBC  |  MBC  ; 
assign pbd = ~PBD; //complement 
assign NDC = ~ndc;  //complement 
assign LBC = ~lbc;  //complement 
assign LBD = ~lbd;  //complement 
assign PDD =  KAD & LBD & LCD & NDC  |  KBD & LCD & NDC  |  KCD & NDC  |  MDC  ; 
assign pdd = ~PDD;  //complement 
assign EPA = TCP & ~APA & ~BPA  |  ZZO & ~APA & BPA  |  tcp & APA & ~BPA  |  TCP & APA & BPA; 
assign epa = ~EPA;  //complement 
assign EPB = TCP & ~APB & ~BPB  |         ZZO & ~APB & BPB  |  tcp & APB & ~BPB  |  TCP & APB & BPB ; 
assign epb = ~EPB;  //complement 
assign CPB =  APA  ; 
assign cpb = ~CPB;  //complement 
assign CPC =  BPB & APA  |  APB  ; 
assign cpc = ~CPC;  //complement 
assign EPC = TCP & ~APC & ~BPC  |  ZZO & ~APC & BPC  |  tcp & APC & ~BPC  |  TCP & APC & BPC; 
assign epc = ~EPC;  //complement 
assign EPD = TCP & ~APD & ~BPD  |         ZZO & ~APD & BPD  |  tcp & APD & ~BPD  |  TCP & APD & BPD ; 
assign epd = ~EPD;  //complement 
assign CPD =  APA & BPB & BPC  |  APB & BPC  |  APC  ; 
assign cpd = ~CPD; //complement 
assign QEG = ~qeg;  //complement 
assign tcp = ~TCP;  //complement 
assign MDC = ~mdc;  //complement 
assign AHA = ~aha;  //complement 
assign bha = ~BHA;  //complement 
assign qca = ~QCA;  //complement 
assign qda = ~QDA;  //complement 
assign RBF = ~rbf;  //complement 
assign SXM = ~sxm;  //complement 
assign tea = ~TEA;  //complement 
assign teb = ~TEB;  //complement 
assign AHB = ~ahb;  //complement 
assign obm = ~OBM;  //complement 
assign obn = ~OBN;  //complement 
assign qec = ~QEC;  //complement 
assign qee = ~QEE;  //complement 
assign qfc = ~QFC;  //complement 
assign qfe = ~QFE;  //complement 
assign QBD = ~qbd;  //complement 
assign AHC = ~ahc;  //complement 
assign QBB = ~qbb;  //complement 
assign SXN = ~sxn;  //complement 
assign SXO = ~sxo;  //complement 
assign SXP = ~sxp;  //complement 
assign rbd = ~RBD;  //complement 
assign RFD = ~rfd;  //complement 
assign sch = ~SCH;  //complement 
assign AHD = ~ahd;  //complement 
assign bhd = ~BHD;  //complement 
assign obo = ~OBO;  //complement 
assign obp = ~OBP;  //complement 
assign QCD = ~qcd;  //complement 
assign qdc = ~QDC;  //complement 
assign qde = ~QDE;  //complement 
assign QDF = ~qdf;  //complement 
assign JBJ =  RFB & rfc & rfd  |  rfb & RFC & rfd  |  rfb & rfc & RFD  |  RFB & RFC & RFD  ; 
assign jbj = ~JBJ; //complement 
assign jcb =  RFB & rfc & rfd  |  rfb & RFC & rfd  |  rfb & rfc & RFD  |  rfb & rfc & rfd  ; 
assign JCB = ~jcb;  //complement 
assign APA = ~apa;  //complement 
assign bpa = ~BPA;  //complement 
assign QCE = ~qce;  //complement 
assign QBE = ~qbe;  //complement 
assign QCB = ~qcb;  //complement 
assign RDF = ~rdf;  //complement 
assign SZM = ~szm;  //complement 
assign QBA = ~qba;  //complement 
assign APB = ~apb;  //complement 
assign bpb = ~BPB;  //complement 
assign odm = ~ODM;  //complement 
assign odn = ~ODN;  //complement 
assign QCC = ~qcc;  //complement 
assign QBC = ~qbc;  //complement 
assign APC = ~apc;  //complement 
assign bpc = ~BPC;  //complement 
assign tec = ~TEC;  //complement 
assign SZN = ~szn;  //complement 
assign SZO = ~szo;  //complement 
assign SZP = ~szp;  //complement 
assign rdd = ~RDD;  //complement 
assign RHD = ~rhd;  //complement 
assign APD = ~apd;  //complement 
assign bpd = ~BPD;  //complement 
assign odo = ~ODO;  //complement 
assign odp = ~ODP;  //complement 
assign JBL =  RHB & rhc & rhd  |  rhb & RHC & rhd  |  rhb & rhc & RHD  |  RHB & RHC & RHD  ; 
assign jbl = ~JBL; //complement 
assign jcd =  RHB & rhc & rhd  |  rhb & RHC & rhd  |  rhb & rhc & RHD  |  rhb & rhc & rhd  ; 
assign JCD = ~jcd;  //complement 
assign iaa = ~IAA; //complement 
assign iab = ~IAB; //complement 
assign iac = ~IAC; //complement 
assign iad = ~IAD; //complement 
assign iae = ~IAE; //complement 
assign iaf = ~IAF; //complement 
assign iag = ~IAG; //complement 
assign iah = ~IAH; //complement 
assign iai = ~IAI; //complement 
assign iaj = ~IAJ; //complement 
assign iak = ~IAK; //complement 
assign ial = ~IAL; //complement 
assign iam = ~IAM; //complement 
assign ian = ~IAN; //complement 
assign iao = ~IAO; //complement 
assign iap = ~IAP; //complement 
assign iba = ~IBA; //complement 
assign ibb = ~IBB; //complement 
assign ibc = ~IBC; //complement 
assign ibd = ~IBD; //complement 
assign ibe = ~IBE; //complement 
assign ibf = ~IBF; //complement 
assign ibg = ~IBG; //complement 
assign ibh = ~IBH; //complement 
assign ibi = ~IBI; //complement 
assign ibj = ~IBJ; //complement 
assign ibk = ~IBK; //complement 
assign ibl = ~IBL; //complement 
assign ibm = ~IBM; //complement 
assign ibn = ~IBN; //complement 
assign ibo = ~IBO; //complement 
assign ibp = ~IBP; //complement 
assign ica = ~ICA; //complement 
assign icb = ~ICB; //complement 
assign icc = ~ICC; //complement 
assign icd = ~ICD; //complement 
assign ice = ~ICE; //complement 
assign icf = ~ICF; //complement 
assign icg = ~ICG; //complement 
assign ich = ~ICH; //complement 
assign ici = ~ICI; //complement 
assign icj = ~ICJ; //complement 
assign ick = ~ICK; //complement 
assign icl = ~ICL; //complement 
assign icm = ~ICM; //complement 
assign icn = ~ICN; //complement 
assign ico = ~ICO; //complement 
assign icp = ~ICP; //complement 
assign ida = ~IDA; //complement 
assign idb = ~IDB; //complement 
assign idc = ~IDC; //complement 
assign idd = ~IDD; //complement 
assign ide = ~IDE; //complement 
assign idf = ~IDF; //complement 
assign idg = ~IDG; //complement 
assign idh = ~IDH; //complement 
assign idi = ~IDI; //complement 
assign idj = ~IDJ; //complement 
assign idk = ~IDK; //complement 
assign idl = ~IDL; //complement 
assign idm = ~IDM; //complement 
assign idn = ~IDN; //complement 
assign ido = ~IDO; //complement 
assign idp = ~IDP; //complement 
assign iga = ~IGA; //complement 
assign ipb = ~IPB; //complement 
assign ipc = ~IPC; //complement 
assign ipd = ~IPD; //complement 
always@(posedge IZZ )
   begin 
 RMA <=  XMA & YMA  |  XPA & YMB  |  XSA & YMC  |  XVA & YMD  ; 
 gaa <=  eaa  |  tda  ; 
 RMB <=  XMB & YMA  |  XPB & YMB  |  XSB & YMC  |  XVB & YMD  ; 
 gab <=  cab & eab  |  CAB & EAB  |  tda  ; 
 vma <=  SWA  |  SWB  |  SWC  |  SWD  ; 
 RMC <=  XMC & YMA  |  XPC & YMB  |  XSC & YMC  |  XVC & YMD  ; 
 gac <=  cac & eac  |  CAC & EAC  |  tda  ; 
 vna <=  SWB & swc  |  SWD  ; 
 voa <=  SWD  |  SWC  ; 
 RMD <=  XMD & YMA  |  XPD & YMB  |  XSD & YMC  |  XVD & YMD  ; 
 gad <=  cad & ead  |  CAD & EAD  |  tda  ; 
 gia <=  eia  |  tda  ; 
 hia <=  EIA  |  tda  ; 
 gib <=  cib & eib  |  CIB & EIB  |  tda  ; 
 hib <=  dib & eib  |  DIB & EIB  |  tda  ; 
 vsa <=  SYA  |  SYB  |  SYC  |  SYD  ; 
 gic <=  cic & eic  |  CIC & EIC  |  tda  ; 
 hic <=  dic & eic  |  DIC & EIC  |  tda  ; 
 vua <=  SYD  |  SYC  ; 
 vta <=  SYB & syc  |  SYD  ; 
 gid <=  cid & eid  |  CID & EID  |  tda  ; 
 hid <=  did & eid  |  DID & EID  |  tda  ; 
 TCA <= QEF ; 
 TDA <= QEA ; 
 TAA <= QDB ; 
 tba <= qdb ; 
 KAB <=  CAE & FAB & FAC & FAD  |  CBE & FAC & FAD  |  CCE & FAD  |  CDE  ; 
 BIB <=  SYB & tba  |  ICB  |  syb & TBA  ; 
 BIF <=  SYB & tba  |  ICB  |  syb & TBA  ; 
 BIC <=  SYC & tba  |  ICC  |  syc & TBA  ; 
 BIG <=  SYC & tba  |  ICC  |  syc & TBA  ; 
 TCI <= QEG ; 
 aaa <=  swa & taa  |  iaa  |  SWA & TAA  ; 
 BAA <=  SWA & taa  |  IAA  |  swa & TAA  ; 
 aab <=  swb & taa  |  iab  |  SWB & TAA  ; 
 BAB <=  SWB & taa  |  IAB  |  swb & TAA  ; 
 OAA <=  GAA  |  XBA  |  RMA  ; 
 aac <=  swc & taa  |  iac  |  SWC & TAA  ; 
 BAC <=  SWC & taa  |  IAC  |  swc & TAA  ; 
 OAC <=  GAC  |  XBC & yac  |  xbc & YAC  |  RMC  ; 
 swb <= iab ; 
 swc <= iac ; 
 swd <= iad ; 
 RAA <=  IAD & iab & iac  |  iad & IAB & iac  |  iad & iab & IAC  |  IAD & IAB & IAC  ;
 rea <=  IAD & iab & iac  |  iad & IAB & iac  |  iad & iab & IAC  |  iad & iab & iac  ;
 aad <=  swd & taa  |  iad  |  SWD & TAA  ; 
 BAD <=  SWD & taa  |  IAD  |  swd & TAA  ; 
 OAD <=  GAD  |  XBD & yad  |  xbd & YAD  |  RMD  ; 
 SAA <=  JAA & jab & jae  |  jaa & JAB & jae  |  jaa & jab & JAE  |  JAA & JAB & JAE  ;
 sba <=  JAA & jab & jae  |  jaa & JAB & jae  |  jaa & jab & JAE  |  jaa & jab & jae  ;
 aia <=  sya & taa  |  ica  |  SYA & TAA  ; 
 BIA <=  SYA & taa  |  ICA  |  sya & TAA  ; 
 aib <=  syb & taa  |  icb  |  SYB & TAA  ; 
 OCA <=  GIA & pca  |  HIA & PCA  ; 
 OCB <=  GIB & pca  |  HIB & PCA  ; 
 aic <=  syc & taa  |  icc  |  SYC & TAA  ; 
 syb <= icb ; 
 syc <= icc ; 
 syd <= icd ; 
 RCA <=  ICD & icb & icc  |  icd & ICB & icc  |  icd & icb & ICC  |  ICD & ICB & ICC  ;
 rga <=  ICD & icb & icc  |  icd & ICB & icc  |  icd & icb & ICC  |  icd & icb & icc  ;
 aid <=  syd & taa  |  icd  |  SYD & TAA  ; 
 BID <=  SYD & taa  |  ICD  |  syd & TAA  ; 
 OCC <=  GIC & pca  |  HIC & PCA  ; 
 OCD <=  GID & pca  |  HID & PCA  ; 
 OAB <=  GAB  |  XBB  |  RMB  ; 
 xmc <=  wmc & vmb  |  wmc & vmd  ; 
 rme <=  ymc & yma  ; 
 rmf <=  ymb & yma  ; 
 gba <=  eba  |  tdb  ; 
 hba <=  EBA  |  tdb  ; 
 xmd <=  vmd  |  vmc  ; 
 xme <=  wma  |  vma  ; 
 gbb <=  cbb & ebb  |  CBB & EBB  |  tdb  ; 
 hbb <=  dbb & ebb  |  DBB & EBB  |  tdb  ; 
 vmb <=  SWE  |  SWF  |  SWG  |  SWH  ; 
 RMG <= YME ; 
 gbc <=  cbc & ebc  |  CBC & EBC  |  tdb  ; 
 hbc <=  dbc & ebc  |  DBC & EBC  |  tdb  ; 
 vob <=  SWH  |  SWG  ; 
 gbd <=  cbd & ebd  |  CBD & EBD  |  tdb  ; 
 hbd <=  dbd & ebd  |  DBD & EBD  |  tdb  ; 
 vnb <=  SWF & swg  |  SWH  ; 
 xsc <=  wsc & vsb  |  wsc & vsd  ; 
 gja <=  eja  |  tdb  ; 
 hja <=  EJA  |  tdb  ; 
 xsd <=  vsd  |  vsc  ; 
 xsf <=  wsa  |  vsa  ; 
 xse <=  wsa  |  vsa  ; 
 gjb <=  cjb & ejb  |  CJB & EJB  |  tdb  ; 
 hjb <=  djb & ejb  |  DJB & EJB  |  tdb  ; 
 vsb <=  SYE  |  SYF  |  SYG  |  SYH  ; 
 vtb <=  SYF & syg  |  SYH  ; 
 gjc <=  cjc & ejc  |  CJC & EJC  |  tdb  ; 
 hjc <=  djc & ejc  |  DJC & EJC  |  tdb  ; 
 vub <=  SYH  |  SYG  ; 
 gjd <=  cjd & ejd  |  CJD & EJD  |  tdb  ; 
 hjd <=  djd & ejd  |  DJD & EJD  |  tdb  ; 
 TCB <= QEF ; 
 TDB <= QEA ; 
 TAB <= QDB ; 
 tbb <= qdb ; 
 maa <=  cae  ; 
 BBB <=  SWF & tbb  |  IAF  |  swf & TBB  ; 
 BBF <=  SWF & tbb  |  IAF  |  swf & TBB  ; 
 BBC <=  SWG & tbb  |  IAG  |  swg & TBB  ; 
 BBG <=  SWG & tbb  |  IAG  |  swg & TBB  ; 
 nca <=  fai  ; 
 KAC <=  CAE & FAB & FAC & FAD  |  CBE & FAC & FAD  |  CCE & FAD  |  CDE  ; 
 BJB <=  SYF & tbb  |  ICF  |  syf & TBB  ; 
 BJF <=  SYF & tbb  |  ICF  |  syf & TBB  ; 
 BJC <=  SYG & tbb  |  ICG  |  syg & TBB  ; 
 BJG <=  SYG & tbb  |  ICG  |  syg & TBB  ; 
 TCJ <= QEG ; 
 mca <=  cie  ; 
 aba <=  swe & tab  |  iae  |  SWE & TAB  ; 
 BBA <=  SWE & tab  |  IAE  |  swe & TAB  ; 
 OAE <=  GBA & pab  |  HBA & PAB  |  XBE & yae  |  xbe & YAE  |  RME  ; 
 swa <= iaa ; 
 swe <= iae ; 
 swi <= iai ; 
 RAE <=  IAA & iae & iai  |  iaa & IAE & iai  |  iaa & iae & IAI  |  IAA & IAE & IAI  ;
 ree <=  IAA & iae & iai  |  iaa & IAE & iai  |  iaa & iae & IAI  |  iaa & iae & iai  ;
 abb <=  swf & tab  |  iaf  |  SWF & TAB  ; 
 OAF <=  GBB & pab  |  HBB & PAB  |  XBF & yaf  |  xbf & YAF  |  RMF  ; 
 SBD <=  JBA & rea & ree  |  jba & REA & ree  |  jba & rea & REE  |  JBA & REA & REE  ;
 sca <=  JBA & rea & ree  |  jba & REA & ree  |  jba & rea & REE  |  jba & rea & ree  ;
 abc <=  swg & tab  |  iag  |  SWG & TAB  ; 
 OAG <=  GBC & pab  |  HBC & PAB  |  XBF & YAF  |  RMG  ; 
 swf <= iaf ; 
 swg <= iag ; 
 swh <= iah ; 
 RAB <=  IAH & iaf & iag  |  iah & IAF & iag  |  iah & iaf & IAG  |  IAH & IAF & IAG  ;
 reb <=  IAH & iaf & iag  |  iah & IAF & iag  |  iah & iaf & IAG  |  iah & iaf & iag  ;
 abd <=  swh & tab  |  iah  |  SWH & TAB  ; 
 BBD <=  SWH & tab  |  IAH  |  swh & TAB  ; 
 OAH <=  GBD & pab  |  HBD & PAB  ; 
 aja <=  sye & tab  |  ice  |  SYE & TAB  ; 
 BJA <=  SYE & tab  |  ICE  |  sye & TAB  ; 
 sya <= ica ; 
 sye <= ice ; 
 syi <= ici ; 
 RCE <=  ICA & ice & ici  |  ica & ICE & ici  |  ica & ice & ICI  |  ICA & ICE & ICI  ;
 rge <=  ICA & ice & ici  |  ica & ICE & ici  |  ica & ice & ICI  |  ica & ice & ici  ;
 ajb <=  syf & tab  |  icf  |  SYF & TAB  ; 
 OCE <=  GJA & pcb  |  HJA & PCB  ; 
 OCF <=  GJB & pcb  |  HJB & PCB  ; 
 VCC <=  UCA & ucd & ucf  |  uca & UCD & ucf  |  uca & ucd & UCF  |  UCA & UCD & UCF  ;
 vda <=  UCA & ucd & ucf  |  uca & UCD & ucf  |  uca & ucd & UCF  |  uca & ucd & ucf  ;
 SBG <=  JBE & rga & rge  |  jbe & RGA & rge  |  jbe & rga & RGE  |  JBE & RGA & RGE  ;
 scd <=  JBE & rga & rge  |  jbe & RGA & rge  |  jbe & rga & RGE  |  jbe & rga & rge  ;
 ajc <=  syg & tab  |  icg  |  SYG & TAB  ; 
 syf <= icf ; 
 syg <= icg ; 
 syh <= ich ; 
 RCB <=  ICH & icf & icg  |  ich & ICF & icg  |  ich & icf & ICG  |  ICH & ICF & ICG  ;
 rgb <=  ICH & icf & icg  |  ich & ICF & icg  |  ich & icf & ICG  |  ich & icf & icg  ;
 ajd <=  syh & tab  |  ich  |  SYH & TAB  ; 
 BJD <=  SYH & tab  |  ICH  |  syh & TAB  ; 
 OCG <=  GJC & pcb  |  HJC & PCB  ; 
 OCH <=  GJD & pcb  |  HJD & PCB  ; 
 gca <=  eca  |  tdc  ; 
 hca <=  ECA  |  tdc  ; 
 XMA <=  WMA & VNA  |  WMB & VNB  |  WMC & VNC  |  vmd & VND  ; 
 XMB <=  WMA & VOA  |  WMB & VOB  |  WMC & VOC  |  vmd & VOD  ; 
 gcb <=  ccb & ecb  |  CCB & ECB  |  tdc  ; 
 hcb <=  dcb & ecb  |  DCB & ECB  |  tdc  ; 
 vmc <=  SWI  |  SWJ  |  SWK  |  SWL  ; 
 gcc <=  ccc & ecc  |  CCC & ECC  |  tdc  ; 
 hcc <=  dcc & ecc  |  DCC & ECC  |  tdc  ; 
 voc <=  SWL  |  SWK  ; 
 gcd <=  ccd & ecd  |  CCD & ECD  |  tdc  ; 
 hcd <=  dcd & ecd  |  DCD & ECD  |  tdc  ; 
 vnc <=  SWJ & swk  |  SWL  ; 
 gka <=  eka  |  tdc  ; 
 hka <=  EKA  |  tdc  ; 
 XSA <=  WSA & VTA  |  WSB & VTB  |  WSC & VTC  |  vsd & VTD  ; 
 XSB <=  WSA & VUA  |  WSB & VUB  |  WSC & VUC  |  vsd & VUD  ; 
 gkb <=  ckb & ekb  |  CKB & EKB  |  tdc  ; 
 hkb <=  dkb & ekb  |  DKB & EKB  |  tdc  ; 
 vsc <=  SYI  |  SYJ  |  SYK  |  SYL  ; 
 gkc <=  ckc & ekc  |  CKC & EKC  |  tdc  ; 
 hkc <=  dkc & ekc  |  DKC & EKC  |  tdc  ; 
 vuc <=  SYL  |  SYK  ; 
 vtc <=  SYJ & syk  |  SYL  ; 
 gkd <=  ckd & ekd  |  CKD & EKD  |  tdc  ; 
 hkd <=  dkd & ekd  |  DKD & EKD  |  tdc  ; 
 TCC <= QEF ; 
 TDC <= QEA ; 
 TAC <= QDB ; 
 tbc <= qdb ; 
 mab <=  cae & cbe & cbe  |  fab & cbe  ; 
 BCB <=  SWJ & tbc  |  IAJ  |  swj & TBC  ; 
 BCF <=  SWJ & tbc  |  IAJ  |  swj & TBC  ; 
 BCC <=  SWK & tbc  |  IAK  |  swk & TBC  ; 
 BCG <=  SWK & tbc  |  IAK  |  swk & TBC  ; 
 ncb <=  fai  |  faj  ; 
 KAD <=  CAE & FAB & FAC & FAD  |  CBE & FAC & FAD  |  CCE & FAD  |  CDE  ; 
 BKB <=  SYJ & tbc  |  ICJ  |  syj & TBC  ; 
 BKF <=  SYJ & tbc  |  ICJ  |  syj & TBC  ; 
 BKC <=  SYK & tbc  |  ICK  |  syk & TBC  ; 
 BKG <=  SYK & tbc  |  ICK  |  syk & TBC  ; 
 TCK <= QEG ; 
 mcb <=  cie & cje & cje  |  fbj & cje  ; 
 aca <=  swi & tac  |  iai  |  SWI & TAC  ; 
 BCA <=  SWI & tac  |  IAI  |  swi & TAC  ; 
 acb <=  swj & tac  |  iaj  |  SWJ & TAC  ; 
 OAI <=  GCA & pac  |  HCA & PAC  ; 
 OAJ <=  GCB & pac  |  HCB & PAC  ; 
 acc <=  swk & tac  |  iak  |  SWK & TAC  ; 
 swj <= iaj ; 
 swk <= iak ; 
 swl <= ial ; 
 RAC <=  IAL & iaj & iak  |  ial & IAJ & iak  |  ial & iaj & IAK  |  IAL & IAJ & IAK  ;
 rec <=  IAL & iaj & iak  |  ial & IAJ & iak  |  ial & iaj & IAK  |  ial & iaj & iak  ;
 SBJ <= JBB ; 
 acd <=  swl & tac  |  ial  |  SWL & TAC  ; 
 BCD <=  SWL & tac  |  IAL  |  swl & TAC  ; 
 OAK <=  GCC & pac  |  HCC & PAC  ; 
 OAL <=  GCD & pac  |  HCD & PAC  ; 
 aka <=  syi & tac  |  ici  |  SYI & TAC  ; 
 BKA <=  SYI & tac  |  ICI  |  syi & TAC  ; 
 VBA <=  UBB & sbj & sbk  |  ubb & SBJ & sbk  |  ubb & sbj & SBK  |  UBB & SBJ & SBK  ;
 vca <=  UBB & sbj & sbk  |  ubb & SBJ & sbk  |  ubb & sbj & SBK  |  ubb & sbj & sbk  ;
 akb <=  syj & tac  |  icj  |  SYJ & TAC  ; 
 OCI <=  GKA & pcc  |  HKA & PCC  ; 
 OCJ <=  GKB & pcc  |  HKB & PCC  ; 
 VDC <=  UDA & udb & udc  |  uda & UDB & udc  |  uda & udb & UDC  |  UDA & UDB & UDC  ;
 vea <=  UDA & udb & udc  |  uda & UDB & udc  |  uda & udb & UDC  |  uda & udb & udc  ;
 VEB <= UEA ; 
 akc <=  syk & tac  |  ick  |  SYK & TAC  ; 
 syj <= icj ; 
 syk <= ick ; 
 syl <= icl ; 
 RCC <=  ICL & icj & ick  |  icl & ICJ & ick  |  icl & icj & ICK  |  ICL & ICJ & ICK  ;
 rgc <=  ICL & icj & ick  |  icl & ICJ & ick  |  icl & icj & ICK  |  icl & icj & ick  ;
 SBK <= JBF ; 
 akd <=  syl & tac  |  icl  |  SYL & TAC  ; 
 BKD <=  SYL & tac  |  ICL  |  syl & TAC  ; 
 OCK <=  GKC & pcc  |  HKC & PCC  ; 
 OCL <=  GKD & pcc  |  HKD & PCC  ; 
 gda <=  eda  |  tdd  ; 
 hda <=  EDA  |  tdd  ; 
 gdb <=  cdb & edb  |  CDB & EDB  |  tdd  ; 
 hdb <=  ddb & edb  |  DDB & EDB  |  tdd  ; 
 vmd <=  SWM  |  SWN  |  SWO  |  SWP  ; 
 gdc <=  cdc & edc  |  CDC & EDC  |  tdd  ; 
 hdc <=  ddc & edc  |  DDC & EDC  |  tdd  ; 
 vod <=  SWP  |  SWO  ; 
 gdd <=  cdd & edd  |  CDD & EDD  |  tdd  ; 
 hdd <=  ddd & edd  |  DDD & EDD  |  tdd  ; 
 vnd <=  SWN & swo  |  SWP  ; 
 gla <=  ela  |  tdd  ; 
 hla <=  ELA  |  tdd  ; 
 glb <=  clb & elb  |  CLB & ELB  |  tdd  ; 
 hlb <=  dlb & elb  |  DLB & ELB  |  tdd  ; 
 vsd <=  SYM  |  SYN  |  SYO  |  SYP  ; 
 glc <=  clc & elc  |  CLC & ELC  |  tdd  ; 
 hlc <=  dlc & elc  |  DLC & ELC  |  tdd  ; 
 vud <=  SYP  |  SYO  ; 
 vtd <=  SYN & syo  |  SYP  ; 
 gld <=  cld & eld  |  CLD & ELD  |  tdd  ; 
 hld <=  dld & eld  |  DLD & ELD  |  tdd  ; 
 TCD <= QEF ; 
 TDD <= QEA ; 
 TAD <= QDB ; 
 tbd <= qdb ; 
 mac <=  ZZI & cae & cbe & cce  |  ZZI & cae & cbe & cce  |  fab & cbe & cce  |  ZZI & fac & cce  ; 
 BDB <=  SWN & tbd  |  IAN  |  swn & TBD  ; 
 BDF <=  SWN & tbd  |  IAN  |  swn & TBD  ; 
 BDC <=  SWO & tbd  |  IAO  |  swo & TBD  ; 
 BDG <=  SWO & tbd  |  IAO  |  swo & TBD  ; 
 ncc <=  fai  |  faj  |  fak  ; 
 KBC <=  CEE & FAF & FAG & FAH  |  CFE & FAG & FAH  |  CGE & FAH  |  CHE  ; 
 BLB <=  SYN & tbd  |  ICN  |  syn & TBD  ; 
 BLF <=  SYN & tbd  |  ICN  |  syn & TBD  ; 
 BLC <=  SYO & tbd  |  ICO  |  syo & TBD  ; 
 BLG <=  SYO & tbd  |  ICO  |  syo & TBD  ; 
 TCL <= QEG ; 
 mcc <=  ZZI & cie & cje & cke  |  ZZI & cie & cje & cke  |  fbj & cje & cke  |  ZZI & fbk & cke  ; 
 ada <=  swm & tad  |  iam  |  SWM & TAD  ; 
 BDA <=  SWM & tad  |  IAM  |  swm & TAD  ; 
 xbf <=  wfa  |  tea  ; 
 xbb <=  tea  |  VBB & VBA  |  vba & vbb  ; 
 raf <= iam ; 
 swm <= iam ; 
 adb <=  swn & tad  |  ian  |  SWN & TAD  ; 
 OAM <=  GDA & pad  |  HDA & PAD  ; 
 OAN <=  GDB & pad  |  HDB & PAD  ; 
 xbc <=  tea  |  WCA & VCD  |  vcd & wca  ; 
 SBE <=  JBC & jbi & rfa  |  jbc & JBI & rfa  |  jbc & jbi & RFA  |  JBC & JBI & RFA  ;
 scb <=  JBC & jbi & rfa  |  jbc & JBI & rfa  |  jbc & jbi & RFA  |  jbc & jbi & rfa  ;
 adc <=  swo & tad  |  iao  |  SWO & TAD  ; 
 XAB <= VBA & VBB ; 
 swn <= ian ; 
 swo <= iao ; 
 swp <= iap ; 
 RAD <=  IAP & ian & iao  |  iap & IAN & iao  |  iap & ian & IAO  |  IAP & IAN & IAO  ;
 red <=  IAP & ian & iao  |  iap & IAN & iao  |  iap & ian & IAO  |  iap & ian & iao  ;
 add <=  swp & tad  |  iap  |  SWP & TAD  ; 
 BDD <=  SWP & tad  |  IAP  |  swp & TAD  ; 
 OAO <=  GDC & pad  |  HDC & PAD  ; 
 OAP <=  GDD & pad  |  HDD & PAD  ; 
 ala <=  sym & tad  |  icm  |  SYM & TAD  ; 
 BLA <=  SYM & tad  |  ICM  |  sym & TAD  ; 
 XAC <= VCD & WCA ; 
 rcf <= icm ; 
 sym <= icm ; 
 xba <=  vaa  |  tec  ; 
 alb <=  syn & tad  |  icn  |  SYN & TAD  ; 
 OCM <=  GLA & pcd  |  HLA & PCD  ; 
 OCN <=  GLB & pcd  |  HLB & PCD  ; 
 SCG <=  JCA & jcc & jcd  |  jca & JCC & jcd  |  jca & jcc & JCD  |  JCA & JCC & JCD  ;
 sda <=  JCA & jcc & jcd  |  jca & JCC & jcd  |  jca & jcc & JCD  |  jca & jcc & jcd  ;
 alc <=  syo & tad  |  ico  |  SYO & TAD  ; 
 syn <= icn ; 
 syo <= ico ; 
 syp <= icp ; 
 RCD <=  ICP & icn & ico  |  icp & ICN & ico  |  icp & icn & ICO  |  ICP & ICN & ICO  ;
 rgd <=  ICP & icn & ico  |  icp & ICN & ico  |  icp & icn & ICO  |  icp & icn & ico  ;
 ald <=  syp & tad  |  icp  |  SYP & TAD  ; 
 BLD <=  SYP & tad  |  ICP  |  syp & TAD  ; 
 OCO <=  GLC & pcd  |  HLC & PCD  ; 
 OCP <=  GLD & pcd  |  HLD & PCD  ; 
 gea <=  eea  |  tde  ; 
 hea <=  EEA  |  tde  ; 
 geb <=  ceb & eeb  |  CEB & EEB  |  tde  ; 
 heb <=  deb & eeb  |  DEB & EEB  |  tde  ; 
 vpa <=  SXA  |  SXB  |  SXC  |  SXD  ; 
 gec <=  cec & eec  |  CEC & EEC  |  tde  ; 
 hec <=  dec & eec  |  DEC & EEC  |  tde  ; 
 vra <=  SXD  |  SXC  ; 
 ged <=  ced & eed  |  CED & EED  |  tde  ; 
 hed <=  ded & eed  |  DED & EED  |  tde  ; 
 vqa <=  SXB & sxc  |  SXD  ; 
 gma <=  ema  |  tde  ; 
 hma <=  EMA  |  tde  ; 
 gmb <=  cmb & emb  |  CMB & EMB  |  tde  ; 
 hmb <=  dmb & emb  |  DMB & EMB  |  tde  ; 
 vva <=  SZA  |  SZB  |  SZC  |  SZD  ; 
 gmc <=  cmc & emc  |  CMC & EMC  |  tde  ; 
 hmc <=  dmc & emc  |  DMC & EMC  |  tde  ; 
 vxa <=  SZD  |  SZC  ; 
 vwa <=  SZB & szc  |  SZD  ; 
 gmd <=  cmd & emd  |  CMD & EMD  |  tde  ; 
 hmd <=  dmd & emd  |  DMD & EMD  |  tde  ; 
 TCE <= QEF ; 
 TDE <= QEA ; 
 TAE <= QDB ; 
 tbe <= qdb ; 
 BEB <=  SXB & tbe  |  IBB  |  sxb & TBE  ; 
 BEF <=  SXB & tbe  |  IBB  |  sxb & TBE  ; 
 BEC <=  SXC & tbe  |  IBC  |  sxc & TBE  ; 
 BEG <=  SXC & tbe  |  IBC  |  sxc & TBE  ; 
 KBD <=  CEE & FAF & FAG & FAH  |  CFE & FAG & FAH  |  CGE & FAH  |  CHE  ; 
 BMB <=  SZB & tbe  |  IDB  |  szb & TBE  ; 
 BMF <=  SZB & tbe  |  IDB  |  szb & TBE  ; 
 BMC <=  SZC & tbe  |  IDC  |  szc & TBE  ; 
 BMG <=  SZC & tbe  |  IDC  |  szc & TBE  ; 
 TCM <= QEG ; 
 aea <=  sxa & tae  |  iba  |  SXA & TAE  ; 
 BEA <=  SXA & tae  |  IBA  |  sxa & TAE  ; 
 xbe <=  tea  |  WEB & WEA  |  wea & web  ; 
 XAD <= WDA & WDB ; 
 aeb <=  sxb & tae  |  ibb  |  SXB & TAE  ; 
 OBA <=  GEA & pba  |  HEA & PBA  ; 
 OBB <=  GEB & pba  |  HEB & PBA  ; 
 xbd <=  tea  |  WDB & WDA  |  wda & wdb  ; 
 aec <=  sxc & tae  |  ibc  |  SXC & TAE  ; 
 XAE <= WEA & WEB ; 
 sxb <= ibb ; 
 sxc <= ibc ; 
 sxd <= ibd ; 
 RBA <=  IBD & ibb & ibc  |  ibd & IBB & ibc  |  ibd & ibb & IBC  |  IBD & IBB & IBC  ;
 rfa <=  IBD & ibb & ibc  |  ibd & IBB & ibc  |  ibd & ibb & IBC  |  ibd & ibb & ibc  ;
 aed <=  sxd & tae  |  ibd  |  SXD & TAE  ; 
 BED <=  SXD & tae  |  IBD  |  sxd & TAE  ; 
 OBC <=  GEC & pba  |  HEC & PBA  ; 
 OBD <=  GED & pba  |  HED & PBA  ; 
 SAB <=  JAC & jaf & jag  |  jac & JAF & jag  |  jac & jaf & JAG  |  JAC & JAF & JAG  ;
 sbb <=  JAC & jaf & jag  |  jac & JAF & jag  |  jac & jaf & JAG  |  jac & jaf & jag  ;
 VAA <= UAA ; 
 ama <=  sza & tae  |  ida  |  SZA & TAE  ; 
 BMA <=  SZA & tae  |  IDA  |  sza & TAE  ; 
 amb <=  szb & tae  |  idb  |  SZB & TAE  ; 
 ODA <=  GMA & pda  |  HMA & PDA  ; 
 ODB <=  GMB & pda  |  HMB & PDA  ; 
 VBB <=  UBA & ubc & ubd  |  uba & UBC & ubd  |  uba & ubc & UBD  |  UBA & UBC & UBD  ;
 vcb <=  UBA & ubc & ubd  |  uba & UBC & ubd  |  uba & ubc & UBD  |  uba & ubc & ubd  ;
 amc <=  szc & tae  |  idc  |  SZC & TAE  ; 
 szb <= idb ; 
 szc <= idc ; 
 szd <= idd ; 
 RDA <=  IDD & idb & idc  |  idd & IDB & idc  |  idd & idb & IDC  |  IDD & IDB & IDC  ;
 rha <=  IDD & idb & idc  |  idd & IDB & idc  |  idd & idb & IDC  |  idd & idb & idc  ;
 amd <=  szd & tae  |  idd  |  SZD & TAE  ; 
 BMD <=  SZD & tae  |  IDD  |  szd & TAE  ; 
 ODC <=  GMC & pda  |  HMC & PDA  ; 
 ODD <=  GMD & pda  |  HMD & PDA  ; 
 SBH <=  JBG & jbk & rha  |  jbg & JBK & rha  |  jbg & jbk & RHA  |  JBG & JBK & RHA  ;
 sce <=  JBG & jbk & rha  |  jbg & JBK & rha  |  jbg & jbk & RHA  |  jbg & jbk & rha  ;
 xpc <=  wpc & vpb  |  wpc & vpd  ; 
 gfa <=  efa  |  tdf  ; 
 hfa <=  EFA  |  tdf  ; 
 xpd <=  vpd  |  vpc  ; 
 xpe <=  wpa  |  vpa  ; 
 gfb <=  cfb & efb  |  CFB & EFB  |  tdf  ; 
 hfb <=  dfb & efb  |  DFB & EFB  |  tdf  ; 
 vpb <=  SXE  |  SXF  |  SXG  |  SXH  ; 
 gfc <=  cfc & efc  |  CFC & EFC  |  tdf  ; 
 hfc <=  dfc & efc  |  DFC & EFC  |  tdf  ; 
 vrb <=  SXH  |  SXG  ; 
 xvc <=  wvc & vvb  |  wvc & vvd  ; 
 gfd <=  cfd & efd  |  CFD & EFD  |  tdf  ; 
 hfd <=  dfd & efd  |  DFD & EFD  |  tdf  ; 
 vqb <=  SXF & sxg  |  SXH  ; 
 gna <=  ena  |  tdf  ; 
 hna <=  ENA  |  tdf  ; 
 xvd <=  vvd  |  vvc  ; 
 xve <=  wva  |  vva  |  tfa  ; 
 xvf <=  wva  |  vva  |  tfa  ; 
 gnb <=  cnb & enb  |  CNB & ENB  |  tdf  ; 
 hnb <=  dnb & enb  |  DNB & ENB  |  tdf  ; 
 vvb <=  SZE  |  SZF  |  SZG  |  SZH  ; 
 gnc <=  cnc & enc  |  CNC & ENC  |  tdf  ; 
 hnc <=  dnc & enc  |  DNC & ENC  |  tdf  ; 
 vxb <=  SZH  |  SZG  ; 
 vwb <=  SZF & szg  |  SZH  ; 
 gnd <=  cnd & endd |  CND & ENDD  |  tdf  ; 
 hnd <=  dnd & endd |  DND & ENDD  |  tdf  ; 
 TCF <= QEF ; 
 TDF <= QEA ; 
 TAF <= QDB ; 
 tbf <= qdb ; 
 mba <=  cee  ; 
 BFB <=  SXF & tbf  |  IBF  |  sxf & TBF  ; 
 BFF <=  SXF & tbf  |  IBF  |  sxf & TBF  ; 
 BFC <=  SXG & tbf  |  IBG  |  sxg & TBF  ; 
 BFG <=  SXG & tbf  |  IBG  |  sxg & TBF  ; 
 nba <=  fae  ; 
 nda <=  fam  ; 
 KCD <=  CIE & FAJ & FAK & FAL  |  CJE & FAK & FAL  |  CKE & FAL  |  CLE  ; 
 BNB <=  SZF & tbf  |  IDF  |  szf & TBF  ; 
 BNF <=  SZF & tbf  |  IDF  |  szf & TBF  ; 
 BNC <=  SZG & tbf  |  IDG  |  szg & TBF  ; 
 BNG <=  SZG & tbf  |  IDG  |  szg & TBF  ; 
 TCN <= QEG ; 
 mda <=  cme  ; 
 afa <=  sxe & taf  |  ibe  |  SXE & TAF  ; 
 BFA <=  SXE & taf  |  IBE  |  sxe & TAF  ; 
 sxa <= iba ; 
 sxe <= ibe ; 
 sxi <= ibi ; 
 RBE <=  IBA & ibe & ibi  |  iba & IBE & ibi  |  iba & ibe & IBI  |  IBA & IBE & IBI  ;
 rfe <=  IBA & ibe & ibi  |  iba & IBE & ibi  |  iba & ibe & IBI  |  iba & ibe & ibi  ;
 afb <=  sxf & taf  |  ibf  |  SXF & TAF  ; 
 OBE <=  GFA & pbb  |  HFA & PBB  ; 
 OBF <=  GFB & pbb  |  HFB & PBB  ; 
 afc <=  sxg & taf  |  ibg  |  SXG & TAF  ; 
 sxf <= ibf ; 
 sxg <= ibg ; 
 sxh <= ibh ; 
 RBB <=  IBH & ibf & ibg  |  ibh & IBF & ibg  |  ibh & ibf & IBG  |  IBH & IBF & IBG  ;
 rfb <=  IBH & ibf & ibg  |  ibh & IBF & ibg  |  ibh & ibf & IBG  |  ibh & ibf & ibg  ;
 afd <=  sxh & taf  |  ibh  |  SXH & TAF  ; 
 BFD <=  SXH & taf  |  IBH  |  sxh & TAF  ; 
 OBG <=  GFC & pbb  |  HFC & PBB  ; 
 OBH <=  GFD & pbb  |  HFD & PBB  ; 
 ana <=  sze & taf  |  ide  |  SZE & TAF  ; 
 BNA <=  SZE & taf  |  IDE  |  sze & TAF  ; 
 sza <= ida ; 
 sze <= ide ; 
 szi <= idi ; 
 RDE <=  IDA & ide & idi  |  ida & IDE & idi  |  ida & ide & IDI  |  IDA & IDE & IDI  ;
 rhe <=  IDA & ide & idi  |  ida & IDE & idi  |  ida & ide & IDI  |  ida & ide & idi  ;
 anb <=  szf & taf  |  idf  |  SZF & TAF  ; 
 ODE <=  GNA & pdb  |  HNA & PDB  ; 
 ODF <=  GNB & pdb  |  HNB & PDB  ; 
 anc <=  szg & taf  |  idg  |  SZG & TAF  ; 
 szf <= idf ; 
 szg <= idg ; 
 szh <= idh ; 
 RDB <=  IDH & idf & idg  |  idh & IDF & idg  |  idh & idf & IDG  |  IDH & IDF & IDG  ;
 rhb <=  IDH & idf & idg  |  idh & IDF & idg  |  idh & idf & IDG  |  idh & idf & idg  ;
 andd  <=  szh & taf  |  idh  |  SZH & TAF  ; 
 BND <=  SZH & taf  |  IDH  |  szh & TAF  ; 
 ODG <=  GNC & pdb  |  HNC & PDB  ; 
 ODH <=  GND & pdb  |  HND & PDB  ; 
 gga <=  ega  |  tdg  ; 
 hga <=  EGA  |  tdg  ; 
 XPA <=  WPA & VQA  |  WPB & VQB  |  WPC & VQC  |  vpd & VQD  ; 
 XPB <=  WPA & VRA  |  WPB & VRB  |  WPC & VRC  |  vpd & VRD  ; 
 ggb <=  cgb & egb  |  CGB & EGB  |  tdg  ; 
 hgb <=  dgb & egb  |  DGB & EGB  |  tdg  ; 
 vpc <=  SXI  |  SXJ  |  SXK  |  SXL  ; 
 ggc <=  cgc & egc  |  CGC & EGC  |  tdg  ; 
 hgc <=  dgc & egc  |  DGC & EGC  |  tdg  ; 
 vrc <=  SXL  |  SXK  ; 
 ggd <=  cgd & egd  |  CGD & EGD  |  tdg  ; 
 hgd <=  dgd & egd  |  DGD & EGD  |  tdg  ; 
 vqc <=  SXJ & sxk  |  SXL  ; 
 goa <=  eoa  |  tdg  ; 
 hoa <=  EOA  |  tdg  ; 
 XVA <=  WVA & VWA  |  WVB & VWB  |  WVC & VWC  |  vvd & VWD  ; 
 XVB <=  WVA & VXA  |  WVB & VXB  |  WVC & VXC  |  vvd & VXD  ; 
 gob <=  cob & eob  |  COB & EOB  |  tdg  ; 
 hob <=  dob & eob  |  DOB & EOB  |  tdg  ; 
 vvc <=  SZI  |  SZJ  |  SZK  |  SZL  ; 
 goc <=  coc & eoc  |  COC & EOC  |  tdg  ; 
 hoc <=  doc & eoc  |  DOC & EOC  |  tdg  ; 
 vxc <=  SZL  |  SZK  ; 
 vwc <=  SZJ & szk  |  SZL  ; 
 god <=  cod & eod  |  COD & EOD  |  tdg  ; 
 hod <=  dod & eod  |  DOD & EOD  |  tdg  ; 
 TCG <= QEF ; 
 TDG <= QEA ; 
 TAG <= QDB ; 
 tbg <= qdb ; 
 mbb <=  cee & cfe & cfe  |  fbf & cfe  ; 
 BGB <=  SXJ & tbg  |  IBJ  |  sxj & TBG  ; 
 BGF <=  SXJ & tbg  |  IBJ  |  sxj & TBG  ; 
 BGC <=  SXK & tbg  |  IBK  |  sxk & TBG  ; 
 BGG <=  SXK & tbg  |  IBK  |  sxk & TBG  ; 
 nbb <=  fae  |  faf  ; 
 ndb <=  fam  |  fan  ; 
 lcd <=  fai  |  faj  |  fak  |  fal  ; 
 BOB <=  SZJ & tbg  |  IDJ  |  szj & TBG  ; 
 BOF <=  SZJ & tbg  |  IDJ  |  szj & TBG  ; 
 BOC <=  SZK & tbg  |  IDK  |  szk & TBG  ; 
 BOG <=  SZK & tbg  |  IDK  |  szk & TBG  ; 
 TCO <= QEG ; 
 mdb <=  cme & cne & cne  |  fbn & cne  ; 
 aga <=  sxi & tag  |  ibi  |  SXI & TAG  ; 
 BGA <=  SXI & tag  |  IBI  |  sxi & TAG  ; 
 agb <=  sxj & tag  |  ibj  |  SXJ & TAG  ; 
 OBI <=  GGA & pbc  |  HGA & PBC  ; 
 OBJ <=  GGB & pbc  |  HGB & PBC  ; 
 SBF <=  JBD & jbj & rfe  |  jbd & JBJ & rfe  |  jbd & jbj & RFE  |  JBD & JBJ & RFE  ;
 scc <=  JBD & jbj & rfe  |  jbd & JBJ & rfe  |  jbd & jbj & RFE  |  jbd & jbj & rfe  ;
 agc <=  sxk & tag  |  ibk  |  SXK & TAG  ; 
 sxj <= ibj ; 
 sxk <= ibk ; 
 sxl <= ibl ; 
 RBC <=  IBL & ibj & ibk  |  ibl & IBJ & ibk  |  ibl & ibj & IBK  |  IBL & IBJ & IBK  ;
 rfc <=  IBL & ibj & ibk  |  ibl & IBJ & ibk  |  ibl & ibj & IBK  |  ibl & ibj & ibk  ;
 agd <=  sxl & tag  |  ibl  |  SXL & TAG  ; 
 BGD <=  SXL & tag  |  IBL  |  sxl & TAG  ; 
 OBK <=  GGC & pbc  |  HGC & PBC  ; 
 OBL <=  GGD & pbc  |  HGD & PBC  ; 
 VCD <=  UCB & ucc & uce  |  ucb & UCC & uce  |  ucb & ucc & UCE  |  UCB & UCC & UCE  ;
 vdb <=  UCB & ucc & uce  |  ucb & UCC & uce  |  ucb & ucc & UCE  |  ucb & ucc & uce  ;
 SAC <=  JAD & jah  |  JAH & jad  ; 
 sbc <=  jah & jah  |  jad & jad  ; 
 aoa <=  szi & tag  |  idi  |  SZI & TAG  ; 
 BOA <=  SZI & tag  |  IDI  |  szi & TAG  ; 
 qaa <= iga ; 
 QAB <= IPB ; 
 QAC <= IPC ; 
 QAD <= IPD ; 
 aob <=  szj & tag  |  idj  |  SZJ & TAG  ; 
 ODI <=  GOA & pdc  |  HOA & PDC  ; 
 ODJ <=  GOB & pdc  |  HOB & PDC  ; 
 aoc <=  szk & tag  |  idk  |  SZK & TAG  ; 
 szj <= idj ; 
 szk <= idk ; 
 szl <= idl ; 
 RDC <=  IDL & idj & idk  |  idl & IDJ & idk  |  idl & idj & IDK  |  IDL & IDJ & IDK  ;
 rhc <=  IDL & idj & idk  |  idl & IDJ & idk  |  idl & idj & IDK  |  idl & idj & idk  ;
 aod <=  szl & tag  |  idl  |  SZL & TAG  ; 
 BOD <=  SZL & tag  |  IDL  |  szl & TAG  ; 
 ODK <=  GOC & pdc  |  HOC & PDC  ; 
 ODL <=  GOD & pdc  |  HOD & PDC  ; 
 SBI <=  JBH & jbl & rhe  |  jbh & JBL & rhe  |  jbh & jbl & RHE  |  JBH & JBL & RHE  ;
 scf <=  JBH & jbl & rhe  |  jbh & JBL & rhe  |  jbh & jbl & RHE  |  jbh & jbl & rhe  ;
 gha <=  eha  |  tdh  ; 
 hha <=  EHA  |  tdh  ; 
 ghb <=  chb & ehb  |  CHB & EHB  |  tdh  ; 
 hhb <=  dhb & ehb  |  DHB & EHB  |  tdh  ; 
 vpd <=  SXM  |  SXN  |  SXO  |  SXP  ; 
 ghc <=  chc & ehc  |  CHC & EHC  |  tdh  ; 
 hhc <=  dhc & ehc  |  DHC & EHC  |  tdh  ; 
 vrd <=  SXP  |  SXO  ; 
 ghd <=  chd & ehd  |  CHD & EHD  |  tdh  ; 
 hhd <=  dhd & ehd  |  DHD & EHD  |  tdh  ; 
 vqd <=  SXN & sxo  |  SXP  ; 
 QDD <= QCD ; 
 QED <= QDD ; 
 TFA <= QED ; 
 TFB <= TFA ; 
 gpa <=  epa  |  tdh  ; 
 hpa <=  EPA  |  tdh  ; 
 gpb <=  cpb & epb  |  CPB & EPB  |  tdh  ; 
 hpb <=  dpb & epb  |  DPB & EPB  |  tdh  ; 
 vvd <=  SZM  |  SZN  |  SZO  |  SZP  ; 
 gpc <=  cpc & epc  |  CPC & EPC  |  tdh  ; 
 hpc <=  dpc & epc  |  DPC & EPC  |  tdh  ; 
 vxd <=  SZP  |  SZO  ; 
 vwd <=  SZN & szo  |  SZP  ; 
 gpd <=  cpd & epd  |  CPD & EPD  |  tdh  ; 
 hpd <=  dpd & epd  |  DPD & EPD  |  tdh  ; 
 QEA <= QDA ; 
 QEF <= QDF ; 
 TCH <= QEF ; 
 TDH <= QEA ; 
 QDB <= QCB ; 
 TAH <= QDB ; 
 tbh <= qdb ; 
 mbc <=  ZZI & cee & cfe & cge  |  ZZI & cee & cfe & cge  |  fbf & cfe & cge  |  ZZI & fbg & cge  ; 
 BHB <=  SXN & tbh  |  IBN  |  sxn & TBH  ; 
 BHF <=  SXN & tbh  |  IBN  |  sxn & TBH  ; 
 BHC <=  SXO & tbh  |  IBO  |  sxo & TBH  ; 
 BHG <=  SXO & tbh  |  IBO  |  sxo & TBH  ; 
 nbc <=  fae  |  faf  |  fag  ; 
 ndc <=  fam  |  fan  |  fao  ; 
 lbc <=  fae  |  faf  |  fag  |  fah  ; 
 lbd <=  fae  |  faf  |  fag  |  fah  ; 
 qeg <= qdf ; 
 TCP <= QEG ; 
 mdc <=  ZZI & cme & cne & coe  |  ZZI & cme & cne & coe  |  fbn & cne & coe  |  ZZI & fbo & coe  ; 
 aha <=  sxm & tah  |  ibm  |  SXM & TAH  ; 
 BHA <=  SXM & tah  |  IBM  |  sxm & TAH  ; 
 QCA <=  QBB  |  QBA  ; 
 QDA <= QCA ; 
 rbf <= ibm ; 
 sxm <= ibm ; 
 TEA <= QFC ; 
 TEB <= TEA ; 
 ahb <=  sxn & tah  |  ibn  |  SXN & TAH  ; 
 OBM <=  GHA & pbd  |  HHA & PBD  ; 
 OBN <=  GHB & pbd  |  HHB & PBD  ; 
 QEC <= QDC ; 
 QEE <= QDE ; 
 QFC <= QEC ; 
 QFE <= QEE ; 
 qbd <=  qac  |  qab  |  qaa  ; 
 ahc <=  sxo & tah  |  ibo  |  SXO & TAH  ; 
 qbb <=  QAC  |  qab  |  qaa  ; 
 sxn <= ibn ; 
 sxo <= ibo ; 
 sxp <= ibp ; 
 RBD <=  IBP & ibn & ibo  |  ibp & IBN & ibo  |  ibp & ibn & IBO  |  IBP & IBN & IBO  ;
 rfd <=  IBP & ibn & ibo  |  ibp & IBN & ibo  |  ibp & ibn & IBO  |  ibp & ibn & ibo  ;
 SCH <= JCB ; 
 ahd <=  sxp & tah  |  ibp  |  SXP & TAH  ; 
 BHD <=  SXP & tah  |  IBP  |  sxp & TAH  ; 
 OBO <=  GHC & pbd  |  HHC & PBD  ; 
 OBP <=  GHD & pbd  |  HHD & PBD  ; 
 qcd <= qbd ; 
 QDC <= QCC ; 
 QDE <= QCE ; 
 qdf <= qcb ; 
 apa <=  szm & tah  |  idm  |  SZM & TAH  ; 
 BPA <=  SZM & tah  |  IDM  |  szm & TAH  ; 
 qce <=  qbc  |  qbe  ; 
 qbe <= qad ; 
 qcb <= qbb ; 
 rdf <= idm ; 
 szm <= idm ; 
 qba <=  QAC  |  QAB  |  qaa  ; 
 apb <=  szn & tah  |  idn  |  SZN & TAH  ; 
 BPB <=  SZN & tah  |  IDN  |  szn & TAH  ; 
 ODM <=  GPA & pdd  |  HPA & PDD  ; 
 ODN <=  GPB & pdd  |  HPB & PDD  ; 
 qcc <=  qbc  |  QBE  ; 
 qbc <=  qac  |  QAB  |  qaa  ; 
 apc <=  szo & tah  |  ido  |  SZO & TAH  ; 
 BPC <=  SZO & tah  |  IDO  |  szo & TAH  ; 
 TEC <=  QFE  |  QFC  ; 
 szn <= idn ; 
 szo <= ido ; 
 szp <= idp ; 
 RDD <=  IDP & idn & ido  |  idp & IDN & ido  |  idp & idn & IDO  |  IDP & IDN & IDO  ;
 rhd <=  IDP & idn & ido  |  idp & IDN & ido  |  idp & idn & IDO  |  idp & idn & ido  ;
 apd <=  szp & tah  |  idp  |  SZP & TAH  ; 
 BPD <=  SZP & tah  |  IDP  |  szp & TAH  ; 
 ODO <=  GPC & pdd  |  HPC & PDD  ; 
 ODP <=  GPD & pdd  |  HPD & PDD  ; 
 end 
endmodule;
