module qb( IZZ,
 IAA, 
 IAB, 
 IAC, 
 IAD, 
 IAE, 
 IAF, 
 IAG, 
 IAH, 
 IAI, 
 IAJ, 
 IAK, 
 IAL, 
 IBA, 
 IBB, 
 IBC, 
 IBD, 
 IBE, 
 IBF, 
 IBG, 
 IBH, 
 IBI, 
 IBJ, 
 IBK, 
 IBL, 
 ICA, 
 ICB, 
 ICC, 
 ICD, 
 ICE, 
 ICF, 
 ICG, 
 ICH, 
 ICI, 
 ICJ, 
 ICK, 
 ICL, 
 IDA, 
 IDB, 
 IDC, 
 IDD, 
 IDE, 
 IDF, 
 IDG, 
 IDH, 
 IDI, 
 IDJ, 
 IDK, 
 IDL, 
 IEA, 
 IEB, 
 IEC, 
 IED, 
 IEE, 
 IEF, 
 IEG, 
 IEH, 
 IEI, 
 IEJ, 
 IEK, 
 IEL, 
 IEM, 
 IEN, 
 IEO, 
 IEP, 
 IEQ, 
 IER, 
 IES, 
 IET, 
 IEU, 
 IEV, 
 IEW, 
 IEX, 
 IFA, 
 IFB, 
 IFC, 
 IFD, 
 IFE, 
 IGA, 
 IGB, 
 IGC, 
 IJA, 
 IJB, 
 IJC, 
 IJD, 
 IJE, 
 IJF, 
 IJG, 
 IJH, 
 IJI, 
 IJJ, 
 IJK, 
 IJL, 
 IJM, 
 IJN, 
 IJO, 
 IJP, 
 IKA, 
 IKB, 
 IKC, 
 IKD, 
 IKE, 
 IKF, 
 IKG, 
 IKH, 
 IKI, 
 IKJ, 
 IKK, 
 IKL, 
 IKM, 
 IKN, 
 IKO, 
 IKP, 
 OAA, 
 OAB, 
 OAC, 
 OAD, 
 OAE, 
 OAF, 
 OAG, 
 OAH, 
 OAI, 
 OAJ, 
 OAK, 
 OAL, 
 OAM, 
 OAN, 
 OAO, 
 OAP, 
 OBA, 
 OBB, 
 OBC, 
 OBD, 
 OBE, 
 OBF, 
 OBG, 
 OBH, 
 OBI, 
 OBJ, 
 OBK, 
 OBL, 
 OBM, 
 OBN, 
 OBO, 
 OBP, 
 ODA, 
 ODB, 
 ODC, 
 ODD, 
 ODE, 
 ODF, 
 ODG, 
 ODH, 
 OEA, 
 OEB, 
 OEC, 
 OED, 
 OEE, 
 OEF, 
 OEG, 
 OEH, 
 OFA, 
 OFB, 
 OFC, 
 OFD, 
 OFE, 
 OGA, 
 OGB, 
 OGC, 
 OGD, 
 OGE, 
 OHA, 
 OHB, 
 OHC, 
 OHD, 
 OHE, 
 OIA, 
 OIB, 
 OIC, 
 OID, 
 OIE, 
 OJA, 
 OJB, 
 OJC, 
 OJD, 
 OJE, 
 OJF, 
 OKA, 
 OKB, 
 OKC, 
 OKD, 
 OKE, 
 OKF, 
 OLA, 
 OLB, 
 OLC, 
 OLD, 
 OLE, 
 OLF, 
 OMA, 
 OMB, 
 OMC, 
 OMD, 
 OME, 
 OMF, 
 ONA, 
 ONB, 
 ONC, 
 OND, 
 ONE, 
 ONF, 
 ONG, 
 ONH, 
 ONI, 
 ONJ, 
 ONK, 
 ONL, 
 ONM, 
 ONN, 
 ONO, 
 ONP, 
 OOA, 
 OOB, 
 OOC, 
 OOD, 
 OOE, 
 OOF, 
 OOG, 
 OOH, 
 OOI, 
 OOJ, 
 OOK, 
 OOL, 
 OOM, 
 OON, 
 OOO, 
 OOP, 
 OPA, 
 OPB, 
 OPC, 
 OPD, 
 OPE, 
 OPF, 
 OPG, 
 OPH, 
 OPI, 
 OPJ, 
 OPK, 
 OPL, 
 OPM, 
 OPN, 
 OPO, 
 OPP, 
 OQA, 
 OQB, 
 OQC, 
 OQD, 
 OQE, 
 OQF, 
 OQG, 
 OQH, 
 OQI, 
 OQJ, 
 OQK, 
 OQL, 
 OQM, 
 OQN, 
OQO ); 
    
 input IZZ; 
 input IAA; 
 input IAB; 
 input IAC; 
 input IAD; 
 input IAE; 
 input IAF; 
 input IAG; 
 input IAH; 
 input IAI; 
 input IAJ; 
 input IAK; 
 input IAL; 
 input IBA; 
 input IBB; 
 input IBC; 
 input IBD; 
 input IBE; 
 input IBF; 
 input IBG; 
 input IBH; 
 input IBI; 
 input IBJ; 
 input IBK; 
 input IBL; 
 input ICA; 
 input ICB; 
 input ICC; 
 input ICD; 
 input ICE; 
 input ICF; 
 input ICG; 
 input ICH; 
 input ICI; 
 input ICJ; 
 input ICK; 
 input ICL; 
 input IDA; 
 input IDB; 
 input IDC; 
 input IDD; 
 input IDE; 
 input IDF; 
 input IDG; 
 input IDH; 
 input IDI; 
 input IDJ; 
 input IDK; 
 input IDL; 
 input IEA; 
 input IEB; 
 input IEC; 
 input IED; 
 input IEE; 
 input IEF; 
 input IEG; 
 input IEH; 
 input IEI; 
 input IEJ; 
 input IEK; 
 input IEL; 
 input IEM; 
 input IEN; 
 input IEO; 
 input IEP; 
 input IEQ; 
 input IER; 
 input IES; 
 input IET; 
 input IEU; 
 input IEV; 
 input IEW; 
 input IEX; 
 input IFA; 
 input IFB; 
 input IFC; 
 input IFD; 
 input IFE; 
 input IGA; 
 input IGB; 
 input IGC; 
 input IJA; 
 input IJB; 
 input IJC; 
 input IJD; 
 input IJE; 
 input IJF; 
 input IJG; 
 input IJH; 
 input IJI; 
 input IJJ; 
 input IJK; 
 input IJL; 
 input IJM; 
 input IJN; 
 input IJO; 
 input IJP; 
 input IKA; 
 input IKB; 
 input IKC; 
 input IKD; 
 input IKE; 
 input IKF; 
 input IKG; 
 input IKH; 
 input IKI; 
 input IKJ; 
 input IKK; 
 input IKL; 
 input IKM; 
 input IKN; 
 input IKO; 
 input IKP; 
 output OAA; 
 output OAB; 
 output OAC; 
 output OAD; 
 output OAE; 
 output OAF; 
 output OAG; 
 output OAH; 
 output OAI; 
 output OAJ; 
 output OAK; 
 output OAL; 
 output OAM; 
 output OAN; 
 output OAO; 
 output OAP; 
 output OBA; 
 output OBB; 
 output OBC; 
 output OBD; 
 output OBE; 
 output OBF; 
 output OBG; 
 output OBH; 
 output OBI; 
 output OBJ; 
 output OBK; 
 output OBL; 
 output OBM; 
 output OBN; 
 output OBO; 
 output OBP; 
 output ODA; 
 output ODB; 
 output ODC; 
 output ODD; 
 output ODE; 
 output ODF; 
 output ODG; 
 output ODH; 
 output OEA; 
 output OEB; 
 output OEC; 
 output OED; 
 output OEE; 
 output OEF; 
 output OEG; 
 output OEH; 
 output OFA; 
 output OFB; 
 output OFC; 
 output OFD; 
 output OFE; 
 output OGA; 
 output OGB; 
 output OGC; 
 output OGD; 
 output OGE; 
 output OHA; 
 output OHB; 
 output OHC; 
 output OHD; 
 output OHE; 
 output OIA; 
 output OIB; 
 output OIC; 
 output OID; 
 output OIE; 
 output OJA; 
 output OJB; 
 output OJC; 
 output OJD; 
 output OJE; 
 output OJF; 
 output OKA; 
 output OKB; 
 output OKC; 
 output OKD; 
 output OKE; 
 output OKF; 
 output OLA; 
 output OLB; 
 output OLC; 
 output OLD; 
 output OLE; 
 output OLF; 
 output OMA; 
 output OMB; 
 output OMC; 
 output OMD; 
 output OME; 
 output OMF; 
 output ONA; 
 output ONB; 
 output ONC; 
 output OND; 
 output ONE; 
 output ONF; 
 output ONG; 
 output ONH; 
 output ONI; 
 output ONJ; 
 output ONK; 
 output ONL; 
 output ONM; 
 output ONN; 
 output ONO; 
 output ONP; 
 output OOA; 
 output OOB; 
 output OOC; 
 output OOD; 
 output OOE; 
 output OOF; 
 output OOG; 
 output OOH; 
 output OOI; 
 output OOJ; 
 output OOK; 
 output OOL; 
 output OOM; 
 output OON; 
 output OOO; 
 output OOP; 
 output OPA; 
 output OPB; 
 output OPC; 
 output OPD; 
 output OPE; 
 output OPF; 
 output OPG; 
 output OPH; 
 output OPI; 
 output OPJ; 
 output OPK; 
 output OPL; 
 output OPM; 
 output OPN; 
 output OPO; 
 output OPP; 
 output OQA; 
 output OQB; 
 output OQC; 
 output OQD; 
 output OQE; 
 output OQF; 
 output OQG; 
 output OQH; 
 output OQI; 
 output OQJ; 
 output OQK; 
 output OQL; 
 output OQM; 
 output OQN; 
 output OQO; 
  
  
reg  AAA ;
reg  AAB ;
reg  AAC ;
reg  AAD ;
reg  AAE ;
reg  AAF ;
reg  AAG ;
reg  AAH ;
reg  AAI ;
reg  AAJ ;
reg  AAK ;
reg  AAL ;
reg  AAM ;
reg  aba ;
reg  abb ;
reg  abc ;
reg  abd ;
reg  abe ;
reg  abf ;
reg  abg ;
reg  abh ;
reg  abi ;
reg  abj ;
reg  abk ;
reg  abl ;
reg  aca ;
reg  acb ;
reg  acc ;
reg  acd ;
reg  ace ;
reg  acf ;
reg  acg ;
reg  ach ;
reg  aci ;
reg  acj ;
reg  ack ;
reg  acl ;
reg  ada ;
reg  adb ;
reg  adc ;
reg  add ;
reg  ade ;
reg  adf ;
reg  adg ;
reg  adh ;
reg  adi ;
reg  adj ;
reg  adk ;
reg  adl ;
reg  AEA ;
reg  AEB ;
reg  AEC ;
reg  AED ;
reg  AEE ;
reg  AEF ;
reg  AEG ;
reg  AEH ;
reg  AEI ;
reg  AEJ ;
reg  AEK ;
reg  AEL ;
reg  baa ;
reg  bab ;
reg  bac ;
reg  bad ;
reg  bae ;
reg  baf ;
reg  bag ;
reg  bah ;
reg  bai ;
reg  baj ;
reg  bak ;
reg  bal ;
reg  caa ;
reg  cab ;
reg  cac ;
reg  cad ;
reg  cae ;
reg  caf ;
reg  cba ;
reg  cbb ;
reg  cbc ;
reg  cbd ;
reg  cbe ;
reg  cbf ;
reg  cbg ;
reg  cbh ;
reg  cca ;
reg  ccb ;
reg  ccc ;
reg  ccd ;
reg  cce ;
reg  ccf ;
reg  ccg ;
reg  cch ;
reg  cci ;
reg  ccj ;
reg  cck ;
reg  ccl ;
reg  DAA ;
reg  DAB ;
reg  DAC ;
reg  DBA ;
reg  DBB ;
reg  DBC ;
reg  DCA ;
reg  DCB ;
reg  DCC ;
reg  DDA ;
reg  DDB ;
reg  DDC ;
reg  DDD ;
reg  DEA ;
reg  DEB ;
reg  DEC ;
reg  DED ;
reg  DFA ;
reg  DFB ;
reg  DFC ;
reg  DFD ;
reg  DGA ;
reg  DGB ;
reg  DGC ;
reg  DGD ;
reg  DHA ;
reg  DHB ;
reg  DHC ;
reg  DHD ;
reg  DIA ;
reg  DIB ;
reg  DIC ;
reg  DID ;
reg  DJA ;
reg  DJB ;
reg  DJC ;
reg  DJD ;
reg  DKA ;
reg  DKB ;
reg  DKC ;
reg  DKD ;
reg  DLA ;
reg  DLB ;
reg  DLC ;
reg  DLD ;
reg  DMA ;
reg  DMB ;
reg  DMC ;
reg  DMD ;
reg  DNA ;
reg  DNB ;
reg  DNC ;
reg  DND ;
reg  DOA ;
reg  DOB ;
reg  DOC ;
reg  DOD ;
reg  DPA ;
reg  DPB ;
reg  DPC ;
reg  DPD ;
reg  DQA ;
reg  DQB ;
reg  DQC ;
reg  DQD ;
reg  DRA ;
reg  DRB ;
reg  DRC ;
reg  DRD ;
reg  GAA ;
reg  GAB ;
reg  GAC ;
reg  GAD ;
reg  GAE ;
reg  GAF ;
reg  GAG ;
reg  GAH ;
reg  GBA ;
reg  GBB ;
reg  GBC ;
reg  GBD ;
reg  GBE ;
reg  GBF ;
reg  GBG ;
reg  GBH ;
reg  GCA ;
reg  GCB ;
reg  GCC ;
reg  GCD ;
reg  GCE ;
reg  GCF ;
reg  GCG ;
reg  GCH ;
reg  GDA ;
reg  GDB ;
reg  GDC ;
reg  GDD ;
reg  GDE ;
reg  GEA ;
reg  GEB ;
reg  GEC ;
reg  GED ;
reg  GEE ;
reg  GEF ;
reg  GEG ;
reg  GEH ;
reg  GFA ;
reg  GFB ;
reg  GFC ;
reg  GFD ;
reg  GFE ;
reg  GFF ;
reg  GFG ;
reg  GFH ;
reg  GGA ;
reg  GGB ;
reg  GGC ;
reg  GGD ;
reg  GGE ;
reg  GGF ;
reg  GGG ;
reg  GGH ;
reg  GHA ;
reg  GHB ;
reg  GHC ;
reg  GHD ;
reg  GHE ;
reg  HAA ;
reg  HAB ;
reg  HAC ;
reg  HAD ;
reg  HAE ;
reg  HAF ;
reg  HBA ;
reg  HBB ;
reg  HBC ;
reg  HBD ;
reg  HBE ;
reg  HBF ;
reg  HCA ;
reg  HCB ;
reg  HCC ;
reg  HCD ;
reg  HCE ;
reg  HCF ;
reg  HDA ;
reg  HDB ;
reg  HDC ;
reg  HDD ;
reg  HDE ;
reg  HDF ;
reg  HEA ;
reg  HEB ;
reg  HEC ;
reg  HED ;
reg  HEE ;
reg  HEF ;
reg  HEG ;
reg  HEH ;
reg  HFA ;
reg  HFB ;
reg  HFC ;
reg  HFD ;
reg  HFE ;
reg  HFF ;
reg  HFG ;
reg  HFH ;
reg  HGA ;
reg  HGB ;
reg  HGC ;
reg  HGD ;
reg  HGE ;
reg  HGF ;
reg  HGG ;
reg  HGH ;
reg  HHA ;
reg  HHB ;
reg  HHC ;
reg  HHD ;
reg  HHE ;
reg  HIA ;
reg  HIB ;
reg  HIC ;
reg  HID ;
reg  HIE ;
reg  HIF ;
reg  HIG ;
reg  HIH ;
reg  HII ;
reg  HIJ ;
reg  HIK ;
reg  HIL ;
reg  HIM ;
reg  HIN ;
reg  HIO ;
reg  HIP ;
reg  HJA ;
reg  HJB ;
reg  HJC ;
reg  HJD ;
reg  HJE ;
reg  HJF ;
reg  HJG ;
reg  HJH ;
reg  HJI ;
reg  HJJ ;
reg  HJK ;
reg  HJL ;
reg  HJM ;
reg  HKA ;
reg  HKB ;
reg  HKC ;
reg  HKD ;
reg  HKE ;
reg  HKF ;
reg  HKG ;
reg  HKH ;
reg  HKI ;
reg  HKJ ;
reg  HKK ;
reg  HKL ;
reg  HKM ;
reg  HKN ;
reg  HKO ;
reg  HKP ;
reg  HLA ;
reg  HLB ;
reg  HLC ;
reg  HLD ;
reg  HLE ;
reg  HLF ;
reg  HLG ;
reg  HLH ;
reg  HLI ;
reg  HLJ ;
reg  HLK ;
reg  HLL ;
reg  HLM ;
reg  NAA ;
reg  NAB ;
reg  NAC ;
reg  NAD ;
reg  NAE ;
reg  NAF ;
reg  NAG ;
reg  NAH ;
reg  NBA ;
reg  NBB ;
reg  NBC ;
reg  NBD ;
reg  NBE ;
reg  NBF ;
reg  NBG ;
reg  NBH ;
reg  NCA ;
reg  NCB ;
reg  NCC ;
reg  NCD ;
reg  NCE ;
reg  NCF ;
reg  NCG ;
reg  NCH ;
reg  NDA ;
reg  NDB ;
reg  NDC ;
reg  NDD ;
reg  NDE ;
reg  NDF ;
reg  NDG ;
reg  NDH ;
reg  OAA ;
reg  OAB ;
reg  OAC ;
reg  OAD ;
reg  OAE ;
reg  OAF ;
reg  OAG ;
reg  OAH ;
reg  OAI ;
reg  OAJ ;
reg  OAK ;
reg  OAL ;
reg  OAM ;
reg  OAN ;
reg  OAO ;
reg  OAP ;
reg  OBA ;
reg  OBB ;
reg  OBC ;
reg  OBD ;
reg  OBE ;
reg  OBF ;
reg  OBG ;
reg  OBH ;
reg  OBI ;
reg  OBJ ;
reg  OBK ;
reg  OBL ;
reg  OBM ;
reg  OBN ;
reg  OBO ;
reg  OBP ;
reg  ODA ;
reg  ODB ;
reg  ODC ;
reg  ODD ;
reg  ODE ;
reg  ODF ;
reg  ODG ;
reg  ODH ;
reg  OEA ;
reg  OEB ;
reg  OEC ;
reg  OED ;
reg  OEE ;
reg  OEF ;
reg  OEG ;
reg  OEH ;
reg  ofa ;
reg  ofb ;
reg  ofc ;
reg  ofd ;
reg  ofe ;
reg  oga ;
reg  ogb ;
reg  ogc ;
reg  ogd ;
reg  oge ;
reg  oha ;
reg  ohb ;
reg  ohc ;
reg  ohd ;
reg  ohe ;
reg  oia ;
reg  oib ;
reg  oic ;
reg  oid ;
reg  oie ;
reg  oja ;
reg  ojb ;
reg  ojc ;
reg  ojd ;
reg  oje ;
reg  ojf ;
reg  oka ;
reg  okb ;
reg  okc ;
reg  okd ;
reg  oke ;
reg  okf ;
reg  ola ;
reg  olb ;
reg  olc ;
reg  old ;
reg  ole ;
reg  olf ;
reg  oma ;
reg  omb ;
reg  omc ;
reg  omd ;
reg  ome ;
reg  omf ;
reg  ona ;
reg  onb ;
reg  onc ;
reg  ond ;
reg  one ;
reg  onf ;
reg  ong ;
reg  onh ;
reg  oni ;
reg  onj ;
reg  onk ;
reg  onl ;
reg  onm ;
reg  onn ;
reg  ono ;
reg  onp ;
reg  ooa ;
reg  oob ;
reg  ooc ;
reg  ood ;
reg  ooe ;
reg  oof ;
reg  oog ;
reg  ooh ;
reg  ooi ;
reg  ooj ;
reg  ook ;
reg  ool ;
reg  oom ;
reg  oon ;
reg  ooo ;
reg  oop ;
reg  OPA ;
reg  OPB ;
reg  OPC ;
reg  OPD ;
reg  OPE ;
reg  OPF ;
reg  OPG ;
reg  OPH ;
reg  OPI ;
reg  OPJ ;
reg  OPK ;
reg  OPL ;
reg  OPM ;
reg  OPN ;
reg  OPO ;
reg  OPP ;
reg  OQA ;
reg  OQB ;
reg  OQC ;
reg  OQD ;
reg  OQE ;
reg  OQF ;
reg  OQG ;
reg  OQH ;
reg  OQI ;
reg  OQJ ;
reg  OQK ;
reg  OQL ;
reg  OQM ;
reg  OQN ;
reg  OQO ;
reg  paa ;
reg  pab ;
reg  pac ;
reg  pad ;
reg  pae ;
reg  paf ;
reg  pag ;
reg  pah ;
reg  pba ;
reg  pbb ;
reg  pbc ;
reg  pbd ;
reg  pbe ;
reg  pbf ;
reg  pbg ;
reg  pbh ;
reg  pca ;
reg  pcb ;
reg  pcc ;
reg  pcd ;
reg  pce ;
reg  pcf ;
reg  pcg ;
reg  pch ;
reg  pda ;
reg  pdb ;
reg  pdc ;
reg  pdd ;
reg  pde ;
reg  pdf ;
reg  pdg ;
reg  pdh ;
reg  QAA ;
reg  QAB ;
reg  QAC ;
reg  QAD ;
reg  qba ;
reg  qbb ;
reg  QBC ;
reg  QBD ;
reg  QCA ;
reg  QCB ;
reg  QCC ;
reg  QCD ;
reg  QDA ;
reg  QDB ;
reg  QDC ;
reg  QDD ;
reg  QEA ;
reg  QEB ;
reg  QEC ;
reg  QED ;
reg  qfa ;
reg  qfb ;
reg  TAA ;
reg  TAB ;
reg  TAC ;
reg  TAD ;
reg  TAE ;
reg  TAF ;
reg  TAG ;
reg  TAH ;
reg  tba ;
reg  tbb ;
reg  tbc ;
reg  tbd ;
reg  tca ;
reg  tcb ;
reg  tcc ;
reg  tcd ;
reg  tda ;
reg  tdb ;
reg  tdc ;
reg  tea ;
reg  teb ;
reg  tec ;
reg  ted ;
reg  tfa ;
reg  tfb ;
reg  tfc ;
reg  tga ;
reg  tgb ;
reg  tgc ;
reg  tha ;
reg  thb ;
reg  thc ;
reg  tia ;
reg  tib ;
reg  tic ;
reg  tja ;
reg  tjb ;
reg  tjc ;
reg  TMA ;
reg  TMB ;
reg  TMC ;
reg  TMD ;
reg  tna ;
reg  tnb ;
reg  tnc ;
reg  waa ;
reg  wab ;
reg  wac ;
reg  wad ;
reg  wae ;
reg  waf ;
reg  wag ;
reg  wah ;
reg  wai ;
reg  waj ;
reg  wak ;
reg  wal ;
reg  wam ;
reg  wan ;
reg  wao ;
reg  wap ;
reg  waq ;
reg  war ;
wire  aaa ;
wire  aab ;
wire  aac ;
wire  aad ;
wire  aae ;
wire  aaf ;
wire  aag ;
wire  aah ;
wire  aai ;
wire  aaj ;
wire  aak ;
wire  aal ;
wire  aam ;
wire  ABA ;
wire  ABB ;
wire  ABC ;
wire  ABD ;
wire  ABE ;
wire  ABF ;
wire  ABG ;
wire  ABH ;
wire  ABI ;
wire  ABJ ;
wire  ABK ;
wire  ABL ;
wire  ACA ;
wire  ACB ;
wire  ACC ;
wire  ACD ;
wire  ACE ;
wire  ACF ;
wire  ACG ;
wire  ACH ;
wire  ACI ;
wire  ACJ ;
wire  ACK ;
wire  ACL ;
wire  ADA ;
wire  ADB ;
wire  ADC ;
wire  ADD ;
wire  ADE ;
wire  ADF ;
wire  ADG ;
wire  ADH ;
wire  ADI ;
wire  ADJ ;
wire  ADK ;
wire  ADL ;
wire  aea ;
wire  aeb ;
wire  aec ;
wire  aed ;
wire  aee ;
wire  aef ;
wire  aeg ;
wire  aeh ;
wire  aei ;
wire  aej ;
wire  aek ;
wire  ael ;
wire  BAA ;
wire  BAB ;
wire  BAC ;
wire  BAD ;
wire  BAE ;
wire  BAF ;
wire  BAG ;
wire  BAH ;
wire  BAI ;
wire  BAJ ;
wire  BAK ;
wire  BAL ;
wire  CAA ;
wire  CAB ;
wire  CAC ;
wire  CAD ;
wire  CAE ;
wire  CAF ;
wire  CBA ;
wire  CBB ;
wire  CBC ;
wire  CBD ;
wire  CBE ;
wire  CBF ;
wire  CBG ;
wire  CBH ;
wire  CCA ;
wire  CCB ;
wire  CCC ;
wire  CCD ;
wire  CCE ;
wire  CCF ;
wire  CCG ;
wire  CCH ;
wire  CCI ;
wire  CCJ ;
wire  CCK ;
wire  CCL ;
wire  daa ;
wire  dab ;
wire  dac ;
wire  dba ;
wire  dbb ;
wire  dbc ;
wire  dca ;
wire  dcb ;
wire  dcc ;
wire  dda ;
wire  ddb ;
wire  ddc ;
wire  ddd ;
wire  dea ;
wire  deb ;
wire  dec ;
wire  ded ;
wire  dfa ;
wire  dfb ;
wire  dfc ;
wire  dfd ;
wire  dga ;
wire  dgb ;
wire  dgc ;
wire  dgd ;
wire  dha ;
wire  dhb ;
wire  dhc ;
wire  dhd ;
wire  dia ;
wire  dib ;
wire  dic ;
wire  did ;
wire  dja ;
wire  djb ;
wire  djc ;
wire  djd ;
wire  dka ;
wire  dkb ;
wire  dkc ;
wire  dkd ;
wire  dla ;
wire  dlb ;
wire  dlc ;
wire  dld ;
wire  dma ;
wire  dmb ;
wire  dmc ;
wire  dmd ;
wire  dna ;
wire  dnb ;
wire  dnc ;
wire  dnd ;
wire  doa ;
wire  dob ;
wire  doc ;
wire  dod ;
wire  dpa ;
wire  dpb ;
wire  dpc ;
wire  dpd ;
wire  dqa ;
wire  dqb ;
wire  dqc ;
wire  dqd ;
wire  dra ;
wire  drb ;
wire  drc ;
wire  drd ;
wire  eaa ;
wire  EAA ;
wire  eab ;
wire  EAB ;
wire  eac ;
wire  EAC ;
wire  ead ;
wire  EAD ;
wire  eae ;
wire  EAE ;
wire  eaf ;
wire  EAF ;
wire  eag ;
wire  EAG ;
wire  eah ;
wire  EAH ;
wire  eba ;
wire  EBA ;
wire  ebb ;
wire  EBB ;
wire  ebc ;
wire  EBC ;
wire  ebd ;
wire  EBD ;
wire  ebe ;
wire  EBE ;
wire  ebf ;
wire  EBF ;
wire  ebg ;
wire  EBG ;
wire  ebh ;
wire  EBH ;
wire  eca ;
wire  ECA ;
wire  ecb ;
wire  ECB ;
wire  ecc ;
wire  ECC ;
wire  ecd ;
wire  ECD ;
wire  ece ;
wire  ECE ;
wire  ecf ;
wire  ECF ;
wire  ecg ;
wire  ECG ;
wire  ech ;
wire  ECH ;
wire  eda ;
wire  EDA ;
wire  edb ;
wire  EDB ;
wire  edc ;
wire  EDC ;
wire  edd ;
wire  EDD ;
wire  ede ;
wire  EDE ;
wire  edf ;
wire  EDF ;
wire  edg ;
wire  EDG ;
wire  edh ;
wire  EDH ;
wire  FAA ;
wire  FAB ;
wire  FAC ;
wire  FAD ;
wire  FAE ;
wire  FAF ;
wire  FAG ;
wire  FAH ;
wire  FAI ;
wire  FBA ;
wire  FBB ;
wire  FBC ;
wire  FBD ;
wire  FBE ;
wire  FBF ;
wire  FBG ;
wire  FBH ;
wire  FBI ;
wire  FCA ;
wire  FCB ;
wire  FCC ;
wire  FCD ;
wire  FCE ;
wire  FCF ;
wire  FCG ;
wire  FCH ;
wire  FCI ;
wire  FDA ;
wire  FDB ;
wire  FDC ;
wire  FDD ;
wire  FDE ;
wire  FDF ;
wire  FDG ;
wire  FDH ;
wire  FDI ;
wire  FEA ;
wire  FEB ;
wire  FEC ;
wire  FED ;
wire  FEE ;
wire  FEF ;
wire  FEG ;
wire  FEH ;
wire  FEI ;
wire  FFA ;
wire  FFB ;
wire  FFC ;
wire  FFD ;
wire  FFE ;
wire  FFF ;
wire  FFG ;
wire  FFH ;
wire  FFI ;
wire  FGA ;
wire  FGB ;
wire  FGC ;
wire  FGD ;
wire  FGE ;
wire  FGF ;
wire  FGG ;
wire  FGH ;
wire  FGI ;
wire  FHA ;
wire  FHB ;
wire  FHC ;
wire  FHD ;
wire  FHE ;
wire  FHF ;
wire  FHG ;
wire  FHH ;
wire  FHI ;
wire  gaa ;
wire  gab ;
wire  gac ;
wire  gad ;
wire  gae ;
wire  gaf ;
wire  gag ;
wire  gah ;
wire  gba ;
wire  gbb ;
wire  gbc ;
wire  gbd ;
wire  gbe ;
wire  gbf ;
wire  gbg ;
wire  gbh ;
wire  gca ;
wire  gcb ;
wire  gcc ;
wire  gcd ;
wire  gce ;
wire  gcf ;
wire  gcg ;
wire  gch ;
wire  gda ;
wire  gdb ;
wire  gdc ;
wire  gdd ;
wire  gde ;
wire  gea ;
wire  geb ;
wire  gec ;
wire  ged ;
wire  gee ;
wire  gef ;
wire  geg ;
wire  geh ;
wire  gfa ;
wire  gfb ;
wire  gfc ;
wire  gfd ;
wire  gfe ;
wire  gff ;
wire  gfg ;
wire  gfh ;
wire  gga ;
wire  ggb ;
wire  ggc ;
wire  ggd ;
wire  gge ;
wire  ggf ;
wire  ggg ;
wire  ggh ;
wire  gha ;
wire  ghb ;
wire  ghc ;
wire  ghd ;
wire  ghe ;
wire  haa ;
wire  hab ;
wire  hac ;
wire  had ;
wire  hae ;
wire  haf ;
wire  hba ;
wire  hbb ;
wire  hbc ;
wire  hbd ;
wire  hbe ;
wire  hbf ;
wire  hca ;
wire  hcb ;
wire  hcc ;
wire  hcd ;
wire  hce ;
wire  hcf ;
wire  hda ;
wire  hdb ;
wire  hdc ;
wire  hdd ;
wire  hde ;
wire  hdf ;
wire  hea ;
wire  heb ;
wire  hec ;
wire  hed ;
wire  hee ;
wire  hef ;
wire  heg ;
wire  heh ;
wire  hfa ;
wire  hfb ;
wire  hfc ;
wire  hfd ;
wire  hfe ;
wire  hff ;
wire  hfg ;
wire  hfh ;
wire  hga ;
wire  hgb ;
wire  hgc ;
wire  hgd ;
wire  hge ;
wire  hgf ;
wire  hgg ;
wire  hgh ;
wire  hha ;
wire  hhb ;
wire  hhc ;
wire  hhd ;
wire  hhe ;
wire  hia ;
wire  hib ;
wire  hic ;
wire  hid ;
wire  hie ;
wire  hif ;
wire  hig ;
wire  hih ;
wire  hii ;
wire  hij ;
wire  hik ;
wire  hil ;
wire  him ;
wire  hin ;
wire  hio ;
wire  hip ;
wire  hja ;
wire  hjb ;
wire  hjc ;
wire  hjd ;
wire  hje ;
wire  hjf ;
wire  hjg ;
wire  hjh ;
wire  hji ;
wire  hjj ;
wire  hjk ;
wire  hjl ;
wire  hjm ;
wire  hka ;
wire  hkb ;
wire  hkc ;
wire  hkd ;
wire  hke ;
wire  hkf ;
wire  hkg ;
wire  hkh ;
wire  hki ;
wire  hkj ;
wire  hkk ;
wire  hkl ;
wire  hkm ;
wire  hkn ;
wire  hko ;
wire  hkp ;
wire  hla ;
wire  hlb ;
wire  hlc ;
wire  hld ;
wire  hle ;
wire  hlf ;
wire  hlg ;
wire  hlh ;
wire  hli ;
wire  hlj ;
wire  hlk ;
wire  hll ;
wire  hlm ;
wire  iaa ;
wire  iab ;
wire  iac ;
wire  iad ;
wire  iae ;
wire  iaf ;
wire  iag ;
wire  iah ;
wire  iai ;
wire  iaj ;
wire  iak ;
wire  ial ;
wire  iba ;
wire  ibb ;
wire  ibc ;
wire  ibd ;
wire  ibe ;
wire  ibf ;
wire  ibg ;
wire  ibh ;
wire  ibi ;
wire  ibj ;
wire  ibk ;
wire  ibl ;
wire  ica ;
wire  icb ;
wire  icc ;
wire  icd ;
wire  ice ;
wire  icf ;
wire  icg ;
wire  ich ;
wire  ici ;
wire  icj ;
wire  ick ;
wire  icl ;
wire  ida ;
wire  idb ;
wire  idc ;
wire  idd ;
wire  ide ;
wire  idf ;
wire  idg ;
wire  idh ;
wire  idi ;
wire  idj ;
wire  idk ;
wire  idl ;
wire  iea ;
wire  ieb ;
wire  iec ;
wire  ied ;
wire  iee ;
wire  ief ;
wire  ieg ;
wire  ieh ;
wire  iei ;
wire  iej ;
wire  iek ;
wire  iel ;
wire  iem ;
wire  ien ;
wire  ieo ;
wire  iep ;
wire  ieq ;
wire  ier ;
wire  ies ;
wire  iet ;
wire  ieu ;
wire  iev ;
wire  iew ;
wire  iex ;
wire  ifa ;
wire  ifb ;
wire  ifc ;
wire  ifd ;
wire  ife ;
wire  iga ;
wire  igb ;
wire  igc ;
wire  ija ;
wire  ijb ;
wire  ijc ;
wire  ijd ;
wire  ije ;
wire  ijf ;
wire  ijg ;
wire  ijh ;
wire  iji ;
wire  ijj ;
wire  ijk ;
wire  ijl ;
wire  ijm ;
wire  ijn ;
wire  ijo ;
wire  ijp ;
wire  ika ;
wire  ikb ;
wire  ikc ;
wire  ikd ;
wire  ike ;
wire  ikf ;
wire  ikg ;
wire  ikh ;
wire  iki ;
wire  ikj ;
wire  ikk ;
wire  ikl ;
wire  ikm ;
wire  ikn ;
wire  iko ;
wire  ikp ;
wire  jaa ;
wire  JAA ;
wire  jab ;
wire  JAB ;
wire  jba ;
wire  JBA ;
wire  jbb ;
wire  JBB ;
wire  jbc ;
wire  JBC ;
wire  jbd ;
wire  JBD ;
wire  jbe ;
wire  JBE ;
wire  jbf ;
wire  JBF ;
wire  jbg ;
wire  JBG ;
wire  jbh ;
wire  JBH ;
wire  jbi ;
wire  JBI ;
wire  jbj ;
wire  JBJ ;
wire  jbk ;
wire  JBK ;
wire  jbl ;
wire  JBL ;
wire  jca ;
wire  JCA ;
wire  jcb ;
wire  JCB ;
wire  jcc ;
wire  JCC ;
wire  jme ;
wire  JME ;
wire  kaa ;
wire  KAA ;
wire  kab ;
wire  KAB ;
wire  kac ;
wire  KAC ;
wire  kba ;
wire  KBA ;
wire  kbb ;
wire  KBB ;
wire  kbc ;
wire  KBC ;
wire  kbd ;
wire  KBD ;
wire  kca ;
wire  KCA ;
wire  kcb ;
wire  KCB ;
wire  kcc ;
wire  KCC ;
wire  kcd ;
wire  KCD ;
wire  laa ;
wire  LAA ;
wire  lab ;
wire  LAB ;
wire  lac ;
wire  LAC ;
wire  lad ;
wire  LAD ;
wire  lae ;
wire  LAE ;
wire  laf ;
wire  LAF ;
wire  lag ;
wire  LAG ;
wire  lah ;
wire  LAH ;
wire  naa ;
wire  nab ;
wire  nac ;
wire  nad ;
wire  nae ;
wire  naf ;
wire  nag ;
wire  nah ;
wire  nba ;
wire  nbb ;
wire  nbc ;
wire  nbd ;
wire  nbe ;
wire  nbf ;
wire  nbg ;
wire  nbh ;
wire  nca ;
wire  ncb ;
wire  ncc ;
wire  ncd ;
wire  nce ;
wire  ncf ;
wire  ncg ;
wire  nch ;
wire  nda ;
wire  ndb ;
wire  ndc ;
wire  ndd ;
wire  nde ;
wire  ndf ;
wire  ndg ;
wire  ndh ;
wire  oaa ;
wire  oab ;
wire  oac ;
wire  oad ;
wire  oae ;
wire  oaf ;
wire  oag ;
wire  oah ;
wire  oai ;
wire  oaj ;
wire  oak ;
wire  oal ;
wire  oam ;
wire  oan ;
wire  oao ;
wire  oap ;
wire  oba ;
wire  obb ;
wire  obc ;
wire  obd ;
wire  obe ;
wire  obf ;
wire  obg ;
wire  obh ;
wire  obi ;
wire  obj ;
wire  obk ;
wire  obl ;
wire  obm ;
wire  obn ;
wire  obo ;
wire  obp ;
wire  oda ;
wire  odb ;
wire  odc ;
wire  odd ;
wire  ode ;
wire  odf ;
wire  odg ;
wire  odh ;
wire  oea ;
wire  oeb ;
wire  oec ;
wire  oed ;
wire  oee ;
wire  oef ;
wire  oeg ;
wire  oeh ;
wire  OFA ;
wire  OFB ;
wire  OFC ;
wire  OFD ;
wire  OFE ;
wire  OGA ;
wire  OGB ;
wire  OGC ;
wire  OGD ;
wire  OGE ;
wire  OHA ;
wire  OHB ;
wire  OHC ;
wire  OHD ;
wire  OHE ;
wire  OIA ;
wire  OIB ;
wire  OIC ;
wire  OID ;
wire  OIE ;
wire  OJA ;
wire  OJB ;
wire  OJC ;
wire  OJD ;
wire  OJE ;
wire  OJF ;
wire  OKA ;
wire  OKB ;
wire  OKC ;
wire  OKD ;
wire  OKE ;
wire  OKF ;
wire  OLA ;
wire  OLB ;
wire  OLC ;
wire  OLD ;
wire  OLE ;
wire  OLF ;
wire  OMA ;
wire  OMB ;
wire  OMC ;
wire  OMD ;
wire  OME ;
wire  OMF ;
wire  ONA ;
wire  ONB ;
wire  ONC ;
wire  OND ;
wire  ONE ;
wire  ONF ;
wire  ONG ;
wire  ONH ;
wire  ONI ;
wire  ONJ ;
wire  ONK ;
wire  ONL ;
wire  ONM ;
wire  ONN ;
wire  ONO ;
wire  ONP ;
wire  OOA ;
wire  OOB ;
wire  OOC ;
wire  OOD ;
wire  OOE ;
wire  OOF ;
wire  OOG ;
wire  OOH ;
wire  OOI ;
wire  OOJ ;
wire  OOK ;
wire  OOL ;
wire  OOM ;
wire  OON ;
wire  OOO ;
wire  OOP ;
wire  opa ;
wire  opb ;
wire  opc ;
wire  opd ;
wire  ope ;
wire  opf ;
wire  opg ;
wire  oph ;
wire  opi ;
wire  opj ;
wire  opk ;
wire  opl ;
wire  opm ;
wire  opn ;
wire  opo ;
wire  opp ;
wire  oqa ;
wire  oqb ;
wire  oqc ;
wire  oqd ;
wire  oqe ;
wire  oqf ;
wire  oqg ;
wire  oqh ;
wire  oqi ;
wire  oqj ;
wire  oqk ;
wire  oql ;
wire  oqm ;
wire  oqn ;
wire  oqo ;
wire  PAA ;
wire  PAB ;
wire  PAC ;
wire  PAD ;
wire  PAE ;
wire  PAF ;
wire  PAG ;
wire  PAH ;
wire  PBA ;
wire  PBB ;
wire  PBC ;
wire  PBD ;
wire  PBE ;
wire  PBF ;
wire  PBG ;
wire  PBH ;
wire  PCA ;
wire  PCB ;
wire  PCC ;
wire  PCD ;
wire  PCE ;
wire  PCF ;
wire  PCG ;
wire  PCH ;
wire  PDA ;
wire  PDB ;
wire  PDC ;
wire  PDD ;
wire  PDE ;
wire  PDF ;
wire  PDG ;
wire  PDH ;
wire  qaa ;
wire  qab ;
wire  qac ;
wire  qad ;
wire  QBA ;
wire  QBB ;
wire  qbc ;
wire  qbd ;
wire  qca ;
wire  qcb ;
wire  qcc ;
wire  qcd ;
wire  qda ;
wire  qdb ;
wire  qdc ;
wire  qdd ;
wire  qea ;
wire  qeb ;
wire  qec ;
wire  qed ;
wire  QFA ;
wire  QFB ;
wire  taa ;
wire  tab ;
wire  tac ;
wire  tad ;
wire  tae ;
wire  taf ;
wire  tag ;
wire  tah ;
wire  TBA ;
wire  TBB ;
wire  TBC ;
wire  TBD ;
wire  TCA ;
wire  TCB ;
wire  TCC ;
wire  TCD ;
wire  TDA ;
wire  TDB ;
wire  TDC ;
wire  TEA ;
wire  TEB ;
wire  TEC ;
wire  TED ;
wire  TFA ;
wire  TFB ;
wire  TFC ;
wire  TGA ;
wire  TGB ;
wire  TGC ;
wire  THA ;
wire  THB ;
wire  THC ;
wire  TIA ;
wire  TIB ;
wire  TIC ;
wire  TJA ;
wire  TJB ;
wire  TJC ;
wire  tma ;
wire  tmb ;
wire  tmc ;
wire  tmd ;
wire  TNA ;
wire  TNB ;
wire  TNC ;
wire  WAA ;
wire  WAB ;
wire  WAC ;
wire  WAD ;
wire  WAE ;
wire  WAF ;
wire  WAG ;
wire  WAH ;
wire  WAI ;
wire  WAJ ;
wire  WAK ;
wire  WAL ;
wire  WAM ;
wire  WAN ;
wire  WAO ;
wire  WAP ;
wire  WAQ ;
wire  WAR ;
wire RAA;
wire RAB;
wire RAC;
wire RAD;
wire RAE;
wire RAF;
wire RAG;
wire RAH;
wire RBA;
wire RBB;
wire RBC;
wire RBD;
wire RBE;
wire RBF;
wire RBG;
wire RBH;
wire RCA;
wire RCB;
wire RCC;
wire RCD;
wire RCE;
wire RCF;
wire RCG;
wire RCH;
wire RDA;
wire RDB;
wire RDC;
wire RDD;
wire RDE;
wire RDF;
wire RDG;
wire RDH;
wire REA;
wire REB;
wire REC;
wire RED;
wire REE;
wire REFF;
wire REG;
wire REH;
wire RFA;
wire RFB;
wire RFC;
wire RFD;
wire RFE;
wire RFF;
wire RFG;
wire RFH;
wire RGA;
wire RGB;
wire RGC;
wire RGD;
wire RGE;
wire RGF;
wire RGG;
wire RGH;
wire RHA;
wire RHB;
wire RHC;
wire RHD;
wire RHE;
wire RHF;
wire RHG;
wire RHH;
wire RIA;
wire RIB;
wire RIC;
wire RID;
wire RIE;
wire RIF;
wire RIG;
wire RIH;
wire RJA;
wire RJB;
wire RJC;
wire RJD;
wire RJE;
wire RJF;
wire RJG;
wire RJH;
wire RKA;
wire RKB;
wire RKC;
wire RKD;
wire RKE;
wire RKF;
wire RKG;
wire RKH;
wire RLA;
wire RLB;
wire RLC;
wire RLD;
wire RLE;
wire RLF;
wire RLG;
wire RLH;
wire RMA;
wire RMB;
wire RMC;
wire RMD;
wire RME;
wire RMF;
wire RMG;
wire RMH;
wire RNA;
wire RNB;
wire RNC;
wire RND;
wire RNE;
wire RNF;
wire RNG;
wire RNH;
wire ROA;
wire ROB;
wire ROC;
wire ROD;
wire ROE;
wire ROF;
wire ROG;
wire ROH;
wire RPA;
wire RPB;
wire RPC;
wire RPD;
wire RQA;
wire RQB;
wire RQC;
wire RQD;
wire RRA;
wire RRB;
wire RRC;
wire RRD; 
wire RPE;
wire RQE;
wire RRE;
   
wire  ZZI ;
wire  ZZO ;
assign ZZI = 1'b1;
assign ZZO = 1'b0;
assign dac = ~DAC;  //complement 
assign dab = ~DAB;  //complement 
assign daa = ~DAA;  //complement 
assign haa = ~HAA;  //complement 
assign hab = ~HAB;  //complement 
assign WAA = ~waa;  //complement 
assign TDB = ~tdb;  //complement 
assign hae = ~HAE;  //complement 
assign haf = ~HAF;  //complement 
assign KAA =  QCD  ; 
assign kaa = ~KAA;  //complement  
assign JCA =  QCD & CAF & cae & CAD  ; 
assign jca = ~JCA;  //complement 
assign CAA = ~caa;  //complement 
assign CAD = ~cad;  //complement 
assign dgb = ~DGB;  //complement 
assign dga = ~DGA;  //complement 
assign dgc = ~DGC;  //complement 
assign dgd = ~DGD;  //complement 
assign hea = ~HEA;  //complement 
assign heb = ~HEB;  //complement 
assign CCI = ~cci;  //complement 
assign THB = ~thb;  //complement 
assign WAG = ~wag;  //complement 
assign TGB = ~tgb;  //complement 
assign WAJ = ~waj;  //complement 
assign hee = ~HEE;  //complement 
assign hef = ~HEF;  //complement 
assign dja = ~DJA;  //complement 
assign djb = ~DJB;  //complement 
assign djc = ~DJC;  //complement 
assign djd = ~DJD;  //complement 
assign hfa = ~HFA;  //complement 
assign hfb = ~HFB;  //complement 
assign KCA =  QED  ; 
assign kca = ~KCA;  //complement  
assign CCA = ~cca;  //complement 
assign CCE = ~cce;  //complement 
assign hfe = ~HFE;  //complement 
assign hff = ~HFF;  //complement 
assign PAA = ~paa;  //complement 
assign EAA =  paa & naa  ; 
assign eaa = ~EAA;  //complement 
assign PBA = ~pba;  //complement 
assign JBA =  ADA & qbc  ; 
assign jba = ~JBA;  //complement 
assign JBG =  ADG & qbd  ; 
assign jbg = ~JBG;  //complement 
assign EBA =  pba & nba  ; 
assign eba = ~EBA;  //complement 
assign PCA = ~pca;  //complement 
assign ECA =  pca & nca  ; 
assign eca = ~ECA;  //complement 
assign PDA = ~pda;  //complement 
assign EDA =  pda & nda  ; 
assign eda = ~EDA;  //complement 
assign ged = ~GED;  //complement 
assign gea = ~GEA;  //complement 
assign geb = ~GEB;  //complement 
assign gec = ~GEC;  //complement 
assign hid = ~HID;  //complement 
assign hia = ~HIA;  //complement 
assign hib = ~HIB;  //complement 
assign hic = ~HIC;  //complement 
assign naa = ~NAA;  //complement 
assign oaa = ~OAA;  //complement 
assign ADA = ~ada;  //complement 
assign ADG = ~adg;  //complement 
assign aag = ~AAG;  //complement 
assign FAA = ~AAI & ~AAH & ~AAG & aam & AAK ; 
assign FAB = ~AAI & ~AAH &  AAG & aam & AAK ; 
assign FAC = ~AAI &  AAH & ~AAG & aam & AAK ; 
assign FAD = ~AAI &  AAH &  AAG & aam & AAK ; 
assign FAE =  AAI & ~AAH & ~AAG & aam & AAK ; 
assign FAF =  AAI & ~AAH &  AAG & aam & AAK ; 
assign FAG =  AAI &  AAH & ~AAG & aam & AAK ; 
assign FAH =  AAI &  AAH &  AAG & aam & AAK ; 
assign FAI = ZZI ; 
assign nba = ~NBA;  //complement 
assign oai = ~OAI;  //complement 
assign aaa = ~AAA;  //complement 
assign laa =  naa & nba & nca & nda  ; 
assign LAA = ~laa;  //complement  
assign nca = ~NCA;  //complement 
assign oba = ~OBA;  //complement 
assign BAA = ~baa;  //complement 
assign BAG = ~bag;  //complement 
assign oda = ~ODA;  //complement 
assign oea = ~OEA;  //complement 
assign nda = ~NDA;  //complement 
assign obi = ~OBI;  //complement 
assign opf = ~OPF;  //complement 
assign gad = ~GAD;  //complement 
assign gaa = ~GAA;  //complement 
assign gab = ~GAB;  //complement 
assign gac = ~GAC;  //complement 
assign OFA = ~ofa;  //complement 
assign OGA = ~oga;  //complement 
assign OIA = ~oia;  //complement 
assign OHA = ~oha;  //complement 
assign ACG = ~acg;  //complement 
assign ABA = ~aba;  //complement 
assign ACA = ~aca;  //complement 
assign ABG = ~abg;  //complement 
assign OJA = ~oja;  //complement 
assign OKA = ~oka;  //complement 
assign OLA = ~ola;  //complement 
assign OMA = ~oma;  //complement 
assign hkd = ~HKD;  //complement 
assign hka = ~HKA;  //complement 
assign hkb = ~HKB;  //complement 
assign hkc = ~HKC;  //complement 
assign opc = ~OPC;  //complement 
assign opd = ~OPD;  //complement 
assign ope = ~OPE;  //complement 
assign ONA = ~ona;  //complement 
assign ONB = ~onb;  //complement 
assign ONC = ~onc;  //complement 
assign dbc = ~DBC;  //complement 
assign dbb = ~DBB;  //complement 
assign dba = ~DBA;  //complement 
assign hac = ~HAC;  //complement 
assign had = ~HAD;  //complement 
assign WAB = ~wab;  //complement 
assign TDC = ~tdc;  //complement 
assign KAB =  QCD & CAD  ; 
assign kab = ~KAB;  //complement  
assign CAB = ~cab;  //complement 
assign CAE = ~cae;  //complement 
assign dka = ~DKA;  //complement 
assign dkb = ~DKB;  //complement 
assign dha = ~DHA;  //complement 
assign dhb = ~DHB;  //complement 
assign dhc = ~DHC;  //complement 
assign dhd = ~DHD;  //complement 
assign hec = ~HEC;  //complement 
assign hed = ~HED;  //complement 
assign CCJ = ~ccj;  //complement 
assign THC = ~thc;  //complement 
assign WAH = ~wah;  //complement 
assign TGC = ~tgc;  //complement 
assign WAK = ~wak;  //complement 
assign heg = ~HEG;  //complement 
assign heh = ~HEH;  //complement 
assign dkc = ~DKC;  //complement 
assign dkd = ~DKD;  //complement 
assign hfc = ~HFC;  //complement 
assign hfd = ~HFD;  //complement 
assign KCB =  QED & CCI  ; 
assign kcb = ~KCB;  //complement  
assign CCB = ~ccb;  //complement 
assign CCF = ~ccf;  //complement 
assign hfg = ~HFG;  //complement 
assign hfh = ~HFH;  //complement 
assign PAB = ~pab;  //complement 
assign EAB =  pab & nab  ; 
assign eab = ~EAB;  //complement 
assign PBB = ~pbb;  //complement 
assign JBB =  ADB & qbc  ; 
assign jbb = ~JBB;  //complement 
assign JBH =  ADH & qbd  ; 
assign jbh = ~JBH;  //complement 
assign EBB =  pbb & nbb  ; 
assign ebb = ~EBB;  //complement 
assign PCB = ~pcb;  //complement 
assign ECB =  pcb & ncb  ; 
assign ecb = ~ECB;  //complement 
assign PDB = ~pdb;  //complement 
assign EDB =  pdb & ndb  ; 
assign edb = ~EDB;  //complement 
assign geh = ~GEH;  //complement 
assign gee = ~GEE;  //complement 
assign gef = ~GEF;  //complement 
assign geg = ~GEG;  //complement 
assign hih = ~HIH;  //complement 
assign hie = ~HIE;  //complement 
assign hif = ~HIF;  //complement 
assign hig = ~HIG;  //complement 
assign nab = ~NAB;  //complement 
assign oab = ~OAB;  //complement 
assign ADB = ~adb;  //complement 
assign ADH = ~adh;  //complement 
assign aah = ~AAH;  //complement 
assign FBA = ~AAI & ~AAH & ~AAG & AAJ & AAK ; 
assign FBB = ~AAI & ~AAH &  AAG & AAJ & AAK ; 
assign FBC = ~AAI &  AAH & ~AAG & AAJ & AAK ; 
assign FBD = ~AAI &  AAH &  AAG & AAJ & AAK ; 
assign FBE =  AAI & ~AAH & ~AAG & AAJ & AAK ; 
assign FBF =  AAI & ~AAH &  AAG & AAJ & AAK ; 
assign FBG =  AAI &  AAH & ~AAG & AAJ & AAK ; 
assign FBH =  AAI &  AAH &  AAG & AAJ & AAK ; 
assign FBI = ZZI ; 
assign nbb = ~NBB;  //complement 
assign oaj = ~OAJ;  //complement 
assign lab =  nab & nbb & ncb & ndb  ; 
assign LAB = ~lab;  //complement  
assign ncb = ~NCB;  //complement 
assign obb = ~OBB;  //complement 
assign ACH = ~ach;  //complement 
assign ABB = ~abb;  //complement 
assign ACB = ~acb;  //complement 
assign ABH = ~abh;  //complement 
assign BAB = ~bab;  //complement 
assign BAH = ~bah;  //complement 
assign odb = ~ODB;  //complement 
assign oeb = ~OEB;  //complement 
assign ndb = ~NDB;  //complement 
assign obj = ~OBJ;  //complement 
assign gah = ~GAH;  //complement 
assign gae = ~GAE;  //complement 
assign gaf = ~GAF;  //complement 
assign gag = ~GAG;  //complement 
assign OFB = ~ofb;  //complement 
assign OGB = ~ogb;  //complement 
assign OHB = ~ohb;  //complement 
assign OIB = ~oib;  //complement 
assign OJB = ~ojb;  //complement 
assign OKB = ~okb;  //complement 
assign OLB = ~olb;  //complement 
assign OMB = ~omb;  //complement 
assign hkh = ~HKH;  //complement 
assign hke = ~HKE;  //complement 
assign hkf = ~HKF;  //complement 
assign hkg = ~HKG;  //complement 
assign aab = ~AAB;  //complement 
assign opj = ~OPJ;  //complement 
assign opg = ~OPG;  //complement 
assign oph = ~OPH;  //complement 
assign opi = ~OPI;  //complement 
assign OND = ~ond;  //complement 
assign ONE = ~one;  //complement 
assign ONF = ~onf;  //complement 
assign dcc = ~DCC;  //complement 
assign dcb = ~DCB;  //complement 
assign dca = ~DCA;  //complement 
assign qcb = ~QCB;  //complement 
assign qcc = ~QCC;  //complement 
assign WAC = ~wac;  //complement 
assign TDA = ~tda;  //complement 
assign qca = ~QCA;  //complement 
assign qcd = ~QCD;  //complement 
assign KAC =  QCD & CAD & CAE  ; 
assign kac = ~KAC;  //complement  
assign CAC = ~cac;  //complement 
assign CAF = ~caf;  //complement 
assign dia = ~DIA;  //complement 
assign dib = ~DIB;  //complement 
assign dic = ~DIC;  //complement 
assign did = ~DID;  //complement 
assign CCK = ~cck;  //complement 
assign THA = ~tha;  //complement 
assign WAI = ~wai;  //complement 
assign TGA = ~tga;  //complement 
assign WAL = ~wal;  //complement 
assign dla = ~DLA;  //complement 
assign dlb = ~DLB;  //complement 
assign dlc = ~DLC;  //complement 
assign dld = ~DLD;  //complement 
assign KCC =  QED & CCI & CCJ  ; 
assign kcc = ~KCC;  //complement  
assign CCC = ~ccc;  //complement 
assign CCG = ~ccg;  //complement 
assign aed = ~AED;  //complement 
assign aea = ~AEA;  //complement 
assign aeb = ~AEB;  //complement 
assign aec = ~AEC;  //complement 
assign PAC = ~pac;  //complement 
assign EAC =  pac & nac  ; 
assign eac = ~EAC;  //complement 
assign aee = ~AEE;  //complement 
assign aef = ~AEF;  //complement 
assign PBC = ~pbc;  //complement 
assign JBC =  ADC & qbc  ; 
assign jbc = ~JBC;  //complement 
assign JBI =  ADI & qbd  ; 
assign jbi = ~JBI;  //complement 
assign EBC =  pbc & nbc  ; 
assign ebc = ~EBC;  //complement 
assign PCC = ~pcc;  //complement 
assign ECC =  pcc & ncc  ; 
assign ecc = ~ECC;  //complement 
assign ECH =  pch & nch  ; 
assign ech = ~ECH;  //complement 
assign PDC = ~pdc;  //complement 
assign EDC =  pdc & ndc  ; 
assign edc = ~EDC;  //complement 
assign EDH =  pdh & ndh  ; 
assign edh = ~EDH;  //complement 
assign gfd = ~GFD;  //complement 
assign gfa = ~GFA;  //complement 
assign gfb = ~GFB;  //complement 
assign gfc = ~GFC;  //complement 
assign hil = ~HIL;  //complement 
assign hii = ~HII;  //complement 
assign hij = ~HIJ;  //complement 
assign hik = ~HIK;  //complement 
assign nac = ~NAC;  //complement 
assign oac = ~OAC;  //complement 
assign ADC = ~adc;  //complement 
assign ADI = ~adi;  //complement 
assign aai = ~AAI;  //complement 
assign FCA = ~AAI & ~AAH & ~AAG & aam & AAL ; 
assign FCB = ~AAI & ~AAH &  AAG & aam & AAL ; 
assign FCC = ~AAI &  AAH & ~AAG & aam & AAL ; 
assign FCD = ~AAI &  AAH &  AAG & aam & AAL ; 
assign FCE =  AAI & ~AAH & ~AAG & aam & AAL ; 
assign FCF =  AAI & ~AAH &  AAG & aam & AAL ; 
assign FCG =  AAI &  AAH & ~AAG & aam & AAL ; 
assign FCH =  AAI &  AAH &  AAG & aam & AAL ; 
assign FCI = ZZI ; 
assign nbc = ~NBC;  //complement 
assign oak = ~OAK;  //complement 
assign aac = ~AAC;  //complement 
assign lac =  nac & nbc & ncc & ndc  ; 
assign LAC = ~lac;  //complement  
assign ncc = ~NCC;  //complement 
assign obc = ~OBC;  //complement 
assign ACI = ~aci;  //complement 
assign ACC = ~acc;  //complement 
assign ABI = ~abi;  //complement 
assign BAC = ~bac;  //complement 
assign BAI = ~bai;  //complement 
assign odc = ~ODC;  //complement 
assign oec = ~OEC;  //complement 
assign ndc = ~NDC;  //complement 
assign obk = ~OBK;  //complement 
assign gbd = ~GBD;  //complement 
assign gba = ~GBA;  //complement 
assign gbb = ~GBB;  //complement 
assign gbc = ~GBC;  //complement 
assign OFC = ~ofc;  //complement 
assign OGC = ~ogc;  //complement 
assign OHC = ~ohc;  //complement 
assign OIC = ~oic;  //complement 
assign OJC = ~ojc;  //complement 
assign OKC = ~okc;  //complement 
assign OLC = ~olc;  //complement 
assign OMC = ~omc;  //complement 
assign hkl = ~HKL;  //complement 
assign hki = ~HKI;  //complement 
assign hkj = ~HKJ;  //complement 
assign hkk = ~HKK;  //complement 
assign opn = ~OPN;  //complement 
assign opk = ~OPK;  //complement 
assign opl = ~OPL;  //complement 
assign opm = ~OPM;  //complement 
assign ONG = ~ong;  //complement 
assign ONH = ~onh;  //complement 
assign ONI = ~oni;  //complement 
assign CCD = ~ccd;  //complement 
assign JCB =  QDD & CBH & CBG & cbf & CBE  ; 
assign jcb = ~JCB;  //complement  
assign CCL = ~ccl;  //complement 
assign qea = ~QEA;  //complement 
assign qed = ~QED;  //complement 
assign qeb = ~QEB;  //complement 
assign qec = ~QEC;  //complement 
assign KCD =  QED & CCI & CCJ & CCK  ; 
assign kcd = ~KCD;  //complement  
assign CCH = ~cch;  //complement 
assign PAD = ~pad;  //complement 
assign EAD =  pad & nad  ; 
assign ead = ~EAD;  //complement 
assign gfe = ~GFE;  //complement 
assign PBD = ~pbd;  //complement 
assign JBD =  ADD & qbc  ; 
assign jbd = ~JBD;  //complement 
assign JBJ =  ADJ & qbd  ; 
assign jbj = ~JBJ;  //complement 
assign EBD =  pbd & nbd  ; 
assign ebd = ~EBD;  //complement 
assign PCD = ~pcd;  //complement 
assign ECD =  pcd & ncd  ; 
assign ecd = ~ECD;  //complement 
assign PDD = ~pdd;  //complement 
assign EDD =  pdd & ndd  ; 
assign edd = ~EDD;  //complement 
assign hip = ~HIP;  //complement 
assign him = ~HIM;  //complement 
assign hin = ~HIN;  //complement 
assign hio = ~HIO;  //complement 
assign gfh = ~GFH;  //complement 
assign gff = ~GFF;  //complement 
assign gfg = ~GFG;  //complement 
assign nad = ~NAD;  //complement 
assign oad = ~OAD;  //complement 
assign ADD = ~add;  //complement 
assign ADJ = ~adj;  //complement 
assign aaj = ~AAJ;  //complement 
assign aam = ~AAM;  //complement 
assign FDA = ~AAI & ~AAH & ~AAG & AAJ & AAL ; 
assign FDB = ~AAI & ~AAH &  AAG & AAJ & AAL ; 
assign FDC = ~AAI &  AAH & ~AAG & AAJ & AAL ; 
assign FDD = ~AAI &  AAH &  AAG & AAJ & AAL ; 
assign FDE =  AAI & ~AAH & ~AAG & AAJ & AAL ; 
assign FDF =  AAI & ~AAH &  AAG & AAJ & AAL ; 
assign FDG =  AAI &  AAH & ~AAG & AAJ & AAL ; 
assign FDH =  AAI &  AAH &  AAG & AAJ & AAL ; 
assign FDI = ZZI ; 
assign nbd = ~NBD;  //complement 
assign oal = ~OAL;  //complement 
assign QBA = ~qba;  //complement 
assign aad = ~AAD;  //complement 
assign lad =  nad & nbd & ncd & ndd  ; 
assign LAD = ~lad;  //complement  
assign ncd = ~NCD;  //complement 
assign obd = ~OBD;  //complement 
assign ACJ = ~acj;  //complement 
assign ABD = ~abd;  //complement 
assign ACD = ~acd;  //complement 
assign ABJ = ~abj;  //complement 
assign BAD = ~bad;  //complement 
assign BAJ = ~baj;  //complement 
assign odd = ~ODD;  //complement 
assign oed = ~OED;  //complement 
assign ndd = ~NDD;  //complement 
assign obl = ~OBL;  //complement 
assign gbh = ~GBH;  //complement 
assign gbe = ~GBE;  //complement 
assign gbf = ~GBF;  //complement 
assign gbg = ~GBG;  //complement 
assign OFD = ~ofd;  //complement 
assign OGD = ~ogd;  //complement 
assign OHD = ~ohd;  //complement 
assign OID = ~oid;  //complement 
assign OJD = ~ojd;  //complement 
assign OKD = ~okd;  //complement 
assign OLD = ~old;  //complement 
assign OMD = ~omd;  //complement 
assign hkp = ~HKP;  //complement 
assign hkm = ~HKM;  //complement 
assign hkn = ~HKN;  //complement 
assign hko = ~HKO;  //complement 
assign oqb = ~OQB;  //complement 
assign opo = ~OPO;  //complement 
assign opp = ~OPP;  //complement 
assign oqa = ~OQA;  //complement 
assign ONJ = ~onj;  //complement 
assign ONK = ~onk;  //complement 
assign dda = ~DDA;  //complement 
assign ddb = ~DDB;  //complement 
assign ddc = ~DDC;  //complement 
assign ddd = ~DDD;  //complement 
assign hba = ~HBA;  //complement 
assign hbb = ~HBB;  //complement 
assign WAD = ~wad;  //complement 
assign TFB = ~tfb;  //complement 
assign EBE =  pbe & nbe  ; 
assign ebe = ~EBE;  //complement 
assign KBA =  QDD  ; 
assign kba = ~KBA;  //complement  
assign CBA = ~cba;  //complement 
assign CBE = ~cbe;  //complement 
assign ECE =  pce & nce  ; 
assign ece = ~ECE;  //complement 
assign hbe = ~HBE;  //complement 
assign hbf = ~HBF;  //complement 
assign hhb = ~HHB;  //complement 
assign dmc = ~DMC;  //complement 
assign dmd = ~DMD;  //complement 
assign hga = ~HGA;  //complement 
assign hgb = ~HGB;  //complement 
assign TJB = ~tjb;  //complement 
assign WAM = ~wam;  //complement 
assign TIB = ~tib;  //complement 
assign WAP = ~wap;  //complement 
assign hge = ~HGE;  //complement 
assign hgf = ~HGF;  //complement 
assign dpa = ~DPA;  //complement 
assign dpb = ~DPB;  //complement 
assign dpc = ~DPC;  //complement 
assign dpd = ~DPD;  //complement 
assign hha = ~HHA;  //complement 
assign JCC =  QED & CCL & CCK & ccj & CCI  ; 
assign jcc = ~JCC;  //complement  
assign dma = ~DMA;  //complement 
assign dmb = ~DMB;  //complement 
assign hhe = ~HHE;  //complement 
assign PAE = ~pae;  //complement 
assign EAE =  pae & nae  ; 
assign eae = ~EAE;  //complement 
assign PBE = ~pbe;  //complement 
assign JBE =  ADE & qbc  ; 
assign jbe = ~JBE;  //complement 
assign JBK =  ADK & qbd  ; 
assign jbk = ~JBK;  //complement 
assign PCE = ~pce;  //complement 
assign PDE = ~pde;  //complement 
assign EDE =  pde & nde  ; 
assign ede = ~EDE;  //complement 
assign ggd = ~GGD;  //complement 
assign gga = ~GGA;  //complement 
assign ggb = ~GGB;  //complement 
assign ggc = ~GGC;  //complement 
assign hjd = ~HJD;  //complement 
assign hja = ~HJA;  //complement 
assign hjb = ~HJB;  //complement 
assign hjc = ~HJC;  //complement 
assign hcf = ~HCF;  //complement 
assign hca = ~HCA;  //complement 
assign hcb = ~HCB;  //complement 
assign hce = ~HCE;  //complement 
assign hdf = ~HDF;  //complement 
assign hda = ~HDA;  //complement 
assign hdb = ~HDB;  //complement 
assign hde = ~HDE;  //complement 
assign nae = ~NAE;  //complement 
assign oae = ~OAE;  //complement 
assign ADE = ~ade;  //complement 
assign ADK = ~adk;  //complement 
assign aak = ~AAK;  //complement 
assign FEA = ~HDC & ~HDB & ~HDA & hdd & HDE ; 
assign FEB = ~HDC & ~HDB &  HDA & hdd & HDE ; 
assign FEC = ~HDC &  HDB & ~HDA & hdd & HDE ; 
assign FED = ~HDC &  HDB &  HDA & hdd & HDE ; 
assign FEE =  HDC & ~HDB & ~HDA & hdd & HDE ; 
assign FEF =  HDC & ~HDB &  HDA & hdd & HDE ; 
assign FEG =  HDC &  HDB & ~HDA & hdd & HDE ; 
assign FEH =  HDC &  HDB &  HDA & hdd & HDE ; 
assign FEI = ZZI ; 
assign nbe = ~NBE;  //complement 
assign oam = ~OAM;  //complement 
assign QBB = ~qbb;  //complement 
assign aae = ~AAE;  //complement 
assign lae =  nae & nbe & nce & nde  ; 
assign LAE = ~lae;  //complement  
assign nce = ~NCE;  //complement 
assign obe = ~OBE;  //complement 
assign ACK = ~ack;  //complement 
assign ABE = ~abe;  //complement 
assign ACE = ~ace;  //complement 
assign ABK = ~abk;  //complement 
assign BAE = ~bae;  //complement 
assign BAK = ~bak;  //complement 
assign ode = ~ODE;  //complement 
assign oee = ~OEE;  //complement 
assign nde = ~NDE;  //complement 
assign obm = ~OBM;  //complement 
assign gcd = ~GCD;  //complement 
assign gca = ~GCA;  //complement 
assign gcb = ~GCB;  //complement 
assign gcc = ~GCC;  //complement 
assign ONL = ~onl;  //complement 
assign ONM = ~onm;  //complement 
assign ONN = ~onn;  //complement 
assign OJE = ~oje;  //complement 
assign OKE = ~oke;  //complement 
assign OLE = ~ole;  //complement 
assign OME = ~ome;  //complement 
assign hld = ~HLD;  //complement 
assign hla = ~HLA;  //complement 
assign hlb = ~HLB;  //complement 
assign hlc = ~HLC;  //complement 
assign oqf = ~OQF;  //complement 
assign oqc = ~OQC;  //complement 
assign oqd = ~OQD;  //complement 
assign oqe = ~OQE;  //complement 
assign ONO = ~ono;  //complement 
assign ONP = ~onp;  //complement 
assign dea = ~DEA;  //complement 
assign deb = ~DEB;  //complement 
assign dec = ~DEC;  //complement 
assign ded = ~DED;  //complement 
assign hbc = ~HBC;  //complement 
assign hbd = ~HBD;  //complement 
assign WAE = ~wae;  //complement 
assign TFC = ~tfc;  //complement 
assign KBB =  QDD & CBE  ; 
assign kbb = ~KBB;  //complement  
assign CBB = ~cbb;  //complement 
assign CBF = ~cbf;  //complement 
assign dqb = ~DQB;  //complement 
assign dna = ~DNA;  //complement 
assign dnb = ~DNB;  //complement 
assign dnc = ~DNC;  //complement 
assign dnd = ~DND;  //complement 
assign hgc = ~HGC;  //complement 
assign hgd = ~HGD;  //complement 
assign TJC = ~tjc;  //complement 
assign WAN = ~wan;  //complement 
assign TIC = ~tic;  //complement 
assign WAQ = ~waq;  //complement 
assign hgg = ~HGG;  //complement 
assign hgh = ~HGH;  //complement 
assign dqa = ~DQA;  //complement 
assign dqc = ~DQC;  //complement 
assign dqd = ~DQD;  //complement 
assign hhc = ~HHC;  //complement 
assign hhd = ~HHD;  //complement 
assign PAF = ~paf;  //complement 
assign EAF =  paf & naf  ; 
assign eaf = ~EAF;  //complement 
assign PBF = ~pbf;  //complement 
assign JBF =  ADF & qbc  ; 
assign jbf = ~JBF;  //complement 
assign JBL =  ADL & qbd  ; 
assign jbl = ~JBL;  //complement 
assign EBF =  pbf & nbf  ; 
assign ebf = ~EBF;  //complement 
assign PCF = ~pcf;  //complement 
assign ECF =  pcf & ncf  ; 
assign ecf = ~ECF;  //complement 
assign PDF = ~pdf;  //complement 
assign EDF =  pdf & ndf  ; 
assign edf = ~EDF;  //complement 
assign ggh = ~GGH;  //complement 
assign gge = ~GGE;  //complement 
assign ggf = ~GGF;  //complement 
assign ggg = ~GGG;  //complement 
assign hjh = ~HJH;  //complement 
assign hje = ~HJE;  //complement 
assign hjf = ~HJF;  //complement 
assign hjg = ~HJG;  //complement 
assign hcc = ~HCC;  //complement 
assign hcd = ~HCD;  //complement 
assign hdc = ~HDC;  //complement 
assign hdd = ~HDD;  //complement 
assign naf = ~NAF;  //complement 
assign oaf = ~OAF;  //complement 
assign ADF = ~adf;  //complement 
assign ADL = ~adl;  //complement 
assign ABL = ~abl;  //complement 
assign aal = ~AAL;  //complement 
assign FFA = ~HDC & ~HDB & ~HDA & HDD & HDE ; 
assign FFB = ~HDC & ~HDB &  HDA & HDD & HDE ; 
assign FFC = ~HDC &  HDB & ~HDA & HDD & HDE ; 
assign FFD = ~HDC &  HDB &  HDA & HDD & HDE ; 
assign FFE =  HDC & ~HDB & ~HDA & HDD & HDE ; 
assign FFF =  HDC & ~HDB &  HDA & HDD & HDE ; 
assign FFG =  HDC &  HDB & ~HDA & HDD & HDE ; 
assign FFH =  HDC &  HDB &  HDA & HDD & HDE ; 
assign FFI = ZZI ; 
assign nbf = ~NBF;  //complement 
assign oan = ~OAN;  //complement 
assign laf =  naf & nbf & ncf & ndf  ; 
assign LAF = ~laf;  //complement  
assign ncf = ~NCF;  //complement 
assign obf = ~OBF;  //complement 
assign BAL = ~bal;  //complement 
assign BAF = ~baf;  //complement 
assign odf = ~ODF;  //complement 
assign oef = ~OEF;  //complement 
assign ndf = ~NDF;  //complement 
assign obn = ~OBN;  //complement 
assign gch = ~GCH;  //complement 
assign gce = ~GCE;  //complement 
assign gcf = ~GCF;  //complement 
assign gcg = ~GCG;  //complement 
assign OFE = ~ofe;  //complement 
assign OGE = ~oge;  //complement 
assign OHE = ~ohe;  //complement 
assign OIE = ~oie;  //complement 
assign ACL = ~acl;  //complement 
assign ABC = ~abc;  //complement 
assign ABF = ~abf;  //complement 
assign ACF = ~acf;  //complement 
assign OJF = ~ojf;  //complement 
assign OKF = ~okf;  //complement 
assign OLF = ~olf;  //complement 
assign OMF = ~omf;  //complement 
assign hlh = ~HLH;  //complement 
assign hle = ~HLE;  //complement 
assign hlf = ~HLF;  //complement 
assign hlg = ~HLG;  //complement 
assign aaf = ~AAF;  //complement 
assign oqj = ~OQJ;  //complement 
assign oqg = ~OQG;  //complement 
assign oqh = ~OQH;  //complement 
assign oqi = ~OQI;  //complement 
assign OOA = ~ooa;  //complement 
assign OOB = ~oob;  //complement 
assign OOC = ~ooc;  //complement 
assign dfa = ~DFA;  //complement 
assign dfb = ~DFB;  //complement 
assign dfc = ~DFC;  //complement 
assign dfd = ~DFD;  //complement 
assign qdb = ~QDB;  //complement 
assign qdc = ~QDC;  //complement 
assign WAF = ~waf;  //complement 
assign TFA = ~tfa;  //complement 
assign qda = ~QDA;  //complement 
assign qdd = ~QDD;  //complement 
assign KBC =  QDD & CBE & CBF  ; 
assign kbc = ~KBC;  //complement  
assign CBC = ~cbc;  //complement 
assign CBG = ~cbg;  //complement 
assign doa = ~DOA;  //complement 
assign dob = ~DOB;  //complement 
assign doc = ~DOC;  //complement 
assign dod = ~DOD;  //complement 
assign TJA = ~tja;  //complement 
assign WAO = ~wao;  //complement 
assign TIA = ~tia;  //complement 
assign WAR = ~war;  //complement 
assign drb = ~DRB;  //complement 
assign dra = ~DRA;  //complement 
assign drc = ~DRC;  //complement 
assign drd = ~DRD;  //complement 
assign aej = ~AEJ;  //complement 
assign aeg = ~AEG;  //complement 
assign aeh = ~AEH;  //complement 
assign aei = ~AEI;  //complement 
assign PAG = ~pag;  //complement 
assign EAG =  pag & nag  ; 
assign eag = ~EAG;  //complement 
assign aek = ~AEK;  //complement 
assign ael = ~AEL;  //complement 
assign PBG = ~pbg;  //complement 
assign EBG =  pbg & nbg  ; 
assign ebg = ~EBG;  //complement 
assign PCG = ~pcg;  //complement 
assign ECG =  pcg & ncg  ; 
assign ecg = ~ECG;  //complement 
assign PDG = ~pdg;  //complement 
assign EDG =  pdg & ndg  ; 
assign edg = ~EDG;  //complement 
assign ghd = ~GHD;  //complement 
assign gha = ~GHA;  //complement 
assign ghb = ~GHB;  //complement 
assign ghc = ~GHC;  //complement 
assign hjl = ~HJL;  //complement 
assign hji = ~HJI;  //complement 
assign hjj = ~HJJ;  //complement 
assign hjk = ~HJK;  //complement 
assign nag = ~NAG;  //complement 
assign oag = ~OAG;  //complement 
assign qbc = ~QBC;  //complement 
assign qbd = ~QBD;  //complement 
assign tad = ~TAD;  //complement 
assign taa = ~TAA;  //complement 
assign tab = ~TAB;  //complement 
assign tac = ~TAC;  //complement 
assign FGA = ~HDC & ~HDB & ~HDA & hdd & HDF ; 
assign FGB = ~HDC & ~HDB &  HDA & hdd & HDF ; 
assign FGC = ~HDC &  HDB & ~HDA & hdd & HDF ; 
assign FGD = ~HDC &  HDB &  HDA & hdd & HDF ; 
assign FGE =  HDC & ~HDB & ~HDA & hdd & HDF ; 
assign FGF =  HDC & ~HDB &  HDA & hdd & HDF ; 
assign FGG =  HDC &  HDB & ~HDA & hdd & HDF ; 
assign FGH =  HDC &  HDB &  HDA & hdd & HDF ; 
assign FGI = ZZI ; 
assign nbg = ~NBG;  //complement 
assign oao = ~OAO;  //complement 
assign JAA =  ACK & qba & qbb  |  ACL & qba & qbb  ; 
assign jaa = ~JAA; //complement 
assign JAB =  ACK & qba & qbb  |  ACL & qba & qbb  ; 
assign jab = ~JAB;  //complement 
assign tah = ~TAH;  //complement 
assign tae = ~TAE;  //complement 
assign taf = ~TAF;  //complement 
assign lag =  nag & nbg & ncg & ndg  ; 
assign LAG = ~lag;  //complement  
assign ncg = ~NCG;  //complement 
assign obg = ~OBG;  //complement 
assign odg = ~ODG;  //complement 
assign oeg = ~OEG;  //complement 
assign ndg = ~NDG;  //complement 
assign obo = ~OBO;  //complement 
assign oqm = ~OQM;  //complement 
assign gdd = ~GDD;  //complement 
assign gda = ~GDA;  //complement 
assign gdb = ~GDB;  //complement 
assign gdc = ~GDC;  //complement 
assign OOD = ~ood;  //complement 
assign OOE = ~ooe;  //complement 
assign OOF = ~oof;  //complement 
assign OOG = ~oog;  //complement 
assign OOH = ~ooh;  //complement 
assign OOI = ~ooi;  //complement 
assign hll = ~HLL;  //complement 
assign hli = ~HLI;  //complement 
assign hlj = ~HLJ;  //complement 
assign hlk = ~HLK;  //complement 
assign tag = ~TAG;  //complement 
assign oqn = ~OQN;  //complement 
assign oqk = ~OQK;  //complement 
assign oql = ~OQL;  //complement 
assign OOJ = ~ooj;  //complement 
assign OOK = ~ook;  //complement 
assign KBD =  QDD & CBE & CBF & CBG  ; 
assign kbd = ~KBD;  //complement  
assign CBD = ~cbd;  //complement 
assign CBH = ~cbh;  //complement 
assign PAH = ~pah;  //complement 
assign EAH =  pah & nah  ; 
assign eah = ~EAH;  //complement 
assign ghe = ~GHE;  //complement 
assign PBH = ~pbh;  //complement 
assign EBH =  pbh & nbh  ; 
assign ebh = ~EBH;  //complement 
assign PCH = ~pch;  //complement 
assign PDH = ~pdh;  //complement 
assign hjm = ~HJM;  //complement 
assign TNA = ~tna;  //complement 
assign TNB = ~tnb;  //complement 
assign TNC = ~tnc;  //complement 
assign tmd = ~TMD;  //complement 
assign tma = ~TMA;  //complement 
assign tmb = ~TMB;  //complement 
assign tmc = ~TMC;  //complement 
assign nah = ~NAH;  //complement 
assign oah = ~OAH;  //complement 
assign QFA = ~qfa;  //complement 
assign QFB = ~qfb;  //complement 
assign qad = ~QAD;  //complement 
assign qaa = ~QAA;  //complement 
assign qab = ~QAB;  //complement 
assign qac = ~QAC;  //complement 
assign FHA = ~HDC & ~HDB & ~HDA & HDD & HDF ; 
assign FHB = ~HDC & ~HDB &  HDA & HDD & HDF ; 
assign FHC = ~HDC &  HDB & ~HDA & HDD & HDF ; 
assign FHD = ~HDC &  HDB &  HDA & HDD & HDF ; 
assign FHE =  HDC & ~HDB & ~HDA & HDD & HDF ; 
assign FHF =  HDC & ~HDB &  HDA & HDD & HDF ; 
assign FHG =  HDC &  HDB & ~HDA & HDD & HDF ; 
assign FHH =  HDC &  HDB &  HDA & HDD & HDF ; 
assign FHI = ZZI ; 
assign nbh = ~NBH;  //complement 
assign oap = ~OAP;  //complement 
assign TBD = ~tbd;  //complement 
assign TBA = ~tba;  //complement 
assign lah =  nah & nbh & nch & ndh  ; 
assign LAH = ~lah;  //complement  
assign jme =  tma  ; 
assign JME = ~jme;  //complement 
assign nch = ~NCH;  //complement 
assign obh = ~OBH;  //complement 
assign TCD = ~tcd;  //complement 
assign TCA = ~tca;  //complement 
assign TCB = ~tcb;  //complement 
assign TCC = ~tcc;  //complement 
assign odh = ~ODH;  //complement 
assign oeh = ~OEH;  //complement 
assign ndh = ~NDH;  //complement 
assign obp = ~OBP;  //complement 
assign TED = ~ted;  //complement 
assign TEA = ~tea;  //complement 
assign TEB = ~teb;  //complement 
assign TEC = ~tec;  //complement 
assign OOL = ~ool;  //complement 
assign OOM = ~oom;  //complement 
assign OON = ~oon;  //complement 
assign gde = ~GDE;  //complement 
assign hlm = ~HLM;  //complement 
assign TBB = ~tbb;  //complement 
assign TBC = ~tbc;  //complement 
assign oqo = ~OQO;  //complement 
assign opa = ~OPA;  //complement 
assign opb = ~OPB;  //complement 
assign OOO = ~ooo;  //complement 
assign OOP = ~oop;  //complement 
assign iaa = ~IAA; //complement 
assign iab = ~IAB; //complement 
assign iac = ~IAC; //complement 
assign iad = ~IAD; //complement 
assign iae = ~IAE; //complement 
assign iaf = ~IAF; //complement 
assign iag = ~IAG; //complement 
assign iah = ~IAH; //complement 
assign iai = ~IAI; //complement 
assign iaj = ~IAJ; //complement 
assign iak = ~IAK; //complement 
assign ial = ~IAL; //complement 
assign iba = ~IBA; //complement 
assign ibb = ~IBB; //complement 
assign ibc = ~IBC; //complement 
assign ibd = ~IBD; //complement 
assign ibe = ~IBE; //complement 
assign ibf = ~IBF; //complement 
assign ibg = ~IBG; //complement 
assign ibh = ~IBH; //complement 
assign ibi = ~IBI; //complement 
assign ibj = ~IBJ; //complement 
assign ibk = ~IBK; //complement 
assign ibl = ~IBL; //complement 
assign ica = ~ICA; //complement 
assign icb = ~ICB; //complement 
assign icc = ~ICC; //complement 
assign icd = ~ICD; //complement 
assign ice = ~ICE; //complement 
assign icf = ~ICF; //complement 
assign icg = ~ICG; //complement 
assign ich = ~ICH; //complement 
assign ici = ~ICI; //complement 
assign icj = ~ICJ; //complement 
assign ick = ~ICK; //complement 
assign icl = ~ICL; //complement 
assign ida = ~IDA; //complement 
assign idb = ~IDB; //complement 
assign idc = ~IDC; //complement 
assign idd = ~IDD; //complement 
assign ide = ~IDE; //complement 
assign idf = ~IDF; //complement 
assign idg = ~IDG; //complement 
assign idh = ~IDH; //complement 
assign idi = ~IDI; //complement 
assign idj = ~IDJ; //complement 
assign idk = ~IDK; //complement 
assign idl = ~IDL; //complement 
assign iea = ~IEA; //complement 
assign ieb = ~IEB; //complement 
assign iec = ~IEC; //complement 
assign ied = ~IED; //complement 
assign iee = ~IEE; //complement 
assign ief = ~IEF; //complement 
assign ieg = ~IEG; //complement 
assign ieh = ~IEH; //complement 
assign iei = ~IEI; //complement 
assign iej = ~IEJ; //complement 
assign iek = ~IEK; //complement 
assign iel = ~IEL; //complement 
assign iem = ~IEM; //complement 
assign ien = ~IEN; //complement 
assign ieo = ~IEO; //complement 
assign iep = ~IEP; //complement 
assign ieq = ~IEQ; //complement 
assign ier = ~IER; //complement 
assign ies = ~IES; //complement 
assign iet = ~IET; //complement 
assign ieu = ~IEU; //complement 
assign iev = ~IEV; //complement 
assign iew = ~IEW; //complement 
assign iex = ~IEX; //complement 
assign ifa = ~IFA; //complement 
assign ifb = ~IFB; //complement 
assign ifc = ~IFC; //complement 
assign ifd = ~IFD; //complement 
assign ife = ~IFE; //complement 
assign iga = ~IGA; //complement 
assign igb = ~IGB; //complement 
assign igc = ~IGC; //complement 
assign ija = ~IJA; //complement 
assign ijb = ~IJB; //complement 
assign ijc = ~IJC; //complement 
assign ijd = ~IJD; //complement 
assign ije = ~IJE; //complement 
assign ijf = ~IJF; //complement 
assign ijg = ~IJG; //complement 
assign ijh = ~IJH; //complement 
assign iji = ~IJI; //complement 
assign ijj = ~IJJ; //complement 
assign ijk = ~IJK; //complement 
assign ijl = ~IJL; //complement 
assign ijm = ~IJM; //complement 
assign ijn = ~IJN; //complement 
assign ijo = ~IJO; //complement 
assign ijp = ~IJP; //complement 
assign ika = ~IKA; //complement 
assign ikb = ~IKB; //complement 
assign ikc = ~IKC; //complement 
assign ikd = ~IKD; //complement 
assign ike = ~IKE; //complement 
assign ikf = ~IKF; //complement 
assign ikg = ~IKG; //complement 
assign ikh = ~IKH; //complement 
assign iki = ~IKI; //complement 
assign ikj = ~IKJ; //complement 
assign ikk = ~IKK; //complement 
assign ikl = ~IKL; //complement 
assign ikm = ~IKM; //complement 
assign ikn = ~IKN; //complement 
assign iko = ~IKO; //complement 
assign ikp = ~IKP; //complement 
always@(posedge IZZ )
   begin 
 DAC <= DAC & tdb |  CAC & TDB ; 
 DAB <= DAB & tdb |  CAB & TDB ; 
 DAA <= DAA & tdb |  CAA & TDB ; 
 HAA <=  RAA & TDA  |  RBA & TDB  |  RCA & TDC  ; 
 HAB <=  RAB & TDA  |  RBB & TDB  |  RCB & TDC  ; 
 waa <= qca ; 
 tdb <= qca ; 
 HAE <=  RAE & TDA  |  RBE & TDB  |  RCE & TDC  ; 
 HAF <=  RAF & TDA  |  RBF & TDB  |  RCF & TDC  ; 
 caa <=  caa & kaa  |  CAA & KAA  |  JCA  |  TMA  ; 
 cad <=  caa & kaa  |  CAA & KAA  |  JCA  |  TMA  ; 
 DGB <=  DGB & tgb  |  CCB & TGB  ; 
 DGA <=  DGA & tgb  |  CCA & TGB  ; 
 DGC <=  DGC & tgb  |  CCC & TGB  ; 
 DGD <=  DGD & tgb  |  CCD & TGB  ; 
 HEA <=  RGA & TGA  |  RHA & TGB  |  RIA & TGC  ; 
 HEB <=  RGB & TGA  |  RHB & TGB  |  RIB & TGC  ; 
 cci <= cce ; 
 thb <= qea ; 
 wag <= qea ; 
 tgb <= qea ; 
 waj <= qea ; 
 HEE <=  RGE & TGA  |  RHE & TGB  |  RIE & TGC  ; 
 HEF <=  RGF & TGA  |  RHF & TGB  |  RIF & TGC  ; 
 DJA <=  DJA & thb  |  CCE & THB  ; 
 DJB <=  DJB & thb  |  CCF & THB  ; 
 DJC <=  DJC & thb  |  CCG & THB  ; 
 DJD <=  DJD & thb  |  CCH & THB  ; 
 HFA <=  RJA & THA  |  RKA & THB  |  RLA & THC  ; 
 HFB <=  RJB & THA  |  RKB & THB  |  RLB & THC  ; 
 cca <=  cca & kca  |  CCA & KCA  |  JCC  |  TNC  ; 
 cce <=  cca & kca  |  CCA & KCA  |  JCC  |  TNC  ; 
 HFE <=  RJE & THA  |  RKE & THB  |  RLE & THC  ; 
 HFF <=  RJF & THA  |  RKF & THB  |  RLF & THC  ; 
 paa <=  paa & naa  |  FEA  |  TMA  ; 
 pba <=  pba & nba  |  FFA  |  TMB  ; 
 pca <=  pca & nca  |  FGA  |  TMC  ; 
 pda <=  pda & nda  |  FHA  |  TMD  ; 
 GED <= GAD ; 
 GEA <= GAA ; 
 GEB <= GAB ; 
 GEC <= GAC ; 
 HID <= HED ; 
 HIA <= HEA ; 
 HIB <= HEB ; 
 HIC <= HEC ; 
 NAA <=  FAA & EAA  ; 
 OAA <=  FAA & EAA  ; 
 ada <= aca ; 
 adg <= acg ; 
 AAG <=  IAG & TAE  |  IBG & TAF  |  ICG & TAG  |  IDG & TAH  |  BAG  ; 
 NBA <=  FBA & EBA  ; 
 OAI <=  FBA & EBA  ; 
 AAA <=  IAA & TAA  |  IBA & TAB  |  ICA & TAC  |  IDA & TAD  |  BAA  ; 
 NCA <=  FCA & ECA  ; 
 OBA <=  FCA & ECA  ; 
 baa <=  aca  |  jaa  ; 
 bag <=  acg  |  jaa  ; 
 ODA <=  LAA & TBA  |  LAB & TBA  |  LAC & TBA  |  LAD & TBA  ; 
 OEA <=  LAA & TBA  |  LAB & TBA  |  LAC & TBA  |  LAD & TBA  ; 
 NDA <=  FDA & EDA  ; 
 OBI <=  FDA & EDA  ; 
 OPF <= HKD ; 
 GAD <= IFD ; 
 GAA <= IFA ; 
 GAB <= IFB ; 
 GAC <= IFC ; 
 ofa <=  aag  |  tca  ; 
 oga <=  aag  |  tcb  ; 
 oia <=  aag  |  tcd  ; 
 oha <=  aag  |  tcc  ; 
 acg <= abg ; 
 aba <= aaa ; 
 aca <= aba ; 
 abg <= aag ; 
 oja <=  haa  |  tea  ; 
 oka <=  haa  |  teb  ; 
 ola <=  haa  |  tec  ; 
 oma <=  haa  |  ted  ; 
 HKD <= HID ; 
 HKA <= HIA ; 
 HKB <= HIB ; 
 HKC <= HIC ; 
 OPC <= HKA ; 
 OPD <= HKB ; 
 OPE <= HKC ; 
 ona <= ija ; 
 onb <= ijb ; 
 onc <= ijc ; 
 DBC <= DBC & tdc |  CAC & TDC ; 
 DBB <= DBB & tdc |  CAB & TDC ; 
 DBA <= DBA & tdc |  CAA & TDC ; 
 HAC <=  RAC & TDA  |  RBC & TDB  |  RCC & TDC  ; 
 HAD <=  RAD & TDA  |  RBD & TDB  |  RCD & TDC  ; 
 wab <= qcb ; 
 tdc <= qcb ; 
 cab <=  cab & kab  |  CAB & KAB  |  JCA  |  TNA  ; 
 cae <=  cab & kab  |  CAB & KAB  |  JCA  |  TNA  ; 
 DKA <=  DKA & thc  |  CCE & THC  ; 
 DKB <=  DKB & thc  |  CCF & THC  ; 
 DHA <=  DHA & tgc  |  CCA & TGC  ; 
 DHB <=  DHB & tgc  |  CCB & TGC  ; 
 DHC <=  DHC & tgc  |  CCC & TGC  ; 
 DHD <=  DHD & tgc  |  CCD & TGC  ; 
 HEC <=  RGC & TGA  |  RHC & TGB  |  RIC & TGC  ; 
 HED <=  RGD & TGA  |  RHD & TGB  |  RID & TGC  ; 
 ccj <= ccf ; 
 thc <= qeb ; 
 wah <= qeb ; 
 tgc <= qeb ; 
 wak <= qeb ; 
 HEG <=  RGG & TGA  |  RHG & TGB  |  RIG & TGC  ; 
 HEH <=  RGH & TGA  |  RHH & TGB  |  RIH & TGC  ; 
 DKC <=  DKC & thc  |  CCG & THC  ; 
 DKD <=  DKD & thc  |  CCH & THC  ; 
 HFC <=  RJC & THA  |  RKC & THB  |  RLC & THC  ; 
 HFD <=  RJD & THA  |  RKD & THB  |  RLD & THC  ; 
 ccb <=  ccb & kcb  |  CCB & KCB  |  JCC  |  TNC  ; 
 ccf <=  ccb & kcb  |  CCB & KCB  |  JCC  |  TNC  ; 
 HFG <=  RJG & THA  |  RKG & THB  |  RLG & THC  ; 
 HFH <=  RJH & THA  |  RKH & THB  |  RLH & THC  ; 
 pab <=  pab & nab  |  FEB  |  TMA  ; 
 pbb <=  pbb & nbb  |  FFB  |  TMB  ; 
 pcb <=  pcb & ncb  |  FGB  |  TMC  ; 
 pdb <=  pdb & ndb  |  FHB  |  TMD  ; 
 GEH <= GAH ; 
 GEE <= GAE ; 
 GEF <= GAF ; 
 GEG <= GAG ; 
 HIH <= HEH ; 
 HIE <= HEE ; 
 HIF <= HEF ; 
 HIG <= HEG ; 
 NAB <=  FAB & EAB  ; 
 OAB <=  FAB & EAB  ; 
 adb <= acb ; 
 adh <= ach ; 
 AAH <=  IAH & TAE  |  IBH & TAF  |  ICH & TAG  |  IDH & TAH  |  BAH  ; 
 NBB <=  FBB & EBB  ; 
 OAJ <=  FBB & EBB  ; 
 NCB <=  FCB & ECB  ; 
 OBB <=  FCB & ECB  ; 
 ach <= abh ; 
 abb <= aab ; 
 acb <= abb ; 
 abh <= aah ; 
 bab <=  acb  |  jaa  ; 
 bah <=  ach  |  jaa  ; 
 ODB <=  LAA & TBB  |  LAB & TBB  |  LAC & TBB  |  LAD & TBB  ; 
 OEB <=  LAA & TBB  |  LAB & TBB  |  LAC & TBB  |  LAD & TBB  ; 
 NDB <=  FDB & EDB  ; 
 OBJ <=  FDB & EDB  ; 
 GAH <= IEC ; 
 GAE <= IFE ; 
 GAF <= IEA ; 
 GAG <= IEB ; 
 ofb <=  aah  |  tca  ; 
 ogb <=  aah  |  tcb  ; 
 ohb <=  aah  |  tcc  ; 
 oib <=  aah  |  tcd  ; 
 ojb <=  hab  |  tea  ; 
 okb <=  hab  |  teb  ; 
 olb <=  hab  |  tec  ; 
 omb <=  hab  |  ted  ; 
 HKH <= HIH ; 
 HKE <= HIE ; 
 HKF <= HIF ; 
 HKG <= HIG ; 
 AAB <=  IAB & TAA  |  IBB & TAB  |  ICB & TAC  |  IDB & TAD  |  BAB  ; 
 OPJ <= HKH ; 
 OPG <= HKE ; 
 OPH <= HKF ; 
 OPI <= HKG ; 
 ond <= ijd ; 
 one <= ije ; 
 onf <= ijf ; 
 DCC <= DCC & tda |  CAC & TDA ; 
 DCB <= DCB & tda |  CAB & TDA ; 
 DCA <= DCA & tda |  CAA & TDA ; 
 QCB <= QCA ; 
 QCC <= QCB ; 
 wac <= qcc ; 
 tda <= qcc ; 
 QCA <=  qcb & qca & tna  ; 
 QCD <=  qcb & qca & tna  ; 
 cac <=  cac & kac  |  CAC & KAC  |  JCA  |  TNA  ; 
 caf <=  cac & kac  |  CAC & KAC  |  JCA  |  TNA  ; 
 DIA <=  DIA & tga  |  CCA & TGA  ; 
 DIB <=  DIB & tga  |  CCB & TGA  ; 
 DIC <=  DIC & tga  |  CCC & TGA  ; 
 DID <=  DID & tga  |  CCD & TGA  ; 
 cck <= ccg ; 
 tha <= qec ; 
 wai <= qec ; 
 tga <= qec ; 
 wal <= qec ; 
 DLA <=  DLA & tha  |  CCE & THA  ; 
 DLB <=  DLB & tha  |  CCF & THA  ; 
 DLC <=  DLC & tha  |  CCG & THA  ; 
 DLD <=  DLD & tha  |  CCH & THA  ; 
 ccc <=  ccc & kcc  |  CCC & KCC  |  JCC  |  TNC  ; 
 ccg <=  ccc & kcc  |  CCC & KCC  |  JCC  |  TNC  ; 
 AED <= JBD ; 
 AEA <= JBA ; 
 AEB <= JBB ; 
 AEC <= JBC ; 
 pac <=  pac & nac  |  FEC  |  TMA  ; 
 AEE <= JBE ; 
 AEF <= JBF ; 
 pbc <=  pbc & nbc  |  FFC  |  TNB  ; 
 pcc <=  pcc & ncc  |  FGC  |  TMC  ; 
 pdc <=  pdc & ndc  |  FHC  |  TMD  ; 
 GFD <= GBD ; 
 GFA <= GBA ; 
 GFB <= GBB ; 
 GFC <= GBC ; 
 HIL <= HFD ; 
 HII <= HFA ; 
 HIJ <= HFB ; 
 HIK <= HFC ; 
 NAC <=  FAC & EAC  ; 
 OAC <=  FAC & EAC  ; 
 adc <= acc ; 
 adi <= aci ; 
 AAI <=  IAI & TAE  |  IBI & TAF  |  ICI & TAG  |  IDI & TAH  |  BAI  ; 
 NBC <=  FBC & EBC  ; 
 OAK <=  FBC & EBC  ; 
 AAC <=  IAC & TAA  |  IBC & TAB  |  ICC & TAC  |  IDC & TAD  |  BAC  ; 
 NCC <=  FCC & ECC  ; 
 OBC <=  FCC & ECC  ; 
 aci <= abi ; 
 acc <= abc ; 
 abi <= aai ; 
 bac <=  acc  |  jaa  ; 
 bai <=  aci  |  jaa  ; 
 ODC <=  LAA & TBC  |  LAB & TBC  |  LAC & TBC  |  LAD & TBC  ; 
 OEC <=  LAA & TBC  |  LAB & TBC  |  LAC & TBC  |  LAD & TBC  ; 
 NDC <=  FDC & EDC  ; 
 OBK <=  FDC & EDC  ; 
 GBD <= IEG ; 
 GBA <= IED ; 
 GBB <= IEE ; 
 GBC <= IEF ; 
 ofc <=  aai  |  tca  ; 
 ogc <=  aai  |  tcb  ; 
 ohc <=  aai  |  tcc  ; 
 oic <=  aai  |  tcd  ; 
 ojc <=  hac  |  tea  ; 
 okc <=  hac  |  teb  ; 
 olc <=  hac  |  tec  ; 
 omc <=  hac  |  ted  ; 
 HKL <= HIL ; 
 HKI <= HII ; 
 HKJ <= HIJ ; 
 HKK <= HIK ; 
 OPN <= HKL ; 
 OPK <= HKI ; 
 OPL <= HKJ ; 
 OPM <= HKK ; 
 ong <= ijg ; 
 onh <= ijh ; 
 oni <= iji ; 
 ccd <=  ccd & kcd  |  CCD & KCD  |  JCC  |  TNC  ; 
 ccl <= cch ; 
 QEA <=  qeb & qea & tnc  ; 
 QED <=  qeb & qea & tnc  ; 
 QEB <= QEA ; 
 QEC <= QEB ; 
 cch <=  ccd & kcd  |  CCD & KCD  |  JCC  |  TNC  ; 
 pad <=  pad & nad  |  FED  |  TMA  ; 
 GFE <= GBE ; 
 pbd <=  pbd & nbd  |  FFD  |  TMB  ; 
 pcd <=  pcd & ncd  |  FGD  |  TMC  ; 
 pdd <=  pdd & ndd  |  FHD  |  TMD  ; 
 HIP <= HFH ; 
 HIM <= HFE ; 
 HIN <= HFF ; 
 HIO <= HFG ; 
 GFH <= GBH ; 
 GFF <= GBF ; 
 GFG <= GBG ; 
 NAD <=  FAD & EAD  ; 
 OAD <=  FAD & EAD  ; 
 add <= acd ; 
 adj <= acj ; 
 AAJ <=  IAJ & TAE  |  IBJ & TAF  |  ICJ & TAG  |  IDJ & TAH  |  BAJ  ; 
 AAM <=  IAJ & TAE  |  IBJ & TAF  |  ICJ & TAG  |  IDJ & TAH  |  BAJ  ; 
 NBD <=  FBD & EBD  ; 
 OAL <=  FBD & EBD  ; 
 qba <=  laa & lab & lac & lad  ; 
 AAD <=  IAD & TAA  |  IBD & TAB  |  ICD & TAC  |  IDD & TAD  |  BAD  ; 
 NCD <=  FCD & ECD  ; 
 OBD <=  FCD & ECD  ; 
 acj <= abj ; 
 abd <= aad ; 
 acd <= abd ; 
 abj <= aaj ; 
 bad <=  acd  |  jaa  ; 
 baj <=  acj  |  jaa  ; 
 ODD <=  LAA & TBD  |  LAB & TBD  |  LAC & TBD  |  LAD & TBD  ; 
 OED <=  LAA & TBD  |  LAB & TBD  |  LAC & TBD  |  LAD & TBD  ; 
 NDD <=  FDD & EDD  ; 
 OBL <=  FDD & EDD  ; 
 GBH <= IEK ; 
 GBE <= IEH ; 
 GBF <= IEI ; 
 GBG <= IEJ ; 
 ofd <=  aaj  |  tca  ; 
 ogd <=  aaj  |  tcb  ; 
 ohd <=  aaj  |  tcc  ; 
 oid <=  aaj  |  tcd  ; 
 ojd <=  had  |  tea  ; 
 okd <=  had  |  teb  ; 
 old <=  had  |  tec  ; 
 omd <=  had  |  ted  ; 
 HKP <= HIP ; 
 HKM <= HIM ; 
 HKN <= HIN ; 
 HKO <= HIO ; 
 OQB <= HKP ; 
 OPO <= HKM ; 
 OPP <= HKN ; 
 OQA <= HKO ; 
 onj <= ijj ; 
 onk <= ijk ; 
 DDA <=  DDA & tfb  |  CBA & TFB  ; 
 DDB <=  DDB & tfb  |  CBB & TFB  ; 
 DDC <=  DDC & tfb  |  CBC & TFB  ; 
 DDD <=  DDD & tfb  |  CBD & TFB  ; 
 HBA <=  RDA & TFA  |  REA & TFB  |  RFA & TFC  ; 
 HBB <=  RDB & TFA  |  REB & TFB  |  RFB & TFC  ; 
 wad <= qda ; 
 tfb <= qda ; 
 cba <=  cba & kba  |  CBA & KBA  |  JCB  |  TMB  ; 
 cbe <=  cba & kba  |  CBA & KBA  |  JCB  |  TMB  ; 
 HBE <=  RDE & TFA  |  REE & TFB  |  RFE & TFC  ; 
 HBF <=  RDF & TFA  |  REFF  & TFB  |  RFF & TFC  ; 
 HHB <=  RPB & TJA  |  RQB & TJB  |  RRB & TJC  ; 
 DMC <=  DMC & tib  |  CCC & TIB  ; 
 DMD <=  DMD & tib  |  CCD & TIB  ; 
 HGA <=  RMA & TIA  |  RNA & TIB  |  ROA & TIC  ; 
 HGB <=  RMB & TIA  |  RNB & TIB  |  ROB & TIC  ; 
 tjb <= qea ; 
 wam <= qea ; 
 tib <= qea ; 
 wap <= qea ; 
 HGE <=  RME & TIA  |  RNE & TIB  |  ROE & TIC  ; 
 HGF <=  RMF & TIA  |  RNF & TIB  |  ROF & TIC  ; 
 DPA <=  DPA & tjb  |  CCE & TJB  ; 
 DPB <=  DPB & tjb  |  CCF & TJB  ; 
 DPC <=  DPC & tjb  |  CCG & TJB  ; 
 DPD <=  DPD & tjb  |  CCH & TJB  ; 
 HHA <=  RPA & TJA  |  RQA & TJB  |  RRA & TJC  ; 
 DMA <=  DMA & tib  |  CCA & TIB  ; 
 DMB <=  DMB & tib  |  CCB & TIB  ; 
 HHE <=  RPE & TJA  |  RQE & TJB  |  RRE & TJC  ; 
 pae <=  pae & nae  |  FEE  |  TMA  ; 
 pbe <=  pbe & nbe  |  FFE  |  TMB  ; 
 pce <=  pce & nce  |  FGE  |  TMC  ; 
 pde <=  pde & nde  |  FHE  |  TMD  ; 
 GGD <= GCD ; 
 GGA <= GCA ; 
 GGB <= GCB ; 
 GGC <= GCC ; 
 HJD <= HGD ; 
 HJA <= HGA ; 
 HJB <= HGB ; 
 HJC <= HGC ; 
 HCF <= HBF ; 
 HCA <= HBA ; 
 HCB <= HBB ; 
 HCE <= HBE ; 
 HDF <= HCF ; 
 HDA <= HCA ; 
 HDB <= HCB ; 
 HDE <= HCE ; 
 NAE <=  FAE & EAE  ; 
 OAE <=  FAE & EAE  ; 
 ade <= ace ; 
 adk <= ack ; 
 AAK <=  IAK & TAE  |  IBK & TAF  |  ICK & TAG  |  IDK & TAH  |  BAK  ; 
 NBE <=  FBE & EBE  ; 
 OAM <=  FBE & EBE  ; 
 qbb <=  lae & laf & lag & lah  ; 
 AAE <=  IAE & TAA  |  IBE & TAB  |  ICE & TAC  |  IDE & TAD  |  BAE  ; 
 NCE <=  FCE & ECE  ; 
 OBE <=  FCE & ECE  ; 
 ack <= abk ; 
 abe <= aae ; 
 ace <= abe ; 
 abk <= aak ; 
 bae <=  ace  |  jaa  ; 
 bak <=  ack  |  jaa  ; 
 ODE <=  LAE & TBA  |  LAF & TBA  |  LAG & TBA  |  LAH & TBA  |  JME  ; 
 OEE <=  LAE & TBA  |  LAF & TBA  |  LAG & TBA  |  LAH & TBA  |  JME  ; 
 NDE <=  FDE & EDE  ; 
 OBM <=  FDE & EDE  ; 
 GCD <= IEO ; 
 GCA <= IEL ; 
 GCB <= IEM ; 
 GCC <= IEN ; 
 onl <= ijl ; 
 onm <= ijm ; 
 onn <= ijn ; 
 oje <=  hae  |  tea  ; 
 oke <=  hae  |  teb  ; 
 ole <=  hae  |  tec  ; 
 ome <=  hae  |  ted  ; 
 HLD <= HJD ; 
 HLA <= HJA ; 
 HLB <= HJB ; 
 HLC <= HJC ; 
 OQF <= HLD ; 
 OQC <= HLA ; 
 OQD <= HLB ; 
 OQE <= HLC ; 
 ono <= ijo ; 
 onp <= ijp ; 
 DEA <=  DEA & tfc  |  CBA & TFC  ; 
 DEB <=  DEB & tfc  |  CBB & TFC  ; 
 DEC <=  DEC & tfc  |  CBC & TFC  ; 
 DED <=  DED & tfc  |  CBD & TFC  ; 
 HBC <=  RDC & TFA  |  REC & TFB  |  RFC & TFC  ; 
 HBD <=  RDD & TFA  |  RED & TFB  |  RFD & TFC  ; 
 wae <= qdb ; 
 tfc <= qdb ; 
 cbb <=  cbb & kbb  |  CBB & KBB  |  JCB  |  TMB  ; 
 cbf <=  cbb & kbb  |  CBB & KBB  |  JCB  |  TMB  ; 
 DQB <=  DQB & tjc  |  CCF & TJC  ; 
 DNA <=  DNA & tic  |  CCA & TIC  ; 
 DNB <=  DNB & tic  |  CCB & TIC  ; 
 DNC <=  DNC & tic  |  CCC & TIC  ; 
 DND <=  DND & tic  |  CCD & TIC  ; 
 HGC <=  RMC & TIA  |  RNC & TIB  |  ROC & TIC  ; 
 HGD <=  RMD & TIA  |  RND & TIB  |  ROD & TIC  ; 
 tjc <= qeb ; 
 wan <= qeb ; 
 tic <= qeb ; 
 waq <= qeb ; 
 HGG <=  RMG & TIA  |  RNG & TIB  |  ROG & TIC  ; 
 HGH <=  RMH & TIA  |  RNH & TIB  |  ROH & TIC  ; 
 DQA <=  DQA & tjc  |  CCE & TJC  ; 
 DQC <=  DQC & tjc  |  CCG & TJC  ; 
 DQD <=  DQD & tjc  |  CCH & TJC  ; 
 HHC <=  RPC & TJA  |  RQC & TJB  |  RRC & TJC  ; 
 HHD <=  RPD & TJA  |  RQD & TJB  |  RRD & TJC  ; 
 paf <=  paf & naf  |  FEF  |  TMA  ; 
 pbf <=  pbf & nbf  |  FFF  |  TMB  ; 
 pcf <=  pcf & ncf  |  FGF  |  TMC  ; 
 pdf <=  pdf & ndf  |  FHF  |  TMD  ; 
 GGH <= GCH ; 
 GGE <= GCE ; 
 GGF <= GCF ; 
 GGG <= GCG ; 
 HJH <= HGH ; 
 HJE <= HGE ; 
 HJF <= HGF ; 
 HJG <= HGG ; 
 HCC <= HBC ; 
 HCD <= HBD ; 
 HDC <= HCC ; 
 HDD <= HCD ; 
 NAF <=  FAF & EAF  ; 
 OAF <=  FAF & EAF  ; 
 adf <= acf ; 
 adl <= acl ; 
 abl <= aal ; 
 AAL <=  IAL & TAE  |  IBL & TAF  |  ICL & TAG  |  IDL & TAH  |  BAL  ; 
 NBF <=  FBF & EBF  ; 
 OAN <=  FBF & EBF  ; 
 NCF <=  FCF & ECF  ; 
 OBF <=  FCF & ECF  ; 
 bal <=  acl  |  jaa  ; 
 baf <=  acf  |  jaa  ; 
 ODF <=  LAE & TBB  |  LAF & TBB  |  LAG & TBB  |  LAH & TBB  |  JME  ; 
 OEF <=  LAE & TBB  |  LAF & TBB  |  LAG & TBB  |  LAH & TBB  |  JME  ; 
 NDF <=  FDF & EDF  ; 
 OBN <=  FDF & EDF  ; 
 GCH <= IES ; 
 GCE <= IEP ; 
 GCF <= IEQ ; 
 GCG <= IER ; 
 ofe <=  aal  |  tca  ; 
 oge <=  aal  |  tcb  ; 
 ohe <=  aal  |  tcc  ; 
 oie <=  aal  |  tcd  ; 
 acl <= abl ; 
 abc <= aac ; 
 abf <= aaf ; 
 acf <= abf ; 
 ojf <=  haf  |  tea  ; 
 okf <=  haf  |  teb  ; 
 olf <=  haf  |  tec  ; 
 omf <=  haf  |  ted  ; 
 HLH <= HJH ; 
 HLE <= HJE ; 
 HLF <= HJF ; 
 HLG <= HJG ; 
 AAF <=  IAF & TAA  |  IBF & TAB  |  ICF & TAC  |  IDF & TAD  |  BAF  ; 
 OQJ <= HLH ; 
 OQG <= HLE ; 
 OQH <= HLF ; 
 OQI <= HLG ; 
 ooa <= ika ; 
 oob <= ikb ; 
 ooc <= ikc ; 
 DFA <=  DFA & tfa  |  CBA & TFA  ; 
 DFB <=  DFB & tfa  |  CBB & TFA  ; 
 DFC <=  DFC & tfa  |  CBC & TFA  ; 
 DFD <=  DFD & tfa  |  CBD & TFA  ; 
 QDB <= QDA ; 
 QDC <= QDB ; 
 waf <= qdc ; 
 tfa <= qdc ; 
 QDA <=  qdb & qda & tnb  ; 
 QDD <=  qdb & qda & tnb  ; 
 cbc <=  cbc & kbc  |  CBC & KBC  |  JCB  |  TNB  ; 
 cbg <=  cbc & kbc  |  CBC & KBC  |  JCB  |  TNB  ; 
 DOA <=  DOA & tia  |  CCA & TIA  ; 
 DOB <=  DOB & tia  |  CCB & TIA  ; 
 DOC <=  DOC & tia  |  CCC & TIA  ; 
 DOD <=  DOD & tia  |  CCD & TIA  ; 
 tja <= qec ; 
 wao <= qec ; 
 tia <= qec ; 
 war <= qec ; 
 DRB <=  DRB & tja  |  CCF & TJA  ; 
 DRA <=  DRA & tja  |  CCE & TJA  ; 
 DRC <=  DRC & tja  |  CCG & TJA  ; 
 DRD <=  DRD & tja  |  CCH & TJA  ; 
 AEJ <= JBJ ; 
 AEG <= JBG ; 
 AEH <= JBH ; 
 AEI <= JBI ; 
 pag <=  pag & nag  |  FEG  |  TMA  ; 
 AEK <= JBK ; 
 AEL <= JBL ; 
 pbg <=  pbg & nbg  |  FFG  |  TMB  ; 
 pcg <=  pcg & ncg  |  FGG  |  TMC  ; 
 pdg <=  pdg & ndg  |  FHG  |  TMD  ; 
 GHD <= GDD ; 
 GHA <= GDA ; 
 GHB <= GDB ; 
 GHC <= GDC ; 
 HJL <= HHD ; 
 HJI <= HHA ; 
 HJJ <= HHB ; 
 HJK <= HHC ; 
 NAG <=  FAG & EAG  ; 
 OAG <=  FAG & EAG  ; 
 QBC <= JAA ; 
 QBD <= JAA ; 
 TAD <= jab & QAC ; 
 TAA <= jab & QAA ; 
 TAB <= jab & QAA ; 
 TAC <= jab & QAB ; 
 NBG <=  FBG & EBG  ; 
 OAO <=  FBG & EBG  ; 
 TAH <= jab & QAC ; 
 TAE <= jab & QAD ; 
 TAF <= jab & QAA ; 
 NCG <=  FCG & ECG  ; 
 OBG <=  FCG & ECG  ; 
 ODG <=  LAE & TBC  |  LAF & TBC  |  LAG & TBC  |  LAH & TBC  |  JME  ; 
 OEG <=  LAE & TBC  |  LAF & TBC  |  LAG & TBC  |  LAH & TBC  |  JME  ; 
 NDG <=  FDG & EDG  ; 
 OBO <=  FDG & EDG  ; 
 OQM <= HLK ; 
 GDD <= IEW ; 
 GDA <= IET ; 
 GDB <= IEU ; 
 GDC <= IEV ; 
 ood <= ikd ; 
 ooe <= ike ; 
 oof <= ikf ; 
 oog <= ikg ; 
 ooh <= ikh ; 
 ooi <= iki ; 
 HLL <= HJL ; 
 HLI <= HJI ; 
 HLJ <= HJJ ; 
 HLK <= HJK ; 
 TAG <= jab & QAB ; 
 OQN <= HLL ; 
 OQK <= HLI ; 
 OQL <= HLJ ; 
 ooj <= ikj ; 
 ook <= ikk ; 
 cbd <=  cbd & kbd  |  CBD & KBD  |  JCB  |  TNB  ; 
 cbh <=  cbd & kbd  |  CBD & KBD  |  JCB  |  TNB  ; 
 pah <=  pah & nah  |  FEH  |  TMA  ; 
 GHE <= GDE ; 
 pbh <=  pbh & nbh  |  FFH  |  TMB  ; 
 pch <=  pch & nch  |  FGH  |  TMC  ; 
 pdh <=  pdh & ndh  |  FHH  |  TMD  ; 
 HJM <= HHE ; 
 tna <=  igc  ; 
 tnb <=  igc  ; 
 tnc <=  igc  ; 
 TMD <= IGA ; 
 TMA <= IGA ; 
 TMB <= IGA ; 
 TMC <= IGA ; 
 NAH <=  FAH & EAH  ; 
 OAH <=  FAH & EAH  ; 
 qfa <=  qab & qad  ; 
 qfb <=  qac & qad  ; 
 QAD <= QAC ; 
 QAA <= IGB ; 
 QAB <= QAA ; 
 QAC <= QAB ; 
 NBH <=  FBH & EBH  ; 
 OAP <=  FBH & EBH  ; 
 tbd <= qaa ; 
 tba <= qab ; 
 NCH <=  FCH & ECH  ; 
 OBH <=  FCH & ECH  ; 
 tcd <= qad ; 
 tca <= qaa ; 
 tcb <= qab ; 
 tcc <= qac ; 
 ODH <=  LAE & TBD  |  LAF & TBD  |  LAG & TBD  |  LAH & TBD  |  JME  ; 
 OEH <=  LAE & TBD  |  LAF & TBD  |  LAG & TBD  |  LAH & TBD  |  JME  ; 
 NDH <=  FDH & EDH  ; 
 OBP <=  FDH & EDH  ; 
 ted <= qab ; 
 tea <= qac ; 
 teb <= qad ; 
 tec <= qaa ; 
 ool <= ikl ; 
 oom <= ikm ; 
 oon <= ikn ; 
 GDE <=  IEX  ; 
 HLM <= HJM ; 
 tbb <= qac ; 
 tbc <= qad ; 
 OQO <= HLM ; 
 OPA <= QFA ; 
 OPB <= QFB ; 
 ooo <= iko ; 
 oop <= ikp ; 
end
ram_16x4 rinst_0(RAA,RAB,RAC,RAD,AEA,AEB,AEC,AED,ZZI,DAC,DAB,DAA, ZZI, WAA, IZZ); 
ram_16x4 rinst_1(RAE,RAF,RAG,RAH,AEE,AEF,ZZI,ZZI,ZZI,DAC,DAB,DAA, ZZI, WAA, IZZ); 
ram_16x4 rinst_2(RGA,RGB,RGC,RGD,GEA,GEB,GEC,GED,DGD,DGC,DGB,DGA, ZZI, WAG, IZZ); 
ram_16x4 rinst_3(RGE,RGF,RGG,RGH,GEE,GEF,GEG,GEH,DGD,DGC,DGB,DGA, ZZI, WAG, IZZ); 
ram_16x4 rinst_4(RJA,RJB,RJC,RJD,GFA,GFB,GFC,GFD,DKD,DKC,DKB,DKA, ZZI, WAJ, IZZ); 
ram_16x4 rinst_5(RJE,RJF,RJG,RJH,GFE,GFF,GFG,GFH,DKD,DKC,DKB,DKA, ZZI, WAJ, IZZ); 
ram_16x4 rinst_6(RBA,RBB,RBC,RBD,AEA,AEB,AEC,AED,ZZI,DBC,DBB,DBA, ZZI, WAB, IZZ); 
ram_16x4 rinst_7(RBE,RBF,RBG,RBH,AEE,AEF,ZZI,ZZI,ZZI,DBC,DBB,DBA, ZZI, WAB, IZZ); 
ram_16x4 rinst_8(RHA,RHB,RHC,RHD,GEA,GEB,GEC,GED,DHD,DHC,DHB,DHA, ZZI, WAH, IZZ); 
ram_16x4 rinst_9(RHE,RHF,RHG,RHH,GEE,GEF,GEG,GEH,DHD,DHC,DHB,DHA, ZZI, WAH, IZZ); 
ram_16x4 rinst_10(RKA,RKB,RKC,RKD,GFA,GFB,GFC,GFD,DKD,DKC,DKB,DKA, ZZI, WAK, IZZ); 
ram_16x4 rinst_11(RKE,RKF,RKG,RKH,GFE,GFF,GFG,GFH,DKD,DKC,DKB,DKA, ZZI, WAK, IZZ); 
ram_16x4 rinst_12(RCA,RCB,RCC,RCD,AEA,AEB,AEC,AED,ZZI,DCC,DCB,DCA, ZZI, WAC, IZZ); 
ram_16x4 rinst_13(RCE,RCF,RCG,RCH,AEE,AEF,ZZI,ZZI,ZZI,DCC,DCB,DCA, ZZI, WAC, IZZ); 
ram_16x4 rinst_14(RIA,RIB,RIC,RID,GEA,GEB,GEC,GED,DID,DIC,DEB,DIA, ZZI, WAI, IZZ); 
ram_16x4 rinst_15(RIE,RIF,RIG,RIH,GEE,GEF,GEG,GEH,DID,DIC,DIB,DIA, ZZI, WAI, IZZ); 
ram_16x4 rinst_16(RLA,RLB,RLC,RLD,GFA,GFB,GFC,GFD,DLD,DLC,DLB,DLA, ZZI, WAL, IZZ); 
ram_16x4 rinst_17(RLE,RLF,RLG,RLH,GFE,GFF,GFG,GFH,DLD,DLC,DLB,DLA, ZZI, WAL, IZZ); 
ram_16x4 rinst_18(RDA,RDB,RDC,RDD,AEG,AEH,AEI,AEJ,DDD,DDC,DDB,DDA, ZZI, WAD, IZZ); 
ram_16x4 rinst_19(RDE,RDF,RDG,RDH,AEK,AEL,ZZI,ZZI,DDD,DDC,DDB,DDA, ZZI, WAD, IZZ); 
ram_16x4 rinst_20(RMA,RMB,RMC,RMD,GGA,GGB,GGC,GGD,DMD,DMC,DMB,DNA, ZZI, WAM, IZZ); 
ram_16x4 rinst_21(RME,RMF,RMG,RMH,GGE,GGF,GGG,GGH,DMD,DMC,DMB,DNA, ZZI, WAM, IZZ); 
ram_16x4 rinst_22(RPA,RPB,RPC,RPD,GHA,GHB,GHC,GHD,DPD,DPC,DPB,DPA, ZZI, WAP, IZZ); 
ram_16x4 rinst_23(REA,REB,REC,RED,AEG,AEH,AEI,AEJ,DED,DEC,DEB,DEA, ZZI, WAE, IZZ); 
ram_16x4 rinst_24(REE,REFF ,REG,REH,AEK,AEL,ZZI,ZZI,DED,DEC,DEB,DEA, ZZI, WAE, IZZ); 
ram_16x4 rinst_25(RNA,RNB,RNC,RND,GGA,GGB,GGC,GGD,DND,DNC,DNB,DNA, ZZI, WAN, IZZ); 
ram_16x4 rinst_26(RNE,RNF,RNG,RNH,GGE,GGF,GGG,GGH,DND,DNC,DNB,DNA, ZZI, WAN, IZZ); 
ram_16x4 rinst_27(RQA,RQB,RQC,RQD,GHA,GHB,GHC,GHD,DQD,DQC,DQB,DQA, ZZI, WAQ, IZZ); 
ram_16x4 rinst_28(RFA,RFB,RFC,RFD,AEG,AEH,AEI,AEJ,DFD,DFC,DFB,DFA, ZZI, WAF, IZZ); 
ram_16x4 rinst_29(RFE,RFF,RFG,RFH,AEK,AEL,ZZI,ZZI,DFD,DFC,DFB,DFA, ZZI, WAF, IZZ); 
ram_16x4 rinst_30(ROA,ROB,ROC,ROD,GGA,GGB,GGC,GGD,DOD,DOC,DOB,DOA, ZZI, WAO, IZZ); 
ram_16x4 rinst_31(ROE,ROF,ROG,ROH,GGE,GGF,GGG,GGH,DOD,DOC,DOB,DOA, ZZI, WAO, IZZ); 
ram_16x4 rinst_32(RRA,RRB,RRC,RRD,GHA,GHB,GHC,GHD, DRD,DRC,DRB,DRA, ZZI, WAR, IZZ); 
endmodule;
