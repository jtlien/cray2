module ra( IZZ,
 IAA, 
 IAB, 
 IAC, 
 IAD, 
 IAE, 
 IAF, 
 IAG, 
 IAH, 
 IAI, 
 IAJ, 
 IAK, 
 IAL, 
 IAM, 
 IAN, 
 IAO, 
 IAP, 
 ICA, 
 ICB, 
 ICC, 
 ICD, 
 ICE, 
 ICF, 
 ICG, 
 ICH, 
 ICI, 
 ICJ, 
 ICK, 
 ICL, 
 ICM, 
 ICN, 
 ICO, 
 ICP, 
 IGA, 
 IJA, 
 IKA, 
 ILA, 
 ILB, 
 ILC, 
 ILD, 
 ILE, 
 ILF, 
 ILG, 
 ILH, 
 ILI, 
 IPA, 
 IPB, 
 IQA, 
 IQB, 
 IQC, 
 IRA, 
 IRB, 
 ISA, 
 OAA, 
 OAB, 
 OAC, 
 OAD, 
 OAE, 
 OAF, 
 OAG, 
 OAH, 
 OAI, 
 OAJ, 
 OAK, 
 OAL, 
 OAM, 
 OAN, 
 OAO, 
 OAP, 
 OAQ, 
 OAR, 
 OAS, 
 OAT, 
 OAU, 
 OAV, 
 OAW, 
 OAX, 
 OAY, 
 OAZ, 
 OBA, 
 OBB, 
 OBC, 
 OBD, 
 OBE, 
 OBF, 
 OBG, 
 OBH, 
 OBI, 
 OBJ, 
 OBK, 
 OBL, 
 OBM, 
 OBN, 
 OBO, 
 OBP, 
 OBQ, 
 OBR, 
 OBS, 
 OBT, 
 OBU, 
 OBV, 
 OBW, 
 OBX, 
 OBY, 
 OBZ, 
 OCA, 
 OCB, 
 OCC, 
 OCD, 
 OCE, 
 OCF, 
 OCG, 
 OCH, 
 OCI, 
 OCJ, 
 OCK, 
 OCL, 
 OCM, 
 OCN, 
 OCO, 
 OCP, 
 OCQ, 
 OCR, 
 OCS, 
 OCT, 
 OCU, 
 OCV, 
 OCW, 
 OCX, 
 OCY, 
 OCZ, 
 ODA, 
 ODB, 
 ODC, 
 ODD, 
 ODE, 
 ODF, 
 ODG, 
 ODH, 
 ODI, 
 ODJ, 
 ODK, 
 ODL, 
 ODM, 
 ODN, 
 ODO, 
 ODP, 
 ODQ, 
 ODR, 
 ODS, 
 ODT, 
 ODU, 
 ODV, 
 ODW, 
 ODX, 
 ODY, 
 ODZ, 
 OEA, 
 OEB, 
 OEC, 
 OED, 
 OEE, 
 OEF, 
 OEG, 
 OEH, 
 OEI, 
 OEJ, 
 OEK, 
 OEL, 
 OEM, 
 OEN, 
 OEO, 
 OEP, 
 OFA, 
 OFB, 
 OFC, 
 OFD, 
 OFE, 
 OFF, 
 OFG, 
 OFH, 
 OFI, 
 OFJ, 
 OFK, 
 OFL, 
 OFM, 
 OFN, 
 OFO, 
 OFP, 
 OGA, 
 OGB, 
 OGC, 
 OGD, 
 OGE, 
 OGF, 
 OGG, 
 OGH, 
 OGI, 
 OGJ, 
 OGK, 
 OGL, 
 OGM, 
 OGN, 
 OGO, 
 OGP, 
 OHA, 
 OHB, 
 OHC, 
 OHD, 
 OHE, 
 OHF, 
 OHG, 
 OHH, 
 OHI, 
 OHJ, 
 OHK, 
 OHL, 
 OHM, 
 OHN, 
 OHO, 
 OHP, 
 OIA, 
 OIB, 
 OIC, 
 OID, 
 OIE, 
 OIF, 
 OIG, 
 OIH, 
 OII, 
 OIJ, 
 OIK, 
 OIL, 
 OIM, 
 OJA, 
 OKA, 
 OKB, 
 OKC, 
 OKD, 
 OKE, 
 OKF, 
 OKG, 
 OLA, 
 OLB, 
 OLC, 
 OLD, 
 OLE, 
 OLF, 
 OLG, 
 OLH, 
 OLI, 
 OMA, 
ONA ); 
    
 input IZZ; 
 input IAA; 
 input IAB; 
 input IAC; 
 input IAD; 
 input IAE; 
 input IAF; 
 input IAG; 
 input IAH; 
 input IAI; 
 input IAJ; 
 input IAK; 
 input IAL; 
 input IAM; 
 input IAN; 
 input IAO; 
 input IAP; 
 input ICA; 
 input ICB; 
 input ICC; 
 input ICD; 
 input ICE; 
 input ICF; 
 input ICG; 
 input ICH; 
 input ICI; 
 input ICJ; 
 input ICK; 
 input ICL; 
 input ICM; 
 input ICN; 
 input ICO; 
 input ICP; 
 input IGA; 
 input IJA; 
 input IKA; 
 input ILA; 
 input ILB; 
 input ILC; 
 input ILD; 
 input ILE; 
 input ILF; 
 input ILG; 
 input ILH; 
 input ILI; 
 input IPA; 
 input IPB; 
 input IQA; 
 input IQB; 
 input IQC; 
 input IRA; 
 input IRB; 
 input ISA; 
 output OAA; 
 output OAB; 
 output OAC; 
 output OAD; 
 output OAE; 
 output OAF; 
 output OAG; 
 output OAH; 
 output OAI; 
 output OAJ; 
 output OAK; 
 output OAL; 
 output OAM; 
 output OAN; 
 output OAO; 
 output OAP; 
 output OAQ; 
 output OAR; 
 output OAS; 
 output OAT; 
 output OAU; 
 output OAV; 
 output OAW; 
 output OAX; 
 output OAY; 
 output OAZ; 
 output OBA; 
 output OBB; 
 output OBC; 
 output OBD; 
 output OBE; 
 output OBF; 
 output OBG; 
 output OBH; 
 output OBI; 
 output OBJ; 
 output OBK; 
 output OBL; 
 output OBM; 
 output OBN; 
 output OBO; 
 output OBP; 
 output OBQ; 
 output OBR; 
 output OBS; 
 output OBT; 
 output OBU; 
 output OBV; 
 output OBW; 
 output OBX; 
 output OBY; 
 output OBZ; 
 output OCA; 
 output OCB; 
 output OCC; 
 output OCD; 
 output OCE; 
 output OCF; 
 output OCG; 
 output OCH; 
 output OCI; 
 output OCJ; 
 output OCK; 
 output OCL; 
 output OCM; 
 output OCN; 
 output OCO; 
 output OCP; 
 output OCQ; 
 output OCR; 
 output OCS; 
 output OCT; 
 output OCU; 
 output OCV; 
 output OCW; 
 output OCX; 
 output OCY; 
 output OCZ; 
 output ODA; 
 output ODB; 
 output ODC; 
 output ODD; 
 output ODE; 
 output ODF; 
 output ODG; 
 output ODH; 
 output ODI; 
 output ODJ; 
 output ODK; 
 output ODL; 
 output ODM; 
 output ODN; 
 output ODO; 
 output ODP; 
 output ODQ; 
 output ODR; 
 output ODS; 
 output ODT; 
 output ODU; 
 output ODV; 
 output ODW; 
 output ODX; 
 output ODY; 
 output ODZ; 
 output OEA; 
 output OEB; 
 output OEC; 
 output OED; 
 output OEE; 
 output OEF; 
 output OEG; 
 output OEH; 
 output OEI; 
 output OEJ; 
 output OEK; 
 output OEL; 
 output OEM; 
 output OEN; 
 output OEO; 
 output OEP; 
 output OFA; 
 output OFB; 
 output OFC; 
 output OFD; 
 output OFE; 
 output OFF; 
 output OFG; 
 output OFH; 
 output OFI; 
 output OFJ; 
 output OFK; 
 output OFL; 
 output OFM; 
 output OFN; 
 output OFO; 
 output OFP; 
 output OGA; 
 output OGB; 
 output OGC; 
 output OGD; 
 output OGE; 
 output OGF; 
 output OGG; 
 output OGH; 
 output OGI; 
 output OGJ; 
 output OGK; 
 output OGL; 
 output OGM; 
 output OGN; 
 output OGO; 
 output OGP; 
 output OHA; 
 output OHB; 
 output OHC; 
 output OHD; 
 output OHE; 
 output OHF; 
 output OHG; 
 output OHH; 
 output OHI; 
 output OHJ; 
 output OHK; 
 output OHL; 
 output OHM; 
 output OHN; 
 output OHO; 
 output OHP; 
 output OIA; 
 output OIB; 
 output OIC; 
 output OID; 
 output OIE; 
 output OIF; 
 output OIG; 
 output OIH; 
 output OII; 
 output OIJ; 
 output OIK; 
 output OIL; 
 output OIM; 
 output OJA; 
 output OKA; 
 output OKB; 
 output OKC; 
 output OKD; 
 output OKE; 
 output OKF; 
 output OKG; 
 output OLA; 
 output OLB; 
 output OLC; 
 output OLD; 
 output OLE; 
 output OLF; 
 output OLG; 
 output OLH; 
 output OLI; 
 output OMA; 
 output ONA; 
  
  
reg  AAA ;
reg  AAB ;
reg  AAC ;
reg  AAD ;
reg  AAE ;
reg  AAF ;
reg  AAG ;
reg  AAH ;
reg  AAI ;
reg  AAJ ;
reg  AAK ;
reg  AAL ;
reg  ABA ;
reg  ABB ;
reg  ABC ;
reg  ABD ;
reg  ABE ;
reg  ABF ;
reg  ABG ;
reg  ABH ;
reg  ABI ;
reg  ABJ ;
reg  ABK ;
reg  ABL ;
reg  ACA ;
reg  ACB ;
reg  ACC ;
reg  ACD ;
reg  ACE ;
reg  ACF ;
reg  ACG ;
reg  ACH ;
reg  ACI ;
reg  ACJ ;
reg  ACK ;
reg  ACL ;
reg  ADB ;
reg  ADC ;
reg  ADD ;
reg  ADE ;
reg  ADF ;
reg  ADG ;
reg  ADH ;
reg  ADI ;
reg  ADJ ;
reg  ADK ;
reg  ADL ;
reg  AEA ;
reg  AEB ;
reg  AEC ;
reg  AED ;
reg  AEE ;
reg  AEF ;
reg  AEG ;
reg  AEH ;
reg  AEI ;
reg  AEJ ;
reg  AEK ;
reg  AEL ;
reg  AFA ;
reg  AFB ;
reg  AFC ;
reg  AFD ;
reg  AFE ;
reg  AFF ;
reg  AFG ;
reg  AFH ;
reg  AFI ;
reg  AFJ ;
reg  AFK ;
reg  AFL ;
reg  agb ;
reg  agc ;
reg  agd ;
reg  age ;
reg  agf ;
reg  agg ;
reg  agh ;
reg  agi ;
reg  agj ;
reg  agk ;
reg  agl ;
reg  aha ;
reg  ahb ;
reg  ahc ;
reg  ahd ;
reg  ahe ;
reg  ahf ;
reg  ahg ;
reg  ahh ;
reg  ahi ;
reg  ahj ;
reg  ahk ;
reg  ahl ;
reg  aia ;
reg  aib ;
reg  aic ;
reg  aid ;
reg  aie ;
reg  aif ;
reg  aig ;
reg  aih ;
reg  aii ;
reg  aij ;
reg  aik ;
reg  ail ;
reg  ajb ;
reg  ajc ;
reg  ajd ;
reg  aje ;
reg  ajf ;
reg  ajg ;
reg  ajh ;
reg  aji ;
reg  ajj ;
reg  ajk ;
reg  ajl ;
reg  aka ;
reg  akb ;
reg  akc ;
reg  akd ;
reg  ake ;
reg  akf ;
reg  akg ;
reg  akh ;
reg  aki ;
reg  akj ;
reg  akk ;
reg  akl ;
reg  ala ;
reg  alb ;
reg  alc ;
reg  ald ;
reg  ale ;
reg  alf ;
reg  alg ;
reg  alh ;
reg  ali ;
reg  alj ;
reg  alk ;
reg  all ;
reg  AMA ;
reg  AMB ;
reg  AMC ;
reg  AMD ;
reg  AME ;
reg  AMF ;
reg  AMG ;
reg  AMH ;
reg  AMI ;
reg  AMJ ;
reg  AMK ;
reg  AML ;
reg  AMM ;
reg  AMN ;
reg  AMO ;
reg  AMP ;
reg  BAK ;
reg  BAL ;
reg  BAM ;
reg  BAN ;
reg  BAO ;
reg  BAP ;
reg  BAQ ;
reg  BAR ;
reg  BAS ;
reg  BAT ;
reg  BAU ;
reg  BAV ;
reg  BAW ;
reg  BAX ;
reg  BAY ;
reg  BAZ ;
reg  bba ;
reg  bbb ;
reg  bbc ;
reg  bbd ;
reg  bbe ;
reg  bbf ;
reg  bbg ;
reg  bbh ;
reg  bbi ;
reg  bbj ;
reg  bbk ;
reg  bbl ;
reg  bbm ;
reg  bbn ;
reg  bbo ;
reg  bbp ;
reg  BCA ;
reg  BCB ;
reg  BCC ;
reg  BCD ;
reg  BCE ;
reg  BCF ;
reg  BCG ;
reg  BCH ;
reg  BCI ;
reg  BCJ ;
reg  BCK ;
reg  BCL ;
reg  BCM ;
reg  BCN ;
reg  BCO ;
reg  BCP ;
reg  BDA ;
reg  BDB ;
reg  BDC ;
reg  BDD ;
reg  BDE ;
reg  BDF ;
reg  BDG ;
reg  BDH ;
reg  BDI ;
reg  BDJ ;
reg  BDK ;
reg  BDL ;
reg  BDM ;
reg  BDN ;
reg  BDO ;
reg  BDP ;
reg  BEA ;
reg  BEB ;
reg  BEC ;
reg  BED ;
reg  BEE ;
reg  BEF ;
reg  BEG ;
reg  BEH ;
reg  BEI ;
reg  BEJ ;
reg  BEK ;
reg  BEL ;
reg  BEM ;
reg  BEN ;
reg  BEO ;
reg  BEP ;
reg  BFA ;
reg  BFB ;
reg  BFC ;
reg  DAA ;
reg  DAB ;
reg  DAC ;
reg  DAD ;
reg  DAE ;
reg  DAF ;
reg  DAG ;
reg  DAH ;
reg  DBA ;
reg  DBB ;
reg  DBC ;
reg  DBD ;
reg  DBE ;
reg  DBF ;
reg  DBG ;
reg  DBH ;
reg  dca ;
reg  dcb ;
reg  dcc ;
reg  dcd ;
reg  dce ;
reg  dcf ;
reg  dcg ;
reg  dch ;
reg  dda ;
reg  ddb ;
reg  ddc ;
reg  ddd ;
reg  dde ;
reg  ddf ;
reg  ddg ;
reg  ddh ;
reg  DIA ;
reg  DIB ;
reg  DIC ;
reg  DID ;
reg  DIE ;
reg  DIF ;
reg  DIG ;
reg  DIH ;
reg  eaa ;
reg  eab ;
reg  eac ;
reg  ead ;
reg  eae ;
reg  eaf ;
reg  eag ;
reg  eah ;
reg  eai ;
reg  eaj ;
reg  eak ;
reg  eal ;
reg  eba ;
reg  ebb ;
reg  ebc ;
reg  ebd ;
reg  ebe ;
reg  ebf ;
reg  ebg ;
reg  ebh ;
reg  ebi ;
reg  ebj ;
reg  ebk ;
reg  ebl ;
reg  eca ;
reg  ecb ;
reg  ecc ;
reg  ecd ;
reg  ece ;
reg  ecf ;
reg  ecg ;
reg  ech ;
reg  eci ;
reg  ecj ;
reg  eck ;
reg  ecl ;
reg  fba ;
reg  fbb ;
reg  fca ;
reg  OAA ;
reg  OAB ;
reg  OAC ;
reg  OAD ;
reg  OAE ;
reg  OAF ;
reg  OAG ;
reg  OAH ;
reg  OAI ;
reg  OAJ ;
reg  OAK ;
reg  OAL ;
reg  OAM ;
reg  OAN ;
reg  OAO ;
reg  OAP ;
reg  OAQ ;
reg  OAR ;
reg  OAS ;
reg  OAT ;
reg  OAU ;
reg  OAV ;
reg  OAW ;
reg  OAX ;
reg  OAY ;
reg  OAZ ;
reg  OBA ;
reg  OBB ;
reg  OBC ;
reg  OBD ;
reg  OBE ;
reg  OBF ;
reg  OBG ;
reg  OBH ;
reg  OBI ;
reg  OBJ ;
reg  OBK ;
reg  OBL ;
reg  OBM ;
reg  OBN ;
reg  OBO ;
reg  OBP ;
reg  OBQ ;
reg  OBR ;
reg  OBS ;
reg  OBT ;
reg  OBU ;
reg  OBV ;
reg  OBW ;
reg  OBX ;
reg  OBY ;
reg  OBZ ;
reg  OCA ;
reg  OCB ;
reg  OCC ;
reg  OCD ;
reg  OCE ;
reg  OCF ;
reg  OCG ;
reg  OCH ;
reg  OCI ;
reg  OCJ ;
reg  OCK ;
reg  OCL ;
reg  OCM ;
reg  OCN ;
reg  OCO ;
reg  OCP ;
reg  OCQ ;
reg  OCR ;
reg  OCS ;
reg  OCT ;
reg  OCU ;
reg  OCV ;
reg  OCW ;
reg  OCX ;
reg  OCY ;
reg  OCZ ;
reg  ODA ;
reg  ODB ;
reg  ODC ;
reg  ODD ;
reg  ODE ;
reg  ODF ;
reg  ODG ;
reg  ODH ;
reg  ODI ;
reg  ODJ ;
reg  ODK ;
reg  ODL ;
reg  ODM ;
reg  ODN ;
reg  ODO ;
reg  ODP ;
reg  ODQ ;
reg  ODR ;
reg  ODS ;
reg  ODT ;
reg  ODU ;
reg  ODV ;
reg  ODW ;
reg  ODX ;
reg  ODY ;
reg  ODZ ;
reg  OEA ;
reg  OEB ;
reg  OEC ;
reg  OED ;
reg  OEE ;
reg  OEF ;
reg  OEG ;
reg  OEH ;
reg  OEI ;
reg  OEJ ;
reg  OEK ;
reg  OEL ;
reg  OEM ;
reg  OEN ;
reg  OEO ;
reg  OEP ;
reg  OFA ;
reg  OFB ;
reg  OFC ;
reg  OFD ;
reg  OFE ;
reg  OFF ;
reg  OFG ;
reg  OFH ;
reg  OFI ;
reg  OFJ ;
reg  OFK ;
reg  OFL ;
reg  OFM ;
reg  OFN ;
reg  OFO ;
reg  OFP ;
reg  oga ;
reg  ogb ;
reg  ogc ;
reg  ogd ;
reg  oge ;
reg  ogf ;
reg  ogg ;
reg  ogh ;
reg  ogi ;
reg  ogj ;
reg  ogk ;
reg  ogl ;
reg  ogm ;
reg  ogn ;
reg  ogo ;
reg  ogp ;
reg  oha ;
reg  ohb ;
reg  ohc ;
reg  ohd ;
reg  ohe ;
reg  ohf ;
reg  ohg ;
reg  ohh ;
reg  ohi ;
reg  ohj ;
reg  ohk ;
reg  ohl ;
reg  ohm ;
reg  ohn ;
reg  oho ;
reg  ohp ;
reg  OIA ;
reg  OIB ;
reg  OIC ;
reg  OID ;
reg  OIE ;
reg  OIF ;
reg  OIG ;
reg  OIH ;
reg  OII ;
reg  OIJ ;
reg  OIK ;
reg  OIL ;
reg  OIM ;
reg  oja ;
reg  OKA ;
reg  OKB ;
reg  OKC ;
reg  OKD ;
reg  OKE ;
reg  OKF ;
reg  OKG ;
reg  OLA ;
reg  OLB ;
reg  OLC ;
reg  OLD ;
reg  OLE ;
reg  OLF ;
reg  OLG ;
reg  OLH ;
reg  OLI ;
reg  OMA ;
reg  ONA ;
reg  paa ;
reg  pab ;
reg  pac ;
reg  pad ;
reg  pae ;
reg  paf ;
reg  pag ;
reg  pah ;
reg  pai ;
reg  paj ;
reg  pak ;
reg  pal ;
reg  pam ;
reg  pan ;
reg  pao ;
reg  pap ;
reg  paq ;
reg  par ;
reg  pas ;
reg  pat ;
reg  pba ;
reg  pbb ;
reg  pbc ;
reg  pbd ;
reg  pbe ;
reg  pbf ;
reg  pbg ;
reg  pbh ;
reg  pbi ;
reg  pbj ;
reg  pbk ;
reg  pbl ;
reg  pbm ;
reg  pbn ;
reg  pbo ;
reg  pbp ;
reg  pbq ;
reg  pbr ;
reg  pbs ;
reg  pbt ;
reg  PCA ;
reg  PCB ;
reg  PCC ;
reg  PCD ;
reg  PCE ;
reg  PCF ;
reg  PCG ;
reg  PCH ;
reg  PCI ;
reg  PCJ ;
reg  PCK ;
reg  PCL ;
reg  PCM ;
reg  PCN ;
reg  PDA ;
reg  PDB ;
reg  PDC ;
reg  PDD ;
reg  PDE ;
reg  PDF ;
reg  PEA ;
reg  PEB ;
reg  QAA ;
reg  QAB ;
reg  QAC ;
reg  QAD ;
reg  QAE ;
reg  QAF ;
reg  QAG ;
reg  QAH ;
reg  QAI ;
reg  QBA ;
reg  QBB ;
reg  QBC ;
reg  QBD ;
reg  QBE ;
reg  QBF ;
reg  QBG ;
reg  QBH ;
reg  QBI ;
reg  QBJ ;
reg  QCB ;
reg  QCD ;
reg  QCF ;
reg  QCH ;
reg  QCJ ;
reg  QDA ;
reg  QDB ;
reg  QDC ;
reg  QDD ;
reg  QDE ;
reg  QDF ;
reg  QDG ;
reg  QDH ;
reg  QDI ;
reg  QDJ ;
reg  QEA ;
reg  QEB ;
reg  qfa ;
reg  qfb ;
reg  QGA ;
reg  QGB ;
reg  QGC ;
reg  QGD ;
reg  QGE ;
reg  QGF ;
reg  QHA ;
reg  QHB ;
reg  QHC ;
reg  QHD ;
reg  qhe ;
reg  qhf ;
reg  qhg ;
reg  qhh ;
reg  qhi ;
reg  qhj ;
reg  qhk ;
reg  qhl ;
reg  qhm ;
reg  qhn ;
reg  qho ;
reg  qhp ;
reg  qhq ;
reg  qhr ;
reg  qhs ;
reg  qht ;
reg  qia ;
reg  qib ;
reg  qic ;
reg  QJA ;
reg  QJB ;
reg  QLA ;
reg  QMA ;
reg  QMB ;
reg  qmc ;
reg  qmd ;
reg  QME ;
reg  QMF ;
reg  QNA ;
reg  QNB ;
reg  QNC ;
reg  QND ;
reg  QNE ;
reg  QNF ;
reg  QNG ;
reg  QPA ;
reg  QPB ;
reg  QQA ;
reg  QQB ;
reg  QQC ;
reg  QRA ;
reg  TBA ;
reg  TBB ;
reg  TBC ;
reg  TBD ;
reg  TBE ;
reg  TBF ;
reg  TBG ;
reg  TBH ;
reg  TCA ;
reg  TCB ;
reg  TDA ;
reg  TDB ;
reg  TEA ;
reg  TEB ;
reg  TEC ;
reg  TED ;
reg  TEE ;
reg  TGA ;
reg  TGB ;
reg  TGC ;
reg  TGD ;
reg  tge ;
reg  tgf ;
reg  tgg ;
reg  tgh ;
reg  THA ;
reg  THB ;
reg  TIA ;
reg  TIB ;
reg  TJA ;
reg  TJB ;
reg  TKA ;
reg  TKB ;
reg  TLA ;
reg  TLB ;
reg  tlc ;
reg  tld ;
reg  TMA ;
reg  TMB ;
reg  tmc ;
reg  tmd ;
reg  TNA ;
reg  TNB ;
reg  tnc ;
reg  tnd ;
reg  TOA ;
reg  TOB ;
reg  toc ;
reg  tod ;
reg  TPA ;
reg  TPB ;
reg  TPC ;
reg  TPD ;
reg  tqa ;
reg  TQB ;
reg  tqc ;
reg  TQD ;
reg  tqe ;
reg  TQF ;
reg  tqg ;
reg  TQH ;
reg  tqi ;
reg  TQJ ;
reg  tqk ;
reg  TQL ;
reg  tqm ;
reg  TQN ;
reg  tqo ;
reg  TQP ;
reg  tqq ;
reg  TQR ;
reg  tqs ;
reg  TQT ;
reg  tra ;
reg  TRB ;
reg  trc ;
reg  TRD ;
reg  tre ;
reg  TRF ;
reg  trg ;
reg  TRH ;
reg  trii ;
reg  TRJ ;
reg  trk ;
reg  TRL ;
reg  trm ;
reg  TRN ;
reg  tro ;
reg  TRP ;
reg  trq ;
reg  TRR ;
reg  trs ;
reg  TRT ;
reg  tsa ;
reg  TSB ;
reg  tsc ;
reg  TSD ;
reg  tse ;
reg  TSF ;
reg  tsg ;
reg  TSH ;
reg  tsi ;
reg  TSJ ;
reg  tsk ;
reg  TSL ;
reg  tsm ;
reg  TSN ;
reg  tso ;
reg  TSP ;
reg  tsq ;
reg  TSR ;
reg  tss ;
reg  TST ;
reg  tta ;
reg  TTB ;
reg  ttc ;
reg  TTD ;
reg  tte ;
reg  TTF ;
reg  ttg ;
reg  TTH ;
reg  tti ;
reg  TTJ ;
reg  ttk ;
reg  TTL ;
reg  ttm ;
reg  TTN ;
reg  tto ;
reg  TTP ;
reg  ttq ;
reg  TTR ;
reg  tts ;
reg  TTT ;
reg  TUA ;
reg  TUB ;
reg  TUC ;
reg  TUD ;
reg  WAA ;
reg  WAB ;
reg  WAC ;
reg  WAD ;
reg  WAE ;
reg  WAF ;
reg  WAG ;
reg  WAH ;
reg  WBA ;
reg  WBB ;
reg  WBC ;
reg  WBD ;
reg  WBE ;
reg  WBF ;
reg  WBG ;
reg  WBH ;
reg  WCA ;
reg  WCB ;
reg  WCC ;
reg  WCD ;
reg  WCE ;
reg  WCF ;
reg  WCG ;
reg  WCH ;
reg  WDA ;
reg  WDB ;
reg  WDC ;
reg  WDD ;
reg  WDE ;
reg  WDF ;
reg  WDG ;
reg  WDH ;
reg  WEA ;
reg  WEB ;
reg  WEC ;
reg  WED ;
reg  WEE ;
reg  WEF ;
reg  WEG ;
reg  WEH ;
wire  aaa ;
wire  aab ;
wire  aac ;
wire  aad ;
wire  aae ;
wire  aaf ;
wire  aag ;
wire  aah ;
wire  aai ;
wire  aaj ;
wire  aak ;
wire  aal ;
wire  aba ;
wire  abb ;
wire  abc ;
wire  abd ;
wire  abe ;
wire  abf ;
wire  abg ;
wire  abh ;
wire  abi ;
wire  abj ;
wire  abk ;
wire  abl ;
wire  aca ;
wire  acb ;
wire  acc ;
wire  acd ;
wire  ace ;
wire  acf ;
wire  acg ;
wire  ach ;
wire  aci ;
wire  acj ;
wire  ack ;
wire  acl ;
wire  adb ;
wire  adc ;
wire  add ;
wire  ade ;
wire  adf ;
wire  adg ;
wire  adh ;
wire  adi ;
wire  adj ;
wire  adk ;
wire  adl ;
wire  aea ;
wire  aeb ;
wire  aec ;
wire  aed ;
wire  aee ;
wire  aef ;
wire  aeg ;
wire  aeh ;
wire  aei ;
wire  aej ;
wire  aek ;
wire  ael ;
wire  afa ;
wire  afb ;
wire  afc ;
wire  afd ;
wire  afe ;
wire  aff ;
wire  afg ;
wire  afh ;
wire  afi ;
wire  afj ;
wire  afk ;
wire  afl ;
wire  AGB ;
wire  AGC ;
wire  AGD ;
wire  AGE ;
wire  AGF ;
wire  AGG ;
wire  AGH ;
wire  AGI ;
wire  AGJ ;
wire  AGK ;
wire  AGL ;
wire  AHA ;
wire  AHB ;
wire  AHC ;
wire  AHD ;
wire  AHE ;
wire  AHF ;
wire  AHG ;
wire  AHH ;
wire  AHI ;
wire  AHJ ;
wire  AHK ;
wire  AHL ;
wire  AIA ;
wire  AIB ;
wire  AIC ;
wire  AID ;
wire  AIE ;
wire  AIF ;
wire  AIG ;
wire  AIH ;
wire  AII ;
wire  AIJ ;
wire  AIK ;
wire  AIL ;
wire  AJB ;
wire  AJC ;
wire  AJD ;
wire  AJE ;
wire  AJF ;
wire  AJG ;
wire  AJH ;
wire  AJI ;
wire  AJJ ;
wire  AJK ;
wire  AJL ;
wire  AKA ;
wire  AKB ;
wire  AKC ;
wire  AKD ;
wire  AKE ;
wire  AKF ;
wire  AKG ;
wire  AKH ;
wire  AKI ;
wire  AKJ ;
wire  AKK ;
wire  AKL ;
wire  ALA ;
wire  ALB ;
wire  ALC ;
wire  ALD ;
wire  ALE ;
wire  ALF ;
wire  ALG ;
wire  ALH ;
wire  ALI ;
wire  ALJ ;
wire  ALK ;
wire  ALL ;
wire  ama ;
wire  amb ;
wire  amc ;
wire  amd ;
wire  ame ;
wire  amf ;
wire  amg ;
wire  amh ;
wire  ami ;
wire  amj ;
wire  amk ;
wire  aml ;
wire  amm ;
wire  amn ;
wire  amo ;
wire  amp ;
wire  bak ;
wire  bal ;
wire  bam ;
wire  ban ;
wire  bao ;
wire  bap ;
wire  baq ;
wire  bar ;
wire  bas ;
wire  bat ;
wire  bau ;
wire  bav ;
wire  baw ;
wire  bax ;
wire  bay ;
wire  baz ;
wire  BBA ;
wire  BBB ;
wire  BBC ;
wire  BBD ;
wire  BBE ;
wire  BBF ;
wire  BBG ;
wire  BBH ;
wire  BBI ;
wire  BBJ ;
wire  BBK ;
wire  BBL ;
wire  BBM ;
wire  BBN ;
wire  BBO ;
wire  BBP ;
wire  bca ;
wire  bcb ;
wire  bcc ;
wire  bcd ;
wire  bce ;
wire  bcf ;
wire  bcg ;
wire  bch ;
wire  bci ;
wire  bcj ;
wire  bck ;
wire  bcl ;
wire  bcm ;
wire  bcn ;
wire  bco ;
wire  bcp ;
wire  bda ;
wire  bdb ;
wire  bdc ;
wire  bdd ;
wire  bde ;
wire  bdf ;
wire  bdg ;
wire  bdh ;
wire  bdi ;
wire  bdj ;
wire  bdk ;
wire  bdl ;
wire  bdm ;
wire  bdn ;
wire  bdo ;
wire  bdp ;
wire  bea ;
wire  beb ;
wire  bec ;
wire  bed ;
wire  bee ;
wire  bef ;
wire  beg ;
wire  beh ;
wire  bei ;
wire  bej ;
wire  bek ;
wire  bel ;
wire  bem ;
wire  ben ;
wire  beo ;
wire  bep ;
wire  bfa ;
wire  bfb ;
wire  bfc ;
wire  caa ;
wire  CAA ;
wire  cab ;
wire  CAB ;
wire  cac ;
wire  CAC ;
wire  cad ;
wire  CAD ;
wire  cae ;
wire  CAE ;
wire  caf ;
wire  CAF ;
wire  cag ;
wire  CAG ;
wire  cah ;
wire  CAH ;
wire  cai ;
wire  CAI ;
wire  caj ;
wire  CAJ ;
wire  cak ;
wire  CAK ;
wire  cal ;
wire  CAL ;
wire  cam ;
wire  CAM ;
wire  can ;
wire  CAN ;
wire  cao ;
wire  CAO ;
wire  cap ;
wire  CAP ;
wire  daa ;
wire  dab ;
wire  dac ;
wire  dad ;
wire  dae ;
wire  daf ;
wire  dag ;
wire  dah ;
wire  dba ;
wire  dbb ;
wire  dbc ;
wire  dbd ;
wire  dbe ;
wire  dbf ;
wire  dbg ;
wire  dbh ;
wire  DCA ;
wire  DCB ;
wire  DCC ;
wire  DCD ;
wire  DCE ;
wire  DCF ;
wire  DCG ;
wire  DCH ;
wire  DDA ;
wire  DDB ;
wire  DDC ;
wire  DDD ;
wire  DDE ;
wire  DDF ;
wire  DDG ;
wire  DDH ;
wire  dia ;
wire  dib ;
wire  dic ;
wire  did ;
wire  die ;
wire  dif ;
wire  dig ;
wire  dih ;
wire  EAA ;
wire  EAB ;
wire  EAC ;
wire  EAD ;
wire  EAE ;
wire  EAF ;
wire  EAG ;
wire  EAH ;
wire  EAI ;
wire  EAJ ;
wire  EAK ;
wire  EAL ;
wire  EBA ;
wire  EBB ;
wire  EBC ;
wire  EBD ;
wire  EBE ;
wire  EBF ;
wire  EBG ;
wire  EBH ;
wire  EBI ;
wire  EBJ ;
wire  EBK ;
wire  EBL ;
wire  ECA ;
wire  ECB ;
wire  ECC ;
wire  ECD ;
wire  ECE ;
wire  ECF ;
wire  ECG ;
wire  ECH ;
wire  ECI ;
wire  ECJ ;
wire  ECK ;
wire  ECL ;
wire  fab ;
wire  FAB ;
wire  fac ;
wire  FAC ;
wire  fad ;
wire  FAD ;
wire  fae ;
wire  FAE ;
wire  faf ;
wire  FAF ;
wire  fag ;
wire  FAG ;
wire  fah ;
wire  FAH ;
wire  fai ;
wire  FAI ;
wire  faj ;
wire  FAJ ;
wire  fak ;
wire  FAK ;
wire  fal ;
wire  FAL ;
wire  FBA ;
wire  FBB ;
wire  FCA ;
wire  iaa ;
wire  iab ;
wire  iac ;
wire  iad ;
wire  iae ;
wire  iaf ;
wire  iag ;
wire  iah ;
wire  iai ;
wire  iaj ;
wire  iak ;
wire  ial ;
wire  iam ;
wire  ian ;
wire  iao ;
wire  iap ;
wire  ica ;
wire  icb ;
wire  icc ;
wire  icd ;
wire  ice ;
wire  icf ;
wire  icg ;
wire  ich ;
wire  ici ;
wire  icj ;
wire  ick ;
wire  icl ;
wire  icm ;
wire  icn ;
wire  ico ;
wire  icp ;
wire  iga ;
wire  ija ;
wire  ika ;
wire  ila ;
wire  ilb ;
wire  ilc ;
wire  ild ;
wire  ile ;
wire  ilf ;
wire  ilg ;
wire  ilh ;
wire  ili ;
wire  ipa ;
wire  ipb ;
wire  iqa ;
wire  iqb ;
wire  iqc ;
wire  ira ;
wire  irb ;
wire  isa ;
wire  naa ;
wire  NAA ;
wire  nab ;
wire  NAB ;
wire  nac ;
wire  NAC ;
wire  nad ;
wire  NAD ;
wire  nae ;
wire  NAE ;
wire  naf ;
wire  NAF ;
wire  nag ;
wire  NAG ;
wire  nah ;
wire  NAH ;
wire  nai ;
wire  NAI ;
wire  naj ;
wire  NAJ ;
wire  nak ;
wire  NAK ;
wire  nal ;
wire  NAL ;
wire  nam ;
wire  NAM ;
wire  nan ;
wire  NAN ;
wire  nao ;
wire  NAO ;
wire  nap ;
wire  NAP ;
wire  naq ;
wire  NAQ ;
wire  nar ;
wire  NAR ;
wire  nas ;
wire  NAS ;
wire  nat ;
wire  NAT ;
wire  nba ;
wire  NBA ;
wire  nbb ;
wire  NBB ;
wire  nbc ;
wire  NBC ;
wire  nbd ;
wire  NBD ;
wire  nbe ;
wire  NBE ;
wire  nbf ;
wire  NBF ;
wire  nbg ;
wire  NBG ;
wire  nbh ;
wire  NBH ;
wire  nbi ;
wire  NBI ;
wire  nbj ;
wire  NBJ ;
wire  nbk ;
wire  NBK ;
wire  nbl ;
wire  NBL ;
wire  nbm ;
wire  NBM ;
wire  nbn ;
wire  NBN ;
wire  nbo ;
wire  NBO ;
wire  nbp ;
wire  NBP ;
wire  nbq ;
wire  NBQ ;
wire  nbr ;
wire  NBR ;
wire  nbs ;
wire  NBS ;
wire  nbt ;
wire  NBT ;
wire  oaa ;
wire  oab ;
wire  oac ;
wire  oad ;
wire  oae ;
wire  oaf ;
wire  oag ;
wire  oah ;
wire  oai ;
wire  oaj ;
wire  oak ;
wire  oal ;
wire  oam ;
wire  oan ;
wire  oao ;
wire  oap ;
wire  oaq ;
wire  oar ;
wire  oas ;
wire  oat ;
wire  oau ;
wire  oav ;
wire  oaw ;
wire  oax ;
wire  oay ;
wire  oaz ;
wire  oba ;
wire  obb ;
wire  obc ;
wire  obd ;
wire  obe ;
wire  obf ;
wire  obg ;
wire  obh ;
wire  obi ;
wire  obj ;
wire  obk ;
wire  obl ;
wire  obm ;
wire  obn ;
wire  obo ;
wire  obp ;
wire  obq ;
wire  obr ;
wire  obs ;
wire  obt ;
wire  obu ;
wire  obv ;
wire  obw ;
wire  obx ;
wire  oby ;
wire  obz ;
wire  oca ;
wire  ocb ;
wire  occ ;
wire  ocd ;
wire  oce ;
wire  ocf ;
wire  ocg ;
wire  och ;
wire  oci ;
wire  ocj ;
wire  ock ;
wire  ocl ;
wire  ocm ;
wire  ocn ;
wire  oco ;
wire  ocp ;
wire  ocq ;
wire  ocr ;
wire  ocs ;
wire  oct ;
wire  ocu ;
wire  ocv ;
wire  ocw ;
wire  ocx ;
wire  ocy ;
wire  ocz ;
wire  oda ;
wire  odb ;
wire  odc ;
wire  odd ;
wire  ode ;
wire  odf ;
wire  odg ;
wire  odh ;
wire  odi ;
wire  odj ;
wire  odk ;
wire  odl ;
wire  odm ;
wire  odn ;
wire  odo ;
wire  odp ;
wire  odq ;
wire  odr ;
wire  ods ;
wire  odt ;
wire  odu ;
wire  odv ;
wire  odw ;
wire  odx ;
wire  ody ;
wire  odz ;
wire  oea ;
wire  oeb ;
wire  oec ;
wire  oed ;
wire  oee ;
wire  oef ;
wire  oeg ;
wire  oeh ;
wire  oei ;
wire  oej ;
wire  oek ;
wire  oel ;
wire  oem ;
wire  oen ;
wire  oeo ;
wire  oep ;
wire  ofa ;
wire  ofb ;
wire  ofc ;
wire  ofd ;
wire  ofe ;
wire  off ;
wire  ofg ;
wire  ofh ;
wire  ofi ;
wire  ofj ;
wire  ofk ;
wire  ofl ;
wire  ofm ;
wire  ofn ;
wire  ofo ;
wire  ofp ;
wire  OGA ;
wire  OGB ;
wire  OGC ;
wire  OGD ;
wire  OGE ;
wire  OGF ;
wire  OGG ;
wire  OGH ;
wire  OGI ;
wire  OGJ ;
wire  OGK ;
wire  OGL ;
wire  OGM ;
wire  OGN ;
wire  OGO ;
wire  OGP ;
wire  OHA ;
wire  OHB ;
wire  OHC ;
wire  OHD ;
wire  OHE ;
wire  OHF ;
wire  OHG ;
wire  OHH ;
wire  OHI ;
wire  OHJ ;
wire  OHK ;
wire  OHL ;
wire  OHM ;
wire  OHN ;
wire  OHO ;
wire  OHP ;
wire  oia ;
wire  oib ;
wire  oic ;
wire  oid ;
wire  oie ;
wire  oif ;
wire  oig ;
wire  oih ;
wire  oii ;
wire  oij ;
wire  oik ;
wire  oil ;
wire  oim ;
wire  OJA ;
wire  oka ;
wire  okb ;
wire  okc ;
wire  okd ;
wire  oke ;
wire  okf ;
wire  okg ;
wire  ola ;
wire  olb ;
wire  olc ;
wire  old ;
wire  ole ;
wire  olf ;
wire  olg ;
wire  olh ;
wire  oli ;
wire  oma ;
wire  ona ;
wire  PAA ;
wire  PAB ;
wire  PAC ;
wire  PAD ;
wire  PAE ;
wire  PAF ;
wire  PAG ;
wire  PAH ;
wire  PAI ;
wire  PAJ ;
wire  PAK ;
wire  PAL ;
wire  PAM ;
wire  PAN ;
wire  PAO ;
wire  PAP ;
wire  PAQ ;
wire  PAR ;
wire  PAS ;
wire  PAT ;
wire  PBA ;
wire  PBB ;
wire  PBC ;
wire  PBD ;
wire  PBE ;
wire  PBF ;
wire  PBG ;
wire  PBH ;
wire  PBI ;
wire  PBJ ;
wire  PBK ;
wire  PBL ;
wire  PBM ;
wire  PBN ;
wire  PBO ;
wire  PBP ;
wire  PBQ ;
wire  PBR ;
wire  PBS ;
wire  PBT ;
wire  pca ;
wire  pcb ;
wire  pcc ;
wire  pcd ;
wire  pce ;
wire  pcf ;
wire  pcg ;
wire  pch ;
wire  pci ;
wire  pcj ;
wire  pck ;
wire  pcl ;
wire  pcm ;
wire  pcn ;
wire  pda ;
wire  pdb ;
wire  pdc ;
wire  pdd ;
wire  pde ;
wire  pdf ;
wire  pea ;
wire  peb ;
wire  qaa ;
wire  qab ;
wire  qac ;
wire  qad ;
wire  qae ;
wire  qaf ;
wire  qag ;
wire  qah ;
wire  qai ;
wire  qba ;
wire  qbb ;
wire  qbc ;
wire  qbd ;
wire  qbe ;
wire  qbf ;
wire  qbg ;
wire  qbh ;
wire  qbi ;
wire  qbj ;
wire  qcb ;
wire  qcd ;
wire  qcf ;
wire  qch ;
wire  qcj ;
wire  qda ;
wire  qdb ;
wire  qdc ;
wire  qdd ;
wire  qde ;
wire  qdf ;
wire  qdg ;
wire  qdh ;
wire  qdi ;
wire  qdj ;
wire  qea ;
wire  qeb ;
wire  QFA ;
wire  QFB ;
wire  qga ;
wire  qgb ;
wire  qgc ;
wire  qgd ;
wire  qge ;
wire  qgf ;
wire  qha ;
wire  qhb ;
wire  qhc ;
wire  qhd ;
wire  QHE ;
wire  QHF ;
wire  QHG ;
wire  QHH ;
wire  QHI ;
wire  QHJ ;
wire  QHK ;
wire  QHL ;
wire  QHM ;
wire  QHN ;
wire  QHO ;
wire  QHP ;
wire  QHQ ;
wire  QHR ;
wire  QHS ;
wire  QHT ;
wire  QIA ;
wire  QIB ;
wire  QIC ;
wire  qja ;
wire  qjb ;
wire  qla ;
wire  qma ;
wire  qmb ;
wire  QMC ;
wire  QMD ;
wire  qme ;
wire  qmf ;
wire  qna ;
wire  qnb ;
wire  qnc ;
wire  qnd ;
wire  qne ;
wire  qnf ;
wire  qng ;
wire  qpa ;
wire  qpb ;
wire  qqa ;
wire  qqb ;
wire  qqc ;
wire  qra ;
wire  tba ;
wire  tbb ;
wire  tbc ;
wire  tbd ;
wire  tbe ;
wire  tbf ;
wire  tbg ;
wire  tbh ;
wire  tca ;
wire  tcb ;
wire  tda ;
wire  tdb ;
wire  tea ;
wire  teb ;
wire  tec ;
wire  ted ;
wire  tee ;
wire  tga ;
wire  tgb ;
wire  tgc ;
wire  tgd ;
wire  TGE ;
wire  TGF ;
wire  TGG ;
wire  TGH ;
wire  tha ;
wire  thb ;
wire  tia ;
wire  tib ;
wire  tja ;
wire  tjb ;
wire  tka ;
wire  tkb ;
wire  tla ;
wire  tlb ;
wire  TLC ;
wire  TLD ;
wire  tma ;
wire  tmb ;
wire  TMC ;
wire  TMD ;
wire  tna ;
wire  tnb ;
wire  TNC ;
wire  TND ;
wire  toa ;
wire  tob ;
wire  TOC ;
wire  TOD ;
wire  tpa ;
wire  tpb ;
wire  tpc ;
wire  tpd ;
wire  TQA ;
wire  tqb ;
wire  TQC ;
wire  tqd ;
wire  TQE ;
wire  tqf ;
wire  TQG ;
wire  tqh ;
wire  TQI ;
wire  tqj ;
wire  TQK ;
wire  tql ;
wire  TQM ;
wire  tqn ;
wire  TQO ;
wire  tqp ;
wire  TQQ ;
wire  tqr ;
wire  TQS ;
wire  tqt ;
wire  TRA ;
wire  trb ;
wire  TRC ;
wire  trd ;
wire  TRE ;
wire  trf ;
wire  TRG ;
wire  trh ;
wire  TRI ;
wire  trj ;
wire  TRK ;
wire  trl ;
wire  TRM ;
wire  trn ;
wire  TRO ;
wire  trp ;
wire  TRQ ;
wire  trr ;
wire  TRS ;
wire  trt ;
wire  TSA ;
wire  tsb ;
wire  TSC ;
wire  tsd ;
wire  TSE ;
wire  tsf ;
wire  TSG ;
wire  tsh ;
wire  TSI ;
wire  tsj ;
wire  TSK ;
wire  tsl ;
wire  TSM ;
wire  tsn ;
wire  TSO ;
wire  tsp ;
wire  TSQ ;
wire  tsr ;
wire  TSS ;
wire  tst ;
wire  TTA ;
wire  ttb ;
wire  TTC ;
wire  ttd ;
wire  TTE ;
wire  ttf ;
wire  TTG ;
wire  tth ;
wire  TTI ;
wire  ttj ;
wire  TTK ;
wire  ttl ;
wire  TTM ;
wire  ttn ;
wire  TTO ;
wire  ttp ;
wire  TTQ ;
wire  ttr ;
wire  TTS ;
wire  ttt ;
wire  tua ;
wire  tub ;
wire  tuc ;
wire  tud ;
wire  waa ;
wire  wab ;
wire  wac ;
wire  wad ;
wire  wae ;
wire  waf ;
wire  wag ;
wire  wah ;
wire  wba ;
wire  wbb ;
wire  wbc ;
wire  wbd ;
wire  wbe ;
wire  wbf ;
wire  wbg ;
wire  wbh ;
wire  wca ;
wire  wcb ;
wire  wcc ;
wire  wcd ;
wire  wce ;
wire  wcf ;
wire  wcg ;
wire  wch ;
wire  wda ;
wire  wdb ;
wire  wdc ;
wire  wdd ;
wire  wde ;
wire  wdf ;
wire  wdg ;
wire  wdh ;
wire  wea ;
wire  web ;
wire  wec ;
wire  wed ;
wire  wee ;
wire  wef ;
wire  weg ;
wire  weh ;
wire  ZZI ;
wire  ZZO ;

wire MAA;
wire MAB;
wire MAC;
wire MAD;
wire MAE;
wire MAF;
wire MAG;
wire MAH;
wire MAI;
wire MAJ;
wire MAK;
wire MAL;
wire MAM;
wire MAN;
wire MAO;
wire MAP;
wire MAQ;
wire MAR;
wire MAS;
wire MAT;
wire MBA;
wire MBB;
wire MBC;
wire MBD;
wire MBE;
wire MBF;
wire MBG;
wire MBH;
wire MBI;
wire MBJ;
wire MBK;
wire MBL;
wire MBM;
wire MBN;
wire MBO;
wire MBP;
wire MBQ;
wire MBR;
wire MBS;
wire MBT;
wire MCA;
wire MCB;
wire MCC;
wire MCD;
wire MCE;
wire MCF;
wire MCG;
wire MCH;
wire MCI;
wire MCJ;
wire MCK;
wire MCL;
wire MCM;
wire MCN;
wire MCO;
wire MCP;
wire MCQ;
wire MCR;
wire MCS;
wire MCT;
wire MDA;
wire MDB;
wire MDC;
wire MDD;
wire MDE;
wire MDF;
wire MDG;
wire MDH;
wire MDI;
wire MDJ;
wire MDK;
wire MDL;
wire MDM;
wire MDN;
wire MDO;
wire MDP;
wire MDQ;
wire MDR;
wire MDS;
wire MDT;
wire MEA;
wire MEB;
wire MEC;
wire MED;
wire MEE;
wire MEF;
wire MEG;
wire MEH;
wire MEI;
wire MEJ;
wire MEK;
wire MEL;
wire MEM;
wire MEN;
wire MEO;
wire MEP;
wire MEQ;
wire MER;
wire MES;
wire MET;
wire MFA;
wire MFB;
wire MFC;
wire MFD;
wire MFE;
wire MFF;
wire MFG;
wire MFH;
wire MFI;
wire MFJ;
wire MFK;
wire MFL;
wire MFM;
wire MFN;
wire MFO;
wire MFP;
wire MFQ;
wire MFR;
wire MFS;
wire MFT;
wire MGA;
wire MGB;
wire MGC;
wire MGD;      
wire MGE;
wire MGF;
wire MGG;
wire MGH;
wire MGI;
wire MGJ;
wire MGK;
wire MGL;
wire MGM;
wire MGN;
wire MGO;
wire MGP;
wire MGQ;
wire MGR;
wire MGS;
wire MGT;
wire MHA;
wire MHB;
wire MHC;
wire MHD;
wire MHE;
wire MHF;
wire MHG;
wire MHH;
wire MHI;
wire MHJ;
wire MHK;
wire MHL;
wire MHM;
wire MHN;
wire MHO;
wire MHP;
wire MHQ;
wire MHR;
wire MHS;
wire MHT;

assign ZZI = 1'b1;
assign ZZO = 1'b0;
assign wde = ~WDE;  //complement 
assign wdf = ~WDF;  //complement 
assign wdg = ~WDG;  //complement 
assign wdh = ~WDH;  //complement 
assign tqt = ~TQT;  //complement 
assign trt = ~TRT;  //complement 
assign tst = ~TST;  //complement 
assign ttt = ~TTT;  //complement 
assign wea = ~WEA;  //complement 
assign web = ~WEB;  //complement 
assign wec = ~WEC;  //complement 
assign wed = ~WED;  //complement 
assign wda = ~WDA;  //complement 
assign wdb = ~WDB;  //complement 
assign wdc = ~WDC;  //complement 
assign wdd = ~WDD;  //complement 
assign pca = ~PCA;  //complement 
assign pdf = ~PDF;  //complement 
assign NBF =  MBF & TQN  |  MDF & TRN  |  MFF & TSN  |  MHF & TTM  ; 
assign nbf = ~NBF;  //complement 
assign wee = ~WEE;  //complement 
assign wef = ~WEF;  //complement 
assign weg = ~WEG;  //complement 
assign weh = ~WEH;  //complement 
assign NBM =  MBM & TQQ  |  MDM & TRQ  |  MFM & TSQ  |  MHM & TTQ  ; 
assign nbm = ~NBM;  //complement 
assign TQO = ~tqo;  //complement 
assign TRO = ~tro;  //complement 
assign TSO = ~tso;  //complement 
assign TTO = ~tto;  //complement 
assign PAA = ~paa;  //complement 
assign PAQ = ~paq;  //complement 
assign PBM = ~pbm;  //complement 
assign QHI = ~qhi;  //complement 
assign QHJ = ~qhj;  //complement 
assign QHE = ~qhe;  //complement 
assign QHF = ~qhf;  //complement 
assign NAQ =  MAQ & TQI  |  MCQ & TRI  |  MEQ & TSI  |  MGQ & TTT  ; 
assign naq = ~NAQ;  //complement 
assign tql = ~TQL;  //complement 
assign trl = ~TRL;  //complement 
assign tsl = ~TSL;  //complement 
assign ttl = ~TTL;  //complement 
assign tqh = ~TQH;  //complement 
assign trh = ~TRH;  //complement 
assign tsh = ~TSH;  //complement 
assign tth = ~TTH;  //complement 
assign NAJ =  MAJ & TQF  |  MCJ & TRF  |  MEJ & TSF  |  MGJ & TTF  ; 
assign naj = ~NAJ;  //complement 
assign PAJ = ~paj;  //complement 
assign PBF = ~pbf;  //complement 
assign CAE =  BAO & TCA  |  AME & TDA  ; 
assign cae = ~CAE;  //complement 
assign CAG =  BAQ & TCA  |  AMG & TDA  ; 
assign cag = ~CAG;  //complement 
assign oaa = ~OAA;  //complement 
assign oba = ~OBA;  //complement 
assign oca = ~OCA;  //complement 
assign oda = ~ODA;  //complement 
assign bao = ~BAO;  //complement 
assign oao = ~OAO;  //complement 
assign obo = ~OBO;  //complement 
assign TLC = ~tlc;  //complement 
assign TLD = ~tld;  //complement 
assign daa = ~DAA;  //complement 
assign dae = ~DAE;  //complement 
assign oig = ~OIG;  //complement 
assign TRC = ~trc;  //complement 
assign baq = ~BAQ;  //complement 
assign oaq = ~OAQ;  //complement 
assign obq = ~OBQ;  //complement 
assign tga = ~TGA;  //complement 
assign tgb = ~TGB;  //complement 
assign tgc = ~TGC;  //complement 
assign tgd = ~TGD;  //complement 
assign amm = ~AMM;  //complement 
assign oem = ~OEM;  //complement 
assign ofm = ~OFM;  //complement 
assign TQC = ~tqc;  //complement 
assign TSC = ~tsc;  //complement 
assign TTC = ~ttc;  //complement 
assign NAA =  MAA & TQA  |  MCA & TRA  |  MEA & TSA  |  MGA & TTA  ; 
assign naa = ~NAA;  //complement 
assign ame = ~AME;  //complement 
assign oee = ~OEE;  //complement 
assign ofe = ~OFE;  //complement 
assign aai = ~AAI;  //complement 
assign abi = ~ABI;  //complement 
assign aci = ~ACI;  //complement 
assign amj = ~AMJ;  //complement 
assign aba = ~ABA;  //complement 
assign aca = ~ACA;  //complement 
assign aae = ~AAE;  //complement 
assign abe = ~ABE;  //complement 
assign ace = ~ACE;  //complement 
assign aaa = ~AAA;  //complement 
assign aab = ~AAB;  //complement 
assign abb = ~ABB;  //complement 
assign acb = ~ACB;  //complement 
assign aaf = ~AAF;  //complement 
assign abf = ~ABF;  //complement 
assign acf = ~ACF;  //complement 
assign waa = ~WAA;  //complement 
assign wab = ~WAB;  //complement 
assign wac = ~WAC;  //complement 
assign wad = ~WAD;  //complement 
assign wae = ~WAE;  //complement 
assign waf = ~WAF;  //complement 
assign wag = ~WAG;  //complement 
assign wah = ~WAH;  //complement 
assign oej = ~OEJ;  //complement 
assign ofj = ~OFJ;  //complement 
assign aaj = ~AAJ;  //complement 
assign abj = ~ABJ;  //complement 
assign acj = ~ACJ;  //complement 
assign dab = ~DAB;  //complement 
assign daf = ~DAF;  //complement 
assign baz = ~BAZ;  //complement 
assign oaz = ~OAZ;  //complement 
assign obz = ~OBZ;  //complement 
assign qpa = ~QPA;  //complement 
assign qpb = ~QPB;  //complement 
assign amd = ~AMD;  //complement 
assign oed = ~OED;  //complement 
assign ofd = ~OFD;  //complement 
assign CAN =  BAX & TCB  |  AMN & TDB  ; 
assign can = ~CAN;  //complement 
assign CAP =  BAZ & TCB  |  AMP & TDB  ; 
assign cap = ~CAP;  //complement 
assign oaj = ~OAJ;  //complement 
assign obj = ~OBJ;  //complement 
assign ocj = ~OCJ;  //complement 
assign odj = ~ODJ;  //complement 
assign bax = ~BAX;  //complement 
assign oax = ~OAX;  //complement 
assign obx = ~OBX;  //complement 
assign tba = ~TBA;  //complement 
assign tbe = ~TBE;  //complement 
assign tpa = ~TPA;  //complement 
assign tua = ~TUA;  //complement 
assign pcb = ~PCB;  //complement 
assign pea = ~PEA;  //complement 
assign pcc = ~PCC;  //complement 
assign pde = ~PDE;  //complement 
assign NBT =  MBT & TQT  |  MDT & TRT  |  MFT & TST  |  MHT & TTT  ; 
assign nbt = ~NBT;  //complement 
assign tqr = ~TQR;  //complement 
assign trr = ~TRR;  //complement 
assign tsr = ~TSR;  //complement 
assign ttr = ~TTR;  //complement 
assign NBK =  MBK & TQO  |  MDK & TRO  |  MFK & TSO  |  MHK & TTO  ; 
assign nbk = ~NBK;  //complement 
assign TQM = ~tqm;  //complement 
assign TRM = ~trm;  //complement 
assign TSM = ~tsm;  //complement 
assign TTM = ~ttm;  //complement 
assign oai = ~OAI;  //complement 
assign PAO = ~pao;  //complement 
assign PBK = ~pbk;  //complement 
assign QHQ = ~qhq;  //complement 
assign QHR = ~qhr;  //complement 
assign QHM = ~qhm;  //complement 
assign QHN = ~qhn;  //complement 
assign NAO =  MAO & TQG  |  MCO & TRG  |  MEO & TSG  |  MGO & TTG  ; 
assign nao = ~NAO;  //complement 
assign TQE = ~tqe;  //complement 
assign TRE = ~tre;  //complement 
assign TSE = ~tse;  //complement 
assign TTE = ~tte;  //complement 
assign ttj = ~TTJ;  //complement 
assign NBD =  MBD & TQL  |  MDD & TRL  |  MFD & TSL  |  MHD & TTL  ; 
assign nbd = ~NBD;  //complement 
assign tqj = ~TQJ;  //complement 
assign trj = ~TRJ;  //complement 
assign tsj = ~TSJ;  //complement 
assign PAH = ~pah;  //complement 
assign PBD = ~pbd;  //complement 
assign PBT = ~pbt;  //complement 
assign ocb = ~OCB;  //complement 
assign qja = ~QJA;  //complement 
assign qjb = ~QJB;  //complement 
assign tca = ~TCA;  //complement 
assign tda = ~TDA;  //complement 
assign ona = ~ONA;  //complement 
assign oco = ~OCO;  //complement 
assign odo = ~ODO;  //complement 
assign tha = ~THA;  //complement 
assign thb = ~THB;  //complement 
assign tla = ~TLA;  //complement 
assign tlb = ~TLB;  //complement 
assign dac = ~DAC;  //complement 
assign dag = ~DAG;  //complement 
assign oie = ~OIE;  //complement 
assign ocq = ~OCQ;  //complement 
assign odq = ~ODQ;  //complement 
assign amo = ~AMO;  //complement 
assign oeo = ~OEO;  //complement 
assign ofo = ~OFO;  //complement 
assign qqc = ~QQC;  //complement 
assign odx = ~ODX;  //complement 
assign amk = ~AMK;  //complement 
assign oek = ~OEK;  //complement 
assign ofk = ~OFK;  //complement 
assign aak = ~AAK;  //complement 
assign abk = ~ABK;  //complement 
assign ack = ~ACK;  //complement 
assign aac = ~AAC;  //complement 
assign abc = ~ABC;  //complement 
assign acc = ~ACC;  //complement 
assign aag = ~AAG;  //complement 
assign abg = ~ABG;  //complement 
assign acg = ~ACG;  //complement 
assign aad = ~AAD;  //complement 
assign abd = ~ABD;  //complement 
assign acd = ~ACD;  //complement 
assign aah = ~AAH;  //complement 
assign abh = ~ABH;  //complement 
assign ach = ~ACH;  //complement 
assign NAH =  MAH & TQD  |  MCH & TRD  |  MEH & TSD  |  MGH & TTD  ; 
assign nah = ~NAH;  //complement 
assign tqb = ~TQB;  //complement 
assign trb = ~TRB;  //complement 
assign tsb = ~TSB;  //complement 
assign ttb = ~TTB;  //complement 
assign amh = ~AMH;  //complement 
assign oeh = ~OEH;  //complement 
assign ofh = ~OFH;  //complement 
assign aal = ~AAL;  //complement 
assign abl = ~ABL;  //complement 
assign acl = ~ACL;  //complement 
assign dad = ~DAD;  //complement 
assign dah = ~DAH;  //complement 
assign ocz = ~OCZ;  //complement 
assign odz = ~ODZ;  //complement 
assign qqb = ~QQB;  //complement 
assign amb = ~AMB;  //complement 
assign oeb = ~OEB;  //complement 
assign ofb = ~OFB;  //complement 
assign tcb = ~TCB;  //complement 
assign tdb = ~TDB;  //complement 
assign oah = ~OAH;  //complement 
assign obh = ~OBH;  //complement 
assign och = ~OCH;  //complement 
assign odh = ~ODH;  //complement 
assign ocx = ~OCX;  //complement 
assign tbb = ~TBB;  //complement 
assign tbf = ~TBF;  //complement 
assign tpb = ~TPB;  //complement 
assign tub = ~TUB;  //complement 
assign qbb = ~QBB;  //complement 
assign qcb = ~QCB;  //complement 
assign qdc = ~QDC;  //complement 
assign qde = ~QDE;  //complement 
assign qea = ~QEA;  //complement 
assign qeb = ~QEB;  //complement 
assign qdd = ~QDD;  //complement 
assign qbd = ~QBD;  //complement 
assign qcd = ~QCD;  //complement 
assign pdd = ~PDD;  //complement 
assign pce = ~PCE;  //complement 
assign NBN =  MBN & TQR  |  MDN & TRR  |  MFN & TSR  |  MHN & TTR  ; 
assign nbn = ~NBN;  //complement 
assign pcd = ~PCD;  //complement 
assign PAB = ~pab;  //complement 
assign PAR = ~par;  //complement 
assign PBN = ~pbn;  //complement 
assign NBE =  MBE & TQM  |  MDE & TRM  |  MFE & TSM  |  MHE & TTM  ; 
assign nbe = ~NBE;  //complement 
assign PAI = ~pai;  //complement 
assign PBE = ~pbe;  //complement 
assign qae = ~QAE;  //complement 
assign qag = ~QAG;  //complement 
assign qbg = ~QBG;  //complement 
assign qbi = ~QBI;  //complement 
assign QIA = ~qia;  //complement 
assign QIB = ~qib;  //complement 
assign QIC = ~qic;  //complement 
assign NAI =  MAI & TQE  |  MCI & TRE  |  MEI & TSE  |  MGI & TTE  ; 
assign nai = ~NAI;  //complement 
assign qbf = ~QBF;  //complement 
assign qcf = ~QCF;  //complement 
assign NAR =  MAR & TQJ  |  MCR & TRJ  |  MER & TSJ  |  MGR & TTJ  ; 
assign nar = ~NAR;  //complement 
assign qbh = ~QBH;  //complement 
assign qch = ~QCH;  //complement 
assign qba = ~QBA;  //complement 
assign qbc = ~QBC;  //complement 
assign qbe = ~QBE;  //complement 
assign qdb = ~QDB;  //complement 
assign qaa = ~QAA;  //complement 
assign qdi = ~QDI;  //complement 
assign qdj = ~QDJ;  //complement 
assign qac = ~QAC;  //complement 
assign qai = ~QAI;  //complement 
assign qab = ~QAB;  //complement 
assign qad = ~QAD;  //complement 
assign qaf = ~QAF;  //complement 
assign qah = ~QAH;  //complement 
assign qdf = ~QDF;  //complement 
assign qdg = ~QDG;  //complement 
assign qdh = ~QDH;  //complement 
assign CAM =  BAW & TCA  |  AMM & TDA  ; 
assign cam = ~CAM;  //complement 
assign CAO =  BAY & TCA  |  AMO & TDA  ; 
assign cao = ~CAO;  //complement 
assign obi = ~OBI;  //complement 
assign oci = ~OCI;  //complement 
assign odi = ~ODI;  //complement 
assign baw = ~BAW;  //complement 
assign oaw = ~OAW;  //complement 
assign obw = ~OBW;  //complement 
assign TMC = ~tmc;  //complement 
assign TMD = ~tmd;  //complement 
assign dba = ~DBA;  //complement 
assign dbe = ~DBE;  //complement 
assign QFA = ~qfa;  //complement 
assign QFB = ~qfb;  //complement 
assign bay = ~BAY;  //complement 
assign oay = ~OAY;  //complement 
assign oby = ~OBY;  //complement 
assign dia = ~DIA;  //complement 
assign ola = ~OLA;  //complement 
assign qla = ~QLA;  //complement 
assign amc = ~AMC;  //complement 
assign oec = ~OEC;  //complement 
assign ofc = ~OFC;  //complement 
assign dib = ~DIB;  //complement 
assign olb = ~OLB;  //complement 
assign oma = ~OMA;  //complement 
assign qda = ~QDA;  //complement 
assign ami = ~AMI;  //complement 
assign oei = ~OEI;  //complement 
assign ofi = ~OFI;  //complement 
assign adi = ~ADI;  //complement 
assign aei = ~AEI;  //complement 
assign afi = ~AFI;  //complement 
assign aea = ~AEA;  //complement 
assign afa = ~AFA;  //complement 
assign ade = ~ADE;  //complement 
assign aee = ~AEE;  //complement 
assign afe = ~AFE;  //complement 
assign adb = ~ADB;  //complement 
assign aeb = ~AEB;  //complement 
assign afb = ~AFB;  //complement 
assign adf = ~ADF;  //complement 
assign aef = ~AEF;  //complement 
assign aff = ~AFF;  //complement 
assign qbj = ~QBJ;  //complement 
assign qcj = ~QCJ;  //complement 
assign NAB =  MAB & TQB  |  MCB & TRB  |  MEB & TSB  |  MGB & TTB  ; 
assign nab = ~NAB;  //complement 
assign oef = ~OEF;  //complement 
assign off = ~OFF;  //complement 
assign adj = ~ADJ;  //complement 
assign aej = ~AEJ;  //complement 
assign afj = ~AFJ;  //complement 
assign dbb = ~DBB;  //complement 
assign dbf = ~DBF;  //complement 
assign oih = ~OIH;  //complement 
assign bar = ~BAR;  //complement 
assign oar = ~OAR;  //complement 
assign obr = ~OBR;  //complement 
assign amn = ~AMN;  //complement 
assign oen = ~OEN;  //complement 
assign ofn = ~OFN;  //complement 
assign CAF =  BAP & TCB  |  AMF & TDB  ; 
assign caf = ~CAF;  //complement 
assign CAH =  BAR & TCB  |  AMH & TDB  ; 
assign cah = ~CAH;  //complement 
assign oab = ~OAB;  //complement 
assign obb = ~OBB;  //complement 
assign odb = ~ODB;  //complement 
assign bap = ~BAP;  //complement 
assign oap = ~OAP;  //complement 
assign obp = ~OBP;  //complement 
assign tbc = ~TBC;  //complement 
assign tbg = ~TBG;  //complement 
assign tpc = ~TPC;  //complement 
assign tuc = ~TUC;  //complement 
assign pcf = ~PCF;  //complement 
assign NBS =  MBS & TQS  |  MDS & TRS  |  MFS & TSS  |  MHS & TTS  ; 
assign nbs = ~NBS;  //complement 
assign NBL =  MBL & TQP  |  MDL & TRP  |  MFL & TSP  |  MHL & TTP  ; 
assign nbl = ~NBL;  //complement 
assign PAG = ~pag;  //complement 
assign PBC = ~pbc;  //complement 
assign PBS = ~pbs;  //complement 
assign FBA = ~fba;  //complement 
assign FCA = ~fca;  //complement 
assign EAC = ~eac;  //complement 
assign EBC = ~ebc;  //complement 
assign ECC = ~ecc;  //complement 
assign NBC =  MBC & TQK  |  MDC & TRK  |  MFC & TSK  |  MHC & TTK  ; 
assign nbc = ~NBC;  //complement 
assign FAJ =  QIB & FBA & EBF & EBG & EBH & EBI  ; 
assign faj = ~FAJ;  //complement  
assign FAI =  QIA & FBA & EBF & EBG & EBH  ; 
assign fai = ~FAI;  //complement  
assign FAG =  QIA & FBA & EBF  ; 
assign fag = ~FAG;  //complement 
assign EAG = ~eag;  //complement 
assign EBG = ~ebg;  //complement 
assign ECG = ~ecg;  //complement 
assign NAP =  MAP & TQH  |  MCP & TRH  |  MEP & TSH  |  MGP & TTH  ; 
assign nap = ~NAP;  //complement 
assign EAH = ~eah;  //complement 
assign EBH = ~ebh;  //complement 
assign ECH = ~ech;  //complement 
assign PAP = ~pap;  //complement 
assign PBL = ~pbl;  //complement 
assign EAD = ~ead;  //complement 
assign EBD = ~ebd;  //complement 
assign ECD = ~ecd;  //complement 
assign oag = ~OAG;  //complement 
assign obg = ~OBG;  //complement 
assign ocg = ~OCG;  //complement 
assign odg = ~ODG;  //complement 
assign ocw = ~OCW;  //complement 
assign odw = ~ODW;  //complement 
assign tia = ~TIA;  //complement 
assign tib = ~TIB;  //complement 
assign tma = ~TMA;  //complement 
assign tmb = ~TMB;  //complement 
assign dbc = ~DBC;  //complement 
assign dbg = ~DBG;  //complement 
assign oim = ~OIM;  //complement 
assign ocy = ~OCY;  //complement 
assign ody = ~ODY;  //complement 
assign dic = ~DIC;  //complement 
assign olc = ~OLC;  //complement 
assign ama = ~AMA;  //complement 
assign oea = ~OEA;  //complement 
assign ofa = ~OFA;  //complement 
assign NAG =  MAG & TQC  |  MCG & TRC  |  MEG & TSC  |  MGG & TTC  ; 
assign nag = ~NAG;  //complement 
assign did = ~DID;  //complement 
assign old = ~OLD;  //complement 
assign amg = ~AMG;  //complement 
assign oeg = ~OEG;  //complement 
assign ofg = ~OFG;  //complement 
assign adk = ~ADK;  //complement 
assign aek = ~AEK;  //complement 
assign afk = ~AFK;  //complement 
assign aml = ~AML;  //complement 
assign odp = ~ODP;  //complement 
assign adc = ~ADC;  //complement 
assign aec = ~AEC;  //complement 
assign afc = ~AFC;  //complement 
assign adg = ~ADG;  //complement 
assign aeg = ~AEG;  //complement 
assign afg = ~AFG;  //complement 
assign add = ~ADD;  //complement 
assign aed = ~AED;  //complement 
assign afd = ~AFD;  //complement 
assign adh = ~ADH;  //complement 
assign aeh = ~AEH;  //complement 
assign afh = ~AFH;  //complement 
assign FAL =  QIC & FCA & FBB & EBJ & EBK  ; 
assign fal = ~FAL;  //complement  
assign FAK =  QIC & FCA & FBB & EBJ  ; 
assign fak = ~FAK;  //complement 
assign EAL = ~eal;  //complement 
assign EBL = ~ebl;  //complement 
assign ECL = ~ecl;  //complement 
assign oel = ~OEL;  //complement 
assign ofl = ~OFL;  //complement 
assign adl = ~ADL;  //complement 
assign ael = ~AEL;  //complement 
assign afl = ~AFL;  //complement 
assign dbd = ~DBD;  //complement 
assign oif = ~OIF;  //complement 
assign dbh = ~DBH;  //complement 
assign ocr = ~OCR;  //complement 
assign odr = ~ODR;  //complement 
assign qqa = ~QQA;  //complement 
assign amp = ~AMP;  //complement 
assign oep = ~OEP;  //complement 
assign ofp = ~OFP;  //complement 
assign EAK = ~eak;  //complement 
assign EBK = ~ebk;  //complement 
assign ECK = ~eck;  //complement 
assign ocp = ~OCP;  //complement 
assign tbd = ~TBD;  //complement 
assign tbh = ~TBH;  //complement 
assign tpd = ~TPD;  //complement 
assign tud = ~TUD;  //complement 
assign bdm = ~BDM;  //complement 
assign EBB = ~ebb;  //complement 
assign pcg = ~PCG;  //complement 
assign NBR =  MBR & TQT  |  MDR & TRT  |  MFR & TST  |  MHR & TTT  ; 
assign nbr = ~NBR;  //complement 
assign pdc = ~PDC;  //complement 
assign pch = ~PCH;  //complement 
assign NBI =  MBI & TQO  |  MDI & TRO  |  MFI & TSO  |  MHI & TTO  ; 
assign nbi = ~NBI;  //complement 
assign bde = ~BDE;  //complement 
assign bce = ~BCE;  //complement 
assign bcm = ~BCM;  //complement 
assign bee = ~BEE;  //complement 
assign bem = ~BEM;  //complement 
assign PAM = ~pam;  //complement 
assign PBI = ~pbi;  //complement 
assign FAE =  QIA & EBA & EBB & EBC & EBD  ; 
assign fae = ~FAE;  //complement  
assign FAC =  QIA & EBA & EBB  ; 
assign fac = ~FAC;  //complement 
assign EAA = ~eaa;  //complement 
assign EBA = ~eba;  //complement 
assign ECA = ~eca;  //complement 
assign FAB =  QIB & EBA  ; 
assign fab = ~FAB;  //complement  
assign FAD =  QIB & EBA & EBB & EBC  ; 
assign fad = ~FAD;  //complement 
assign NAM =  MAM & TQG  |  MCM & TRG  |  MEM & TSG  |  MGM & TTG  ; 
assign nam = ~NAM;  //complement 
assign EAE = ~eae;  //complement 
assign EBE = ~ebe;  //complement 
assign ECE = ~ece;  //complement 
assign NBB =  MBB & TQL  |  MDB & TRL  |  MFB & TSL  |  MHB & TTL  ; 
assign nbb = ~NBB;  //complement 
assign EAF = ~eaf;  //complement 
assign EBF = ~ebf;  //complement 
assign ECF = ~ecf;  //complement 
assign PAF = ~paf;  //complement 
assign PBB = ~pbb;  //complement 
assign PBR = ~pbr;  //complement 
assign EAB = ~eab;  //complement 
assign ECB = ~ecb;  //complement 
assign bdd = ~BDD;  //complement 
assign bdj = ~BDJ;  //complement 
assign FAF =  QIB & EBA & EBB & EBC & EBD & EBE  ; 
assign faf = ~FAF;  //complement  
assign bcd = ~BCD;  //complement 
assign bcj = ~BCJ;  //complement 
assign bed = ~BED;  //complement 
assign bej = ~BEJ;  //complement 
assign CAC =  BAM & TCA  |  AMC & TDA  ; 
assign cac = ~CAC;  //complement 
assign CAI =  BAS & TCA  |  AMI & TDA  ; 
assign cai = ~CAI;  //complement 
assign EAI = ~eai;  //complement 
assign EBI = ~ebi;  //complement 
assign ECI = ~eci;  //complement 
assign bam = ~BAM;  //complement 
assign oam = ~OAM;  //complement 
assign obm = ~OBM;  //complement 
assign TNC = ~tnc;  //complement 
assign TND = ~tnd;  //complement 
assign DCA = ~dca;  //complement 
assign DCE = ~dce;  //complement 
assign oic = ~OIC;  //complement 
assign bas = ~BAS;  //complement 
assign oas = ~OAS;  //complement 
assign obs = ~OBS;  //complement 
assign BBE = ~bbe;  //complement 
assign BBM = ~bbm;  //complement 
assign die = ~DIE;  //complement 
assign ole = ~OLE;  //complement 
assign OGM = ~ogm;  //complement 
assign OHM = ~ohm;  //complement 
assign FBB = ~fbb;  //complement 
assign bal = ~BAL;  //complement 
assign OGE = ~oge;  //complement 
assign OHE = ~ohe;  //complement 
assign AGI = ~agi;  //complement 
assign AHI = ~ahi;  //complement 
assign AII = ~aii;  //complement 
assign AHA = ~aha;  //complement 
assign AIA = ~aia;  //complement 
assign AHE = ~ahe;  //complement 
assign AIE = ~aie;  //complement 
assign AGE = ~age;  //complement 
assign OHD = ~ohd;  //complement 
assign AGB = ~agb;  //complement 
assign AHB = ~ahb;  //complement 
assign AIB = ~aib;  //complement 
assign AGF = ~agf;  //complement 
assign AHF = ~ahf;  //complement 
assign AIF = ~aif;  //complement 
assign NAF =  MAF & TQD  |  MCF & TRD  |  MEF & TSD  |  MGF & TTD  ; 
assign naf = ~NAF;  //complement 
assign EAJ = ~eaj;  //complement 
assign EBJ = ~ebj;  //complement 
assign ECJ = ~ecj;  //complement 
assign OGJ = ~ogj;  //complement 
assign OHJ = ~ohj;  //complement 
assign AGJ = ~agj;  //complement 
assign AHJ = ~ahj;  //complement 
assign AIJ = ~aij;  //complement 
assign DCB = ~dcb;  //complement 
assign DCF = ~dcf;  //complement 
assign oil = ~OIL;  //complement 
assign bav = ~BAV;  //complement 
assign oav = ~OAV;  //complement 
assign obv = ~OBV;  //complement 
assign BBD = ~bbd;  //complement 
assign BBJ = ~bbj;  //complement 
assign dif = ~DIF;  //complement 
assign olf = ~OLF;  //complement 
assign OGD = ~ogd;  //complement 
assign CAB =  BAL & TCB  |  AMB & TDB  ; 
assign cab = ~CAB;  //complement 
assign CAL =  BAV & TCB  |  AML & TDB  ; 
assign cal = ~CAL;  //complement 
assign oaf = ~OAF;  //complement 
assign obf = ~OBF;  //complement 
assign ocf = ~OCF;  //complement 
assign odf = ~ODF;  //complement 
assign oal = ~OAL;  //complement 
assign obl = ~OBL;  //complement 
assign oka = ~OKA;  //complement 
assign pci = ~PCI;  //complement 
assign NBH =  MBH & TQN  |  MDH & TRN  |  MFH & TSN  |  MHH & TTN  ; 
assign nbh = ~NBH;  //complement 
assign pdb = ~PDB;  //complement 
assign pcj = ~PCJ;  //complement 
assign NBO =  MBO & TQQ  |  MDO & TRQ  |  MFO & TSQ  |  MHO & TTQ  ; 
assign nbo = ~NBO;  //complement 
assign bdk = ~BDK;  //complement 
assign bdo = ~BDO;  //complement 
assign bck = ~BCK;  //complement 
assign bco = ~BCO;  //complement 
assign bek = ~BEK;  //complement 
assign beo = ~BEO;  //complement 
assign qhc = ~QHC;  //complement 
assign qhd = ~QHD;  //complement 
assign PAC = ~pac;  //complement 
assign PAS = ~pas;  //complement 
assign PBO = ~pbo;  //complement 
assign qga = ~QGA;  //complement 
assign qgc = ~QGC;  //complement 
assign qge = ~QGE;  //complement 
assign NAS =  MAS & TQE  |  MCS & TRI  |  MES & TST  |  MGS & TTI  ; 
assign nas = ~NAS;  //complement 
assign qgb = ~QGB;  //complement 
assign qgd = ~QGD;  //complement 
assign qgf = ~QGF;  //complement 
assign NAL =  MAL & TQF  |  MCL & TRF  |  MEL & TSF  |  MGL & TTF  ; 
assign nal = ~NAL;  //complement 
assign PAL = ~pal;  //complement 
assign PBH = ~pbh;  //complement 
assign bfa = ~BFA;  //complement 
assign bfb = ~BFB;  //complement 
assign bfc = ~BFC;  //complement 
assign qmb = ~QMB;  //complement 
assign bdb = ~BDB;  //complement 
assign bdh = ~BDH;  //complement 
assign qma = ~QMA;  //complement 
assign bcb = ~BCB;  //complement 
assign bch = ~BCH;  //complement 
assign beb = ~BEB;  //complement 
assign beh = ~BEH;  //complement 
assign qha = ~QHA;  //complement 
assign qhb = ~QHB;  //complement 
assign oac = ~OAC;  //complement 
assign obc = ~OBC;  //complement 
assign occ = ~OCC;  //complement 
assign odc = ~ODC;  //complement 
assign ocm = ~OCM;  //complement 
assign odm = ~ODM;  //complement 
assign tja = ~TJA;  //complement 
assign tjb = ~TJB;  //complement 
assign tna = ~TNA;  //complement 
assign tnb = ~TNB;  //complement 
assign DCC = ~dcc;  //complement 
assign DCG = ~dcg;  //complement 
assign oii = ~OII;  //complement 
assign ocs = ~OCS;  //complement 
assign ods = ~ODS;  //complement 
assign BBK = ~bbk;  //complement 
assign BBO = ~bbo;  //complement 
assign dig = ~DIG;  //complement 
assign olg = ~OLG;  //complement 
assign OGO = ~ogo;  //complement 
assign OHO = ~oho;  //complement 
assign NAC =  MAC & TQA  |  MCC & TRA  |  MEC & TSA  |  MGC & TTA  ; 
assign nac = ~NAC;  //complement 
assign BBB = ~bbb;  //complement 
assign BBH = ~bbh;  //complement 
assign dih = ~DIH;  //complement 
assign olh = ~OLH;  //complement 
assign OGK = ~ogk;  //complement 
assign OHK = ~ohk;  //complement 
assign AGK = ~agk;  //complement 
assign AHK = ~ahk;  //complement 
assign AIK = ~aik;  //complement 
assign AGC = ~agc;  //complement 
assign AHC = ~ahc;  //complement 
assign AIC = ~aic;  //complement 
assign AGG = ~agg;  //complement 
assign AHG = ~ahg;  //complement 
assign AIG = ~aig;  //complement 
assign AGD = ~agd;  //complement 
assign AHD = ~ahd;  //complement 
assign AID = ~aid;  //complement 
assign AGH = ~agh;  //complement 
assign AHH = ~ahh;  //complement 
assign AIH = ~aih;  //complement 
assign OGH = ~ogh;  //complement 
assign OHH = ~ohh;  //complement 
assign AGL = ~agl;  //complement 
assign AHL = ~ahl;  //complement 
assign AIL = ~ail;  //complement 
assign DCD = ~dcd;  //complement 
assign DCH = ~dch;  //complement 
assign oib = ~OIB;  //complement 
assign tea = ~TEA;  //complement 
assign ocv = ~OCV;  //complement 
assign odv = ~ODV;  //complement 
assign OGB = ~ogb;  //complement 
assign OHB = ~ohb;  //complement 
assign qna = ~QNA;  //complement 
assign qnb = ~QNB;  //complement 
assign qnc = ~QNC;  //complement 
assign qnd = ~QND;  //complement 
assign tec = ~TEC;  //complement 
assign ted = ~TED;  //complement 
assign ocl = ~OCL;  //complement 
assign odl = ~ODL;  //complement 
assign okb = ~OKB;  //complement 
assign okc = ~OKC;  //complement 
assign peb = ~PEB;  //complement 
assign pck = ~PCK;  //complement 
assign NBQ =  MBQ & TQS  |  MDQ & TRS  |  MFQ & TSS  |  MHQ & TTS  ; 
assign nbq = ~NBQ;  //complement 
assign TQQ = ~tqq;  //complement 
assign TRQ = ~trq;  //complement 
assign TSQ = ~tsq;  //complement 
assign TTQ = ~ttq;  //complement 
assign NBJ =  MBJ & TQP  |  MDJ & TRP  |  MFJ & TSP  |  MHJ & TTP  ; 
assign nbj = ~NBJ;  //complement 
assign tqn = ~TQN;  //complement 
assign trn = ~TRN;  //complement 
assign tsn = ~TSN;  //complement 
assign ttn = ~TTN;  //complement 
assign bdc = ~BDC;  //complement 
assign bdi = ~BDI;  //complement 
assign bcc = ~BCC;  //complement 
assign bci = ~BCI;  //complement 
assign bec = ~BEC;  //complement 
assign bei = ~BEI;  //complement 
assign PAE = ~pae;  //complement 
assign PBA = ~pba;  //complement 
assign PBQ = ~pbq;  //complement 
assign QHK = ~qhk;  //complement 
assign QHL = ~qhl;  //complement 
assign QHG = ~qhg;  //complement 
assign QHH = ~qhh;  //complement 
assign NBA =  MBA & TQK  |  MDA & TRK  |  MFA & TSK  |  MHA & TTK  ; 
assign nba = ~NBA;  //complement 
assign TQI = ~tqi;  //complement 
assign TRI = ~trii;  //complement 
assign TSI = ~tsi;  //complement 
assign TTI = ~tti;  //complement 
assign amf = ~AMF;  //complement 
assign NAN =  MAN & TQH  |  MCN & TRH  |  MEN & TSH  |  MGN & TTH  ; 
assign nan = ~NAN;  //complement 
assign tqf = ~TQF;  //complement 
assign trf = ~TRF;  //complement 
assign tsf = ~TSF;  //complement 
assign ttf = ~TTF;  //complement 
assign PAN = ~pan;  //complement 
assign PBJ = ~pbj;  //complement 
assign oli = ~OLI;  //complement 
assign QMC = ~qmc;  //complement 
assign QMD = ~qmd;  //complement 
assign bdf = ~BDF;  //complement 
assign bdn = ~BDN;  //complement 
assign bcf = ~BCF;  //complement 
assign bcn = ~BCN;  //complement 
assign bef = ~BEF;  //complement 
assign ben = ~BEN;  //complement 
assign CAA =  BAK & TCA  |  AMA & TDA  ; 
assign caa = ~CAA;  //complement 
assign CAK =  BAU & TCA  |  AMK & TDA  ; 
assign cak = ~CAK;  //complement 
assign oae = ~OAE;  //complement 
assign obe = ~OBE;  //complement 
assign oce = ~OCE;  //complement 
assign ode = ~ODE;  //complement 
assign bak = ~BAK;  //complement 
assign oak = ~OAK;  //complement 
assign obk = ~OBK;  //complement 
assign TOC = ~toc;  //complement 
assign TOD = ~tod;  //complement 
assign DDA = ~dda;  //complement 
assign DDE = ~dde;  //complement 
assign oik = ~OIK;  //complement 
assign bau = ~BAU;  //complement 
assign oau = ~OAU;  //complement 
assign obu = ~OBU;  //complement 
assign BBC = ~bbc;  //complement 
assign BBI = ~bbi;  //complement 
assign OJA = ~oja;  //complement 
assign qra = ~QRA;  //complement 
assign OGC = ~ogc;  //complement 
assign OHC = ~ohc;  //complement 
assign NAE =  MAE & TQC  |  MCE & TRC  |  MEE & TSC  |  MGE & TTC  ; 
assign nae = ~NAE;  //complement 
assign obn = ~OBN;  //complement 
assign OGI = ~ogi;  //complement 
assign OHI = ~ohi;  //complement 
assign AJI = ~aji;  //complement 
assign AKI = ~aki;  //complement 
assign ALI = ~ali;  //complement 
assign AKA = ~aka;  //complement 
assign ALA = ~ala;  //complement 
assign AJE = ~aje;  //complement 
assign AKE = ~ake;  //complement 
assign ALE = ~ale;  //complement 
assign AJB = ~ajb;  //complement 
assign AKB = ~akb;  //complement 
assign ALB = ~alb;  //complement 
assign AJF = ~ajf;  //complement 
assign AKF = ~akf;  //complement 
assign ALF = ~alf;  //complement 
assign TQA = ~tqa;  //complement 
assign TRA = ~tra;  //complement 
assign TSA = ~tsa;  //complement 
assign TTA = ~tta;  //complement 
assign BBF = ~bbf;  //complement 
assign BBN = ~bbn;  //complement 
assign teb = ~TEB;  //complement 
assign tee = ~TEE;  //complement 
assign OGF = ~ogf;  //complement 
assign OHF = ~ohf;  //complement 
assign AJJ = ~ajj;  //complement 
assign AKJ = ~akj;  //complement 
assign ALJ = ~alj;  //complement 
assign DDB = ~ddb;  //complement 
assign DDF = ~ddf;  //complement 
assign oid = ~OID;  //complement 
assign bat = ~BAT;  //complement 
assign oat = ~OAT;  //complement 
assign obt = ~OBT;  //complement 
assign CAD =  BAN & TCB  |  AMD & TDB  ; 
assign cad = ~CAD;  //complement 
assign OGN = ~ogn;  //complement 
assign OHN = ~ohn;  //complement 
assign CAJ =  BAT & TCB  |  AMJ & TDB  ; 
assign caj = ~CAJ;  //complement 
assign qne = ~QNE;  //complement 
assign qng = ~QNG;  //complement 
assign ban = ~BAN;  //complement 
assign oan = ~OAN;  //complement 
assign okd = ~OKD;  //complement 
assign oke = ~OKE;  //complement 
assign NBP =  MBP & TQR  |  MDP & TRR  |  MFP & TSR  |  MHP & TTR  ; 
assign nbp = ~NBP;  //complement 
assign tqp = ~TQP;  //complement 
assign tsp = ~TSP;  //complement 
assign ttp = ~TTP;  //complement 
assign pcl = ~PCL;  //complement 
assign pda = ~PDA;  //complement 
assign pcm = ~PCM;  //complement 
assign pcn = ~PCN;  //complement 
assign TQS = ~tqs;  //complement 
assign TRS = ~trs;  //complement 
assign TSS = ~tss;  //complement 
assign TTS = ~tts;  //complement 
assign trp = ~TRP;  //complement 
assign NBG =  MBG & TQM  |  MDG & TRM  |  MFG & TSM  |  MHG & TTM  ; 
assign nbg = ~NBG;  //complement 
assign bda = ~BDA;  //complement 
assign bdg = ~BDG;  //complement 
assign bca = ~BCA;  //complement 
assign bcg = ~BCG;  //complement 
assign bea = ~BEA;  //complement 
assign beg = ~BEG;  //complement 
assign PAK = ~pak;  //complement 
assign PBG = ~pbg;  //complement 
assign TQK = ~tqk;  //complement 
assign QHS = ~qhs;  //complement 
assign QHT = ~qht;  //complement 
assign QHO = ~qho;  //complement 
assign QHP = ~qhp;  //complement 
assign TRK = ~trk;  //complement 
assign TSK = ~tsk;  //complement 
assign TTK = ~ttk;  //complement 
assign TQG = ~tqg;  //complement 
assign TRG = ~trg;  //complement 
assign TSG = ~tsg;  //complement 
assign TTG = ~ttg;  //complement 
assign NAK =  MAK & TQE  |  MCK & TRE  |  MEK & TSE  |  MGK & TTE  ; 
assign nak = ~NAK;  //complement 
assign wbe = ~WBE;  //complement 
assign wbf = ~WBF;  //complement 
assign wbg = ~WBG;  //complement 
assign wbh = ~WBH;  //complement 
assign wca = ~WCA;  //complement 
assign wcb = ~WCB;  //complement 
assign wcc = ~WCC;  //complement 
assign wcd = ~WCD;  //complement 
assign wce = ~WCE;  //complement 
assign wcf = ~WCF;  //complement 
assign wcg = ~WCG;  //complement 
assign wch = ~WCH;  //complement 
assign NAT =  MAT & TQJ  |  MCT & TRJ  |  MET & TSJ  |  MGT & TTJ  ; 
assign nat = ~NAT;  //complement 
assign wba = ~WBA;  //complement 
assign wbb = ~WBB;  //complement 
assign wbc = ~WBC;  //complement 
assign wbd = ~WBD;  //complement 
assign PAD = ~pad;  //complement 
assign PAT = ~pat;  //complement 
assign PBP = ~pbp;  //complement 
assign qme = ~QME;  //complement 
assign bdl = ~BDL;  //complement 
assign bdp = ~BDP;  //complement 
assign qmf = ~QMF;  //complement 
assign bcl = ~BCL;  //complement 
assign bcp = ~BCP;  //complement 
assign bel = ~BEL;  //complement 
assign bep = ~BEP;  //complement 
assign ock = ~OCK;  //complement 
assign odk = ~ODK;  //complement 
assign tka = ~TKA;  //complement 
assign tkb = ~TKB;  //complement 
assign toa = ~TOA;  //complement 
assign tob = ~TOB;  //complement 
assign DDC = ~ddc;  //complement 
assign DDG = ~ddg;  //complement 
assign oia = ~OIA;  //complement 
assign ocu = ~OCU;  //complement 
assign odu = ~ODU;  //complement 
assign BBA = ~bba;  //complement 
assign BBG = ~bbg;  //complement 
assign OGA = ~oga;  //complement 
assign OHA = ~oha;  //complement 
assign BBL = ~bbl;  //complement 
assign BBP = ~bbp;  //complement 
assign TGE = ~tge;  //complement 
assign FAH =  QIB & FBA & EBF & EBG  ; 
assign fah = ~FAH;  //complement  
assign OGG = ~ogg;  //complement 
assign OHG = ~ohg;  //complement 
assign AJK = ~ajk;  //complement 
assign AKK = ~akk;  //complement 
assign ALK = ~alk;  //complement 
assign OGL = ~ogl;  //complement 
assign AJC = ~ajc;  //complement 
assign AKC = ~akc;  //complement 
assign ALC = ~alc;  //complement 
assign AJG = ~ajg;  //complement 
assign AKG = ~akg;  //complement 
assign ALG = ~alg;  //complement 
assign TGF = ~tgf;  //complement 
assign TGG = ~tgg;  //complement 
assign TGH = ~tgh;  //complement 
assign AJD = ~ajd;  //complement 
assign AKD = ~akd;  //complement 
assign ALD = ~ald;  //complement 
assign AJH = ~ajh;  //complement 
assign AKH = ~akh;  //complement 
assign ALH = ~alh;  //complement 
assign tqd = ~TQD;  //complement 
assign trd = ~TRD;  //complement 
assign tsd = ~TSD;  //complement 
assign ttd = ~TTD;  //complement 
assign NAD =  MAD & TQB  |  MCD & TRB  |  MED & TSB  |  MGD & TTB  ; 
assign nad = ~NAD;  //complement 
assign OHL = ~ohl;  //complement 
assign AJL = ~ajl;  //complement 
assign AKL = ~akl;  //complement 
assign ALL = ~all;  //complement 
assign DDD = ~ddd;  //complement 
assign DDH = ~ddh;  //complement 
assign oij = ~OIJ;  //complement 
assign oct = ~OCT;  //complement 
assign odt = ~ODT;  //complement 
assign OGP = ~ogp;  //complement 
assign OHP = ~ohp;  //complement 
assign qnf = ~QNF;  //complement 
assign oad = ~OAD;  //complement 
assign obd = ~OBD;  //complement 
assign ocd = ~OCD;  //complement 
assign odd = ~ODD;  //complement 
assign ocn = ~OCN;  //complement 
assign odn = ~ODN;  //complement 
assign okf = ~OKF;  //complement 
assign okg = ~OKG;  //complement 
assign iaa = ~IAA; //complement 
assign iab = ~IAB; //complement 
assign iac = ~IAC; //complement 
assign iad = ~IAD; //complement 
assign iae = ~IAE; //complement 
assign iaf = ~IAF; //complement 
assign iag = ~IAG; //complement 
assign iah = ~IAH; //complement 
assign iai = ~IAI; //complement 
assign iaj = ~IAJ; //complement 
assign iak = ~IAK; //complement 
assign ial = ~IAL; //complement 
assign iam = ~IAM; //complement 
assign ian = ~IAN; //complement 
assign iao = ~IAO; //complement 
assign iap = ~IAP; //complement 
assign ica = ~ICA; //complement 
assign icb = ~ICB; //complement 
assign icc = ~ICC; //complement 
assign icd = ~ICD; //complement 
assign ice = ~ICE; //complement 
assign icf = ~ICF; //complement 
assign icg = ~ICG; //complement 
assign ich = ~ICH; //complement 
assign ici = ~ICI; //complement 
assign icj = ~ICJ; //complement 
assign ick = ~ICK; //complement 
assign icl = ~ICL; //complement 
assign icm = ~ICM; //complement 
assign icn = ~ICN; //complement 
assign ico = ~ICO; //complement 
assign icp = ~ICP; //complement 
assign iga = ~IGA; //complement 
assign ija = ~IJA; //complement 
assign ika = ~IKA; //complement 
assign ila = ~ILA; //complement 
assign ilb = ~ILB; //complement 
assign ilc = ~ILC; //complement 
assign ild = ~ILD; //complement 
assign ile = ~ILE; //complement 
assign ilf = ~ILF; //complement 
assign ilg = ~ILG; //complement 
assign ilh = ~ILH; //complement 
assign ili = ~ILI; //complement 
assign ipa = ~IPA; //complement 
assign ipb = ~IPB; //complement 
assign iqa = ~IQA; //complement 
assign iqb = ~IQB; //complement 
assign iqc = ~IQC; //complement 
assign ira = ~IRA; //complement 
assign irb = ~IRB; //complement 
assign isa = ~ISA; //complement 
always@(posedge IZZ )
   begin 
 WDE <= QEA & QBD ; 
 WDF <= QEA & QBD ; 
 WDG <= QEA & QBD ; 
 WDH <= QEA & QBD ; 
 TQT <= QHE ; 
 TRT <= QHI ; 
 TST <= QHM ; 
 TTT <= QHQ ; 
 WEA <= QEA & QBB ; 
 WEB <= QEA & QBB ; 
 WEC <= QEA & QBB ; 
 WED <= QEA & QBB ; 
 WDA <= QEA & QBD ; 
 WDB <= QEA & QBD ; 
 WDC <= QEA & QBD ; 
 WDD <= QEA & QBD ; 
 PCA <=  PBM & paq & paa  |  pbm & PAQ & paa  |  pbm & paq & PAA  |  PBM & PAQ & PAA  ;
 PDF <= PCA ; 
 WEE <= QEA & QBB ; 
 WEF <= QEA & QBB ; 
 WEG <= QEA & QBB ; 
 WEH <= QEA & QBB ; 
 tqo <= qhe ; 
 tro <= qhi ; 
 tso <= qhm ; 
 tto <= qhq ; 
 paa <= naa ; 
 paq <= naq ; 
 pbm <= nbm ; 
 qhi <=  qgc  |  QGD  |  qja  ; 
 qhj <=  qgc  |  QGD  |  qja  ; 
 qhe <=  QGC  |  QGD  |  qja  ; 
 qhf <=  QGC  |  QGD  |  qja  ; 
 TQL <= QHE ; 
 TRL <= QHI ; 
 TSL <= QHM ; 
 TTL <= QHQ ; 
 TQH <= QHE ; 
 TRH <= QHI ; 
 TSH <= QHM ; 
 TTH <= QHQ ; 
 paj <= naj ; 
 pbf <= nbf ; 
 OAA <= NAA ; 
 OBA <= NAA ; 
 OCA <= NAA ; 
 ODA <= NAA ; 
 BAO <=  NAO  |  IAE & TBA  |  CAE  ; 
 OAO <=  NAO  |  IAE & TBA  |  CAE  ; 
 OBO <=  NAO  |  IAE & TBA  |  CAE  ; 
 tlc <=  qha  |  QFB  |  ira  ; 
 tld <=  qha  |  QFB  |  IRA  ; 
 DAA <= DIA ; 
 DAE <= DIE ; 
 OIG <= NBM ; 
 trc <= qhi ; 
 BAQ <=  NAQ  |  IAG & TBA  |  CAG  ; 
 OAQ <=  NAQ  |  IAG & TBA  |  CAG  ; 
 OBQ <=  NAQ  |  IAG & TBA  |  CAG  ; 
 TGA <= QFA ; 
 TGB <= QFA ; 
 TGC <= QFA ; 
 TGD <= QFA ; 
 AMM <=  ICM & TPA  |  BEM & TUA  ; 
 OEM <=  ICM & TPA  |  BEM & TUA  ; 
 OFM <=  ICM & TPA  |  BEM & TUA  ; 
 tqc <= qhe ; 
 tsc <= qhm ; 
 ttc <= qhq ; 
 AME <=  ICE & TPA  |  BEE & TUA  ; 
 OEE <=  ICE & TPA  |  BEE & TUA  ; 
 OFE <=  ICE & TPA  |  BEE & TUA  ; 
 AAI <=  ICM & TLA  |  AAI & THA  |  ECI & TGA  ; 
 ABI <=  ICM & TLA  |  AAI & THA  |  ECI & TGA  ; 
 ACI <=  ICM & TLA  |  AAI & THA  |  ECI & TGA  ; 
 AMJ <=  ICJ & TPA  |  BEJ & TUA  ; 
 ABA <=  ICE & TLC  |  IGA & TLD  |  ABA & THA  |  ECA & TGA  ; 
 ACA <=  ICE & TLC  |  IGA & TLD  |  ABA & THA  |  ECA & TGA  ; 
 AAE <=  ICI & TLA  |  AAE & THA  |  ECE & TGA  ; 
 ABE <=  ICI & TLA  |  AAE & THA  |  ECE & TGA  ; 
 ACE <=  ICI & TLA  |  AAE & THA  |  ECE & TGA  ; 
 AAA <=  ICE & TLC  |  IGA & TLD  |  AAA & THA  |  ECA & TGA  ; 
 AAB <=  ICF & TLA  |  AAB & THA  |  ECB & TGA  ; 
 ABB <=  ICF & TLA  |  AAB & THA  |  ECB & TGA  ; 
 ACB <=  ICF & TLA  |  AAB & THA  |  ECB & TGA  ; 
 AAF <=  ICJ & TLA  |  AAF & THA  |  ECF & TGA  ; 
 ABF <=  ICJ & TLA  |  AAF & THA  |  ECF & TGA  ; 
 ACF <=  ICJ & TLA  |  AAF & THA  |  ECF & TGA  ; 
 WAA <= QEA & QBJ ; 
 WAB <= QEA & QBJ ; 
 WAC <= QEA & QBJ ; 
 WAD <= QEA & QBJ ; 
 WAE <= QEA & QBJ ; 
 WAF <= QEA & QBJ ; 
 WAG <= QEA & QBJ ; 
 WAH <= QEA & QBJ ; 
 OEJ <=  ICJ & TPA  |  BEJ & TUA  ; 
 OFJ <=  ICJ & TPA  |  BEJ & TUA  ; 
 AAJ <=  ICN & TLA  |  AAJ & THA  |  ECJ & TGA  ; 
 ABJ <=  ICN & TLA  |  AAJ & THA  |  ECJ & TGA  ; 
 ACJ <=  ICN & TLA  |  AAJ & THA  |  ECJ & TGA  ; 
 DAB <= DIB ; 
 DAF <= DIF ; 
 BAZ <=  NBF  |  IAP & TBA  |  CAP  ; 
 OAZ <=  NBF  |  IAP & TBA  |  CAP  ; 
 OBZ <=  NBF  |  IAP & TBA  |  CAP  ; 
 QPA <= IPA ; 
 QPB <= IPB ; 
 AMD <=  ICD & TPA  |  BED & TUA  ; 
 OED <=  ICD & TPA  |  BED & TUA  ; 
 OFD <=  ICD & TPA  |  BED & TUA  ; 
 OAJ <= NAJ ; 
 OBJ <= NAJ ; 
 OCJ <= NAJ ; 
 ODJ <= NAJ ; 
 BAX <=  NBD  |  IAN & TBA  |  CAN  ; 
 OAX <=  NBD  |  IAN & TBA  |  CAN  ; 
 OBX <=  NBD  |  IAN & TBA  |  CAN  ; 
 TBA <= QQA ; 
 TBE <= QQA ; 
 TPA <= QPA ; 
 TUA <= QPB ; 
 PCB <=  PBT & pah & pbd  |  pbt & PAH & pbd  |  pbt & pah & PBD  |  PBT & PAH & PBD  ;
 PEA <=  PDD & pde & pdf  |  pdd & PDE & pdf  |  pdd & pde & PDF  |  PDD & PDE & PDF  ;
 PCC <=  PBK & pao & pbf  |  pbk & PAO & pbf  |  pbk & pao & PBF  |  PBK & PAO & PBF  ;
 PDE <= PCB ; 
 TQR <= QHF ; 
 TRR <= QHJ ; 
 TSR <= QHN ; 
 TTR <= QHR ; 
 tqm <= qhf ; 
 trm <= qhj ; 
 tsm <= qhn ; 
 ttm <= qhr ; 
 OAI <= NAI ; 
 pao <= nao ; 
 pbk <= nbk ; 
 qhq <=  qgc  |  qgd  |  qja  ; 
 qhr <=  qgc  |  qgd  |  qja  ; 
 qhm <=  QGC  |  qgd  |  qja  ; 
 qhn <=  QGC  |  qgd  |  qja  ; 
 tqe <= qhf ; 
 tre <= qhj ; 
 tse <= qhn ; 
 tte <= qhr ; 
 TTJ <= QHR ; 
 TQJ <= QHF ; 
 TRJ <= QHJ ; 
 TSJ <= QHN ; 
 pah <= nah ; 
 pbd <= nbd ; 
 pbt <= nbt ; 
 OCB <= NAB ; 
 QJA <= IJA ; 
 QJB <= IJA ; 
 TCA <= QQB ; 
 TDA <= QQC ; 
 ONA <=  PEA & peb  |  pea & PEB  ; 
 OCO <=  NAO  |  IAE & TBB  |  CAE  ; 
 ODO <=  NAO  |  IAE & TBB  |  CAE  ; 
 THA <= qfb & qha ; 
 THB <= qfb & qha ; 
 TLA <= qfb & QHA ; 
 TLB <= qfb & QHA ; 
 DAC <= DIC ; 
 DAG <= DIG ; 
 OIE <= NBK ; 
 OCQ <=  NAQ  |  IAG & TBB  |  CAG  ; 
 ODQ <=  NAQ  |  IAG & TBB  |  CAG  ; 
 AMO <=  ICO & TPB  |  BEO & TUB  ; 
 OEO <=  ICO & TPB  |  BEO & TUB  ; 
 OFO <=  ICO & TPB  |  BEO & TUB  ; 
 QQC <= IQC ; 
 ODX <=  NBD  |  IAN & TBB  |  CAN  ; 
 AMK <=  ICK & TPB  |  BEK & TUB  ; 
 OEK <=  ICK & TPB  |  BEK & TUB  ; 
 OFK <=  ICK & TPB  |  BEK & TUB  ; 
 AAK <=  ICO & TLB  |  AAK & THB  |  ECK & TGB  ; 
 ABK <=  ICO & TLB  |  AAK & THB  |  ECK & TGB  ; 
 ACK <=  ICO & TLB  |  AAK & THB  |  ECK & TGB  ; 
 AAC <=  ICG & TLB  |  AAC & THB  |  ECC & TGB  ; 
 ABC <=  ICG & TLB  |  AAC & THB  |  ECC & TGB  ; 
 ACC <=  ICG & TLB  |  AAC & THB  |  ECC & TGB  ; 
 AAG <=  ICK & TLB  |  AAG & THB  |  ECG & TGB  ; 
 ABG <=  ICK & TLB  |  AAG & THB  |  ECG & TGB  ; 
 ACG <=  ICK & TLB  |  AAG & THB  |  ECG & TGB  ; 
 AAD <=  ICH & TLB  |  AAD & THB  |  ECD & TGB  ; 
 ABD <=  ICH & TLB  |  AAD & THB  |  ECD & TGB  ; 
 ACD <=  ICH & TLB  |  AAD & THB  |  ECD & TGB  ; 
 AAH <=  ICL & TLB  |  AAH & THB  |  ECH & TGB  ; 
 ABH <=  ICL & TLB  |  AAH & THB  |  ECH & TGB  ; 
 ACH <=  ICL & TLB  |  AAH & THB  |  ECH & TGB  ; 
 TQB <= QHF ; 
 TRB <= QHJ ; 
 TSB <= QHM ; 
 TTB <= QHR ; 
 AMH <=  ICH & TPB  |  BEH & TUB  ; 
 OEH <=  ICH & TPB  |  BEH & TUB  ; 
 OFH <=  ICH & TPB  |  BEH & TUB  ; 
 AAL <=  QRA & TLB  |  AAL & THB  |  ECL & TGB  ; 
 ABL <=  QRA & TLB  |  AAL & THB  |  ECL & TGB  ; 
 ACL <=  QRA & TLB  |  AAL & THB  |  ECL & TGB  ; 
 DAD <= DID ; 
 DAH <= DIH ; 
 OCZ <=  NBF  |  IAP & TBB  |  CAP  ; 
 ODZ <=  NBF  |  IAP & TBB  |  CAP  ; 
 QQB <= IQB ; 
 AMB <=  ICB & TPB  |  BEB & TUB  ; 
 OEB <=  ICB & TPB  |  BEB & TUB  ; 
 OFB <=  ICB & TPB  |  BEB & TUB  ; 
 TCB <= QQB ; 
 TDB <= QQC ; 
 OAH <= NAH ; 
 OBH <= NAH ; 
 OCH <= NAH ; 
 ODH <= NAH ; 
 OCX <=  NBD  |  IAN & TBB  |  CAN  ; 
 TBB <= QQA ; 
 TBF <= QQA ; 
 TPB <= QPA ; 
 TUB <= QPB ; 
 QBB <=  QBA  |  QCB & qbc  |  QDF  ; 
 QCB <=  QBA  |  QCB & qbc  |  QDF  ; 
 QDC <= QDB ; 
 QDE <= QDD ; 
 QEA <=  QAD  |  QAE  |  QAF  |  QAG  ; 
 QEB <=  QAD  |  QAE  |  QAF  |  QAG  ; 
 QDD <= QDC ; 
 QBD <=  QCD & qbe & qdj  |  QBC  ; 
 QCD <=  QCD & qbe & qdj  |  QBC  ; 
 PDD <=  PCE & pcd & pcc  |  pce & PCD & pcc  |  pce & pcd & PCC  |  PCE & PCD & PCC  ;
 PCE <=  PAJ & pbe & pai  |  paj & PBE & pai  |  paj & pbe & PAI  |  PAJ & PBE & PAI  ;
 PCD <=  PBN & par & pab  |  pbn & PAR & pab  |  pbn & par & PAB  |  PBN & PAR & PAB  ;
 pab <= nab ; 
 par <= nar ; 
 pbn <= nbn ; 
 pai <= nai ; 
 pbe <= nbe ; 
 QAE <= qdi & QAD ; 
 QAG <= qdi & QAF ; 
 QBG <= QAI & QCF ; 
 QBI <= QAI & QCH ; 
 qia <= qba ; 
 qib <= qba ; 
 qic <= qba ; 
 QBF <=  QCF & qbg & qdj  |  QBE  ; 
 QCF <=  QCF & qbg & qdj  |  QBE  ; 
 QBH <=  QCH & qbi & qdj  |  QBG  ; 
 QCH <=  QCH & qbi & qdj  |  QBG  ; 
 QBA <= QAI & QCJ ; 
 QBC <= QAI & QCB ; 
 QBE <= QAI & QCD ; 
 QDB <= QDA ; 
 QAA <= QDA & QLA ; 
 QDI <= QDA & qde ; 
 QDJ <= QDA & qde ; 
 QAC <= qdi & QAB ; 
 QAI <= qdi & QAH ; 
 QAB <= qdi & QAA ; 
 QAD <= qdi & QAC ; 
 QAF <= qdi & QAE ; 
 QAH <= qdi & QAG ; 
 QDF <= qde & QDD ; 
 QDG <= qde & QDD ; 
 QDH <= qde & QDD ; 
 OBI <= NAI ; 
 OCI <= NAI ; 
 ODI <= NAI ; 
 BAW <=  NBC  |  IAM & TBC  |  CAM  ; 
 OAW <=  NBC  |  IAM & TBC  |  CAM  ; 
 OBW <=  NBC  |  IAM & TBC  |  CAM  ; 
 tmc <=  qhb  |  QFB  |  ira  ; 
 tmd <=  qhb  |  QFB  |  IRA  ; 
 DBA <= DIA ; 
 DBE <= DIE ; 
 qfa <= qda ; 
 qfb <= qda ; 
 BAY <=  NBE  |  IAO & TBC  |  CAO  ; 
 OAY <=  NBE  |  IAO & TBC  |  CAO  ; 
 OBY <=  NBE  |  IAO & TBC  |  CAO  ; 
 DIA <= ILA ; 
 OLA <= ILA ; 
 QLA <= ILI ; 
 AMC <=  ICC & TPC  |  BEC & TUC  ; 
 OEC <=  ICC & TPC  |  BEC & TUC  ; 
 OFC <=  ICC & TPC  |  BEC & TUC  ; 
 DIB <= ILB ; 
 OLB <= ILB ; 
 OMA <= IKA ; 
 QDA <= IKA ; 
 AMI <=  ICI & TPC  |  BEI & TUC  ; 
 OEI <=  ICI & TPC  |  BEI & TUC  ; 
 OFI <=  ICI & TPC  |  BEI & TUC  ; 
 ADI <=  ICM & TMA  |  ADI & TIA  |  ECI & TGC  ; 
 AEI <=  ICM & TMA  |  ADI & TIA  |  ECI & TGC  ; 
 AFI <=  ICM & TMA  |  ADI & TIA  |  ECI & TGC  ; 
 AEA <=  ICE & TMC  |  IGA & TMD  |  AEA & TIA  |  ECA & TGC  ; 
 AFA <=  ICE & TMC  |  IGA & TMD  |  AEA & TIA  |  ECA & TGC  ; 
 ADE <=  ICI & TMA  |  ADE & TIA  |  ECE & TGC  ; 
 AEE <=  ICI & TMA  |  ADE & TIA  |  ECE & TGC  ; 
 AFE <=  ICI & TMA  |  ADE & TIA  |  ECE & TGC  ; 
 ADB <=  ICF & TMA  |  ADB & TIA  |  ECB & TGC  ; 
 AEB <=  ICF & TMA  |  ADB & TIA  |  ECB & TGC  ; 
 AFB <=  ICF & TMA  |  ADB & TIA  |  ECB & TGC  ; 
 ADF <=  ICJ & TMA  |  ADF & TIA  |  ECF & TGC  ; 
 AEF <=  ICJ & TMA  |  ADF & TIA  |  ECF & TGC  ; 
 AFF <=  ICJ & TMA  |  ADF & TIA  |  ECF & TGC  ; 
 QBJ <=  QCJ & qba & qdj  |  QBI  ; 
 QCJ <=  QCJ & qba & qdj  |  QBI  ; 
 OEF <=  ICF & TPC  |  BEF & TUC  ; 
 OFF <=  ICF & TPC  |  BEF & TUC  ; 
 ADJ <=  ICN & TMA  |  ADJ & TIA  |  ECJ & TGC  ; 
 AEJ <=  ICN & TMA  |  ADJ & TIA  |  ECJ & TGC  ; 
 AFJ <=  ICN & TMA  |  ADJ & TIA  |  ECJ & TGC  ; 
 DBB <= DIB ; 
 DBF <= DIF ; 
 OIH <= MBN ; 
 BAR <=  NAR  |  IAH & TBC  |  CAH  ; 
 OAR <=  NAR  |  IAH & TBC  |  CAH  ; 
 OBR <=  NAR  |  IAH & TBC  |  CAH  ; 
 AMN <=  ICN & TPC  |  BEN & TUC  ; 
 OEN <=  ICN & TPC  |  BEN & TUC  ; 
 OFN <=  ICN & TPC  |  BEN & TUC  ; 
 OAB <= NAB ; 
 OBB <= NAB ; 
 ODB <= NAB ; 
 BAP <=  NAP  |  IAF & TBC  |  CAF  ; 
 OAP <=  NAP  |  IAF & TBC  |  CAF  ; 
 OBP <=  NAP  |  IAF & TBC  |  CAF  ; 
 TBC <= QQA ; 
 TBG <= QQA ; 
 TPC <= QPA ; 
 TUC <= QPB ; 
 PCF <=  PBS & pbc & pag  |  pbs & PBC & pag  |  pbs & pbc & PAG  |  PBS & PBC & PAG  ;
 pag <= nag ; 
 pbc <= nbc ; 
 pbs <= nbs ; 
 fba <=  eaa  |  eab  |  eac  |  ead  |  eae  ; 
 fca <=  eaa  |  eab  |  eac  |  ead  |  eae  ; 
 eac <=  EAC & FAC  |  eac & fac  |  QDG  ; 
 ebc <=  EAC & FAC  |  eac & fac  |  QDG  ; 
 ecc <=  EAC & FAC  |  eac & fac  |  QDG  ; 
 eag <=  EAG & FAG  |  eag & fag  |  QDG  ; 
 ebg <=  EAG & FAG  |  eag & fag  |  QDG  ; 
 ecg <=  EAG & FAG  |  eag & fag  |  QDG  ; 
 eah <=  EAH & FAH  |  eah & fah  |  QDG  ; 
 ebh <=  EAH & FAH  |  eah & fah  |  QDG  ; 
 ech <=  EAH & FAH  |  eah & fah  |  QDG  ; 
 pap <= nap ; 
 pbl <= nbl ; 
 ead <=  EAD & FAD  |  ead & fad  |  QDG  ; 
 ebd <=  EAD & FAD  |  ead & fad  |  QDG  ; 
 ecd <=  EAD & FAD  |  ead & fad  |  QDG  ; 
 OAG <= NAG ; 
 OBG <= NAG ; 
 OCG <= NAG ; 
 ODG <= NAG ; 
 OCW <=  NBC  |  IAM & TBD  |  CAM  ; 
 ODW <=  NBC  |  IAM & TBD  |  CAM  ; 
 TIA <= qfb & qhb ; 
 TIB <= qfb & qhb ; 
 TMA <= qfb & QHB ; 
 TMB <= qfb & QHB ; 
 DBC <= DIC ; 
 DBG <= DIG ; 
 OIM <= NBS ; 
 OCY <=  NBE  |  IAO & TBD  |  CAO  ; 
 ODY <=  NBE  |  IAO & TBD  |  CAO  ; 
 DIC <= ILC ; 
 OLC <= ILC ; 
 AMA <=  ICA & TPD  |  BEA & TUD  ; 
 OEA <=  ICA & TPD  |  BEA & TUD  ; 
 OFA <=  ICA & TPD  |  BEA & TUD  ; 
 DID <= ILD ; 
 OLD <= ILD ; 
 AMG <=  ICG & TPD  |  BEG & TUD  ; 
 OEG <=  ICG & TPD  |  BEG & TUD  ; 
 OFG <=  ICG & TPD  |  BEG & TUD  ; 
 ADK <=  ICO & TMB  |  ADK & TIB  |  ECK & TGD  ; 
 AEK <=  ICO & TMB  |  ADK & TIB  |  ECK & TGD  ; 
 AFK <=  ICO & TMB  |  ADK & TIB  |  ECK & TGD  ; 
 AML <=  ICL & TPD  |  BEL & TUD  ; 
 ODP <=  NAP  |  IAF & TBD  |  CAF  ; 
 ADC <=  ICG & TMB  |  ADC & TIB  |  ECC & TGD  ; 
 AEC <=  ICG & TMB  |  ADC & TIB  |  ECC & TGD  ; 
 AFC <=  ICG & TMB  |  ADC & TIB  |  ECC & TGD  ; 
 ADG <=  ICK & TMB  |  ADG & TIB  |  ECG & TGD  ; 
 AEG <=  ICK & TMB  |  ADG & TIB  |  ECG & TGD  ; 
 AFG <=  ICK & TMB  |  ADG & TIB  |  ECG & TGD  ; 
 ADD <=  ICH & TMB  |  ADD & TIB  |  ECD & TGD  ; 
 AED <=  ICH & TMB  |  ADD & TIB  |  ECD & TGD  ; 
 AFD <=  ICH & TMB  |  ADD & TIB  |  ECD & TGD  ; 
 ADH <=  ICL & TMB  |  ADH & TIB  |  ECH & TGD  ; 
 AEH <=  ICL & TMB  |  ADH & TIB  |  ECH & TGD  ; 
 AFH <=  ICL & TMB  |  ADH & TIB  |  ECH & TGD  ; 
 eal <=  EAL & FAL  |  eal & fal  |  QDG  ; 
 ebl <=  EAL & FAL  |  eal & fal  |  QDG  ; 
 ecl <=  EAL & FAL  |  eal & fal  |  QDG  ; 
 OEL <=  ICL & TPD  |  BEL & TUD  ; 
 OFL <=  ICL & TPD  |  BEL & TUD  ; 
 ADL <=  QRA & TMB  |  ADL & TIB  |  ECL & TGD  ; 
 AEL <=  QRA & TMB  |  ADL & TIB  |  ECL & TGD  ; 
 AFL <=  QRA & TMB  |  ADL & TIB  |  ECL & TGD  ; 
 DBD <= DID ; 
 OIF <= NBL ; 
 DBH <= DIH ; 
 OCR <=  NAR  |  IAH & TBD  |  CAH  ; 
 ODR <=  NAR  |  IAH & TBD  |  CAH  ; 
 QQA <= IQA ; 
 AMP <=  ICP & TPD  |  BEP & TUD  ; 
 OEP <=  ICP & TPD  |  BEP & TUD  ; 
 OFP <=  ICP & TPD  |  BEP & TUD  ; 
 eak <=  EAK & FAK  |  eak & fak  |  QDG  ; 
 ebk <=  EAK & FAK  |  eak & fak  |  QDG  ; 
 eck <=  EAK & FAK  |  eak & fak  |  QDG  ; 
 OCP <=  NAP  |  IAF & TBD  |  CAF  ; 
 TBD <= QQA ; 
 TBH <= QQA ; 
 TPD <= QPA ; 
 TUD <= QPB ; 
 BDM <= BCM ; 
 ebb <=  EAB & FAB  |  eab & fab  |  QDH  ; 
 PCG <=  PBR & pbb & paf  |  pbr & PBB & paf  |  pbr & pbb & PAF  |  PBR & PBB & PAF  ;
 PDC <=  PCH & pcg & pcf  |  pch & PCG & pcf  |  pch & pcg & PCF  |  PCH & PCG & PCF  ;
 PCH <=  PBI & pam & pbl  |  pbi & PAM & pbl  |  pbi & pam & PBL  |  PBI & PAM & PBL  ;
 BDE <= BCE ; 
 BCE <= BBE ; 
 BCM <= BBM ; 
 BEE <= BDE ; 
 BEM <= BDM ; 
 pam <= nam ; 
 pbi <= nbi ; 
 eaa <=  EAA & QIA  |  eaa & qia  |  QDH  ; 
 eba <=  EAA & QIA  |  eaa & qia  |  QDH  ; 
 eca <=  EAA & QIA  |  eaa & qia  |  QDH  ; 
 eae <=  EAE & FAE  |  eae & fae  |  QDH  ; 
 ebe <=  EAE & FAE  |  eae & fae  |  QDH  ; 
 ece <=  EAE & FAE  |  eae & fae  |  QDH  ; 
 eaf <=  EAF & FAF  |  eaf & faf  |  QDH  ; 
 ebf <=  EAF & FAF  |  eaf & faf  |  QDH  ; 
 ecf <=  EAF & FAF  |  eaf & faf  |  QDH  ; 
 paf <= naf ; 
 pbb <= nbb ; 
 pbr <= nbr ; 
 eab <=  EAB & FAB  |  eab & fab  |  QDH  ; 
 ecb <=  EAB & FAB  |  eab & fab  |  QDH  ; 
 BDD <= BCD ; 
 BDJ <= BCJ ; 
 BCD <= BBD ; 
 BCJ <= BBJ ; 
 BED <= BDD ; 
 BEJ <= BDJ ; 
 eai <=  EAI & FAI  |  eai & fai  |  QDH  ; 
 ebi <=  EAI & FAI  |  eai & fai  |  QDH  ; 
 eci <=  EAI & FAI  |  eai & fai  |  QDH  ; 
 BAM <=  NAM  |  IAC & TBE  |  CAC  ; 
 OAM <=  NAM  |  IAC & TBE  |  CAC  ; 
 OBM <=  NAM  |  IAC & TBE  |  CAC  ; 
 tnc <=  qhc  |  QFB  |  ira  ; 
 tnd <=  qhc  |  QFB  |  IRA  ; 
 dca <= dia ; 
 dce <= die ; 
 OIC <= NBI ; 
 BAS <=  NAS  |  IAI & TBE  |  CAI  ; 
 OAS <=  NAS  |  IAI & TBE  |  CAI  ; 
 OBS <=  NAS  |  IAI & TBE  |  CAI  ; 
 bbe <= ice ; 
 bbm <= icm ; 
 DIE <= ILE ; 
 OLE <= ILE ; 
 ogm <=  icm & tua  |  bem & tpa  |  tpa & tua  ; 
 ohm <=  icm & tua  |  bem & tpa  |  tpa & tua  ; 
 fbb <=  eaf  |  eag  |  eah  |  eai  ; 
 BAL <=  NAL  |  IAB & TBE  |  CAB  ; 
 oge <=  ice & tua  |  bee & tpa  |  tpa & tua  ; 
 ohe <=  ice & tua  |  bee & tpa  |  tpa & tua  ; 
 agi <=  icm & TNA  |  agi & TJA  |  eci & TGE  ; 
 ahi <=  icm & TNA  |  agi & TJA  |  eci & TGE  ; 
 aii <=  icm & TNA  |  agi & TJA  |  eci & TGE  ; 
 aha <=  ice & TNC  |  iga & TND  |  aha & TJA  |  eca & TGE  ; 
 aia <=  ice & TNC  |  iga & TND  |  aha & TJA  |  eca & TGE  ; 
 ahe <=  ici & TNA  |  age & TJA  |  ece & TGE  ; 
 aie <=  ici & TNA  |  age & TJA  |  ece & TGE  ; 
 age <=  ici & TNA  |  age & TJA  |  ece & TGE  ; 
 ohd <=  icd & tua  |  bed & tpa  |  tpa & tua  ; 
 agb <=  icf & TNA  |  agb & TJA  |  ecb & TGE  ; 
 ahb <=  icf & TNA  |  agb & TJA  |  ecb & TGE  ; 
 aib <=  icf & TNA  |  agb & TJA  |  ecb & TGE  ; 
 agf <=  icj & TNA  |  agf & TJA  |  ecf & TGE  ; 
 ahf <=  icj & TNA  |  agf & TJA  |  ecf & TGE  ; 
 aif <=  icj & TNA  |  agf & TJA  |  ecf & TGE  ; 
 eaj <=  EAJ & FAJ  |  eaj & faj  |  QDH  ; 
 ebj <=  EAJ & FAJ  |  eaj & faj  |  QDH  ; 
 ecj <=  EAJ & FAJ  |  eaj & faj  |  QDH  ; 
 ogj <=  icj & tua  |  bej & tpa  |  tpa & tua  ; 
 ohj <=  icj & tua  |  bej & tpa  |  tpa & tua  ; 
 agj <=  icn & TNA  |  agj & TJA  |  ecj & TGE  ; 
 ahj <=  icn & TNA  |  agj & TJA  |  ecj & TGE  ; 
 aij <=  icn & TNA  |  agj & TJA  |  ecj & TGE  ; 
 dcb <= dib ; 
 dcf <= dif ; 
 OIL <= NBR ; 
 BAV <=  NBB  |  IAL & TBE  |  CAL  ; 
 OAV <=  NBB  |  IAL & TBE  |  CAL  ; 
 OBV <=  NBB  |  IAL & TBE  |  CAL  ; 
 bbd <= icd ; 
 bbj <= icj ; 
 DIF <= ILF ; 
 OLF <= ILF ; 
 ogd <=  icd & tua  |  bed & tpa  |  tpa & tua  ; 
 OAF <= NAF ; 
 OBF <= NAF ; 
 OCF <= NAF ; 
 ODF <= NAF ; 
 OAL <=  NAL  |  IAB & TBE  |  CAB  ; 
 OBL <=  NAL  |  IAB & TBE  |  CAB  ; 
 OKA <=  BFA & TEA  ; 
 PCI <=  PBH & pal & pap  |  pbh & PAL & pap  |  pbh & pal & PAP  |  PBH & PAL & PAP  ;
 PDB <=  PCK & pcj & pci  |  pck & PCJ & pci  |  pck & pcj & PCI  |  PCK & PCJ & PCI  ;
 PCJ <=  PBO & pas & pac  |  pbo & PAS & pac  |  pbo & pas & PAC  |  PBO & PAS & PAC  ;
 BDK <= BCK ; 
 BDO <= BCO ; 
 BCK <= BBK ; 
 BCO <= BBO ; 
 BEK <= BDK ; 
 BEO <= BDO ; 
 QHC <=  qga & QGB  ; 
 QHD <=  QGA & QGB  ; 
 pac <= nac ; 
 pas <= nas ; 
 pbo <= nbo ; 
 QGA <=  qga & qfa  ; 
 QGC <=  qga & qfa  ; 
 QGE <=  qga & qfa  ; 
 QGB <=  QGB & qga & qfa  |  qgb & QGA  ; 
 QGD <=  QGB & qga & qfa  |  qgb & QGA  ; 
 QGF <=  QGB & qga & qfa  |  qgb & QGA  ; 
 pal <= nal ; 
 pbh <= nbh ; 
 BFA <= BDA & bdd |  bda & BDD ; 
 BFB <= BDB & bdd |  bdb & BDD ; 
 BFC <= BDC & bdd |  bdc & BDD ; 
 QMB <=  BBN & bbo  ; 
 BDB <= BCB ; 
 BDH <= BCH ; 
 QMA <= BBO ; 
 BCB <= BBB ; 
 BCH <= BBH ; 
 BEB <= BDB ; 
 BEH <= BDH ; 
 QHA <=  qga & qgb  ; 
 QHB <=  QGA & qgb  ; 
 OAC <= NAC ; 
 OBC <= NAC ; 
 OCC <= NAC ; 
 ODC <= NAC ; 
 OCM <=  NAM  |  IAC & TBF  |  CAC  ; 
 ODM <=  NAM  |  IAC & TBF  |  CAC  ; 
 TJA <= qfb & qhc ; 
 TJB <= qfb & qhc ; 
 TNA <= qfb & QHC ; 
 TNB <= qfb & QHC ; 
 dcc <= dic ; 
 dcg <= dig ; 
 OII <= NBO ; 
 OCS <=  NAS  |  IAI & TBF  |  CAI  ; 
 ODS <=  NAS  |  IAI & TBF  |  CAI  ; 
 bbk <= ick ; 
 bbo <= ico ; 
 DIG <= ILG ; 
 OLG <= ILG ; 
 ogo <=  ico & tub  |  beo & tpb  |  tpb & tub  ; 
 oho <=  ico & tub  |  beo & tpb  |  tpb & tub  ; 
 bbb <= icb ; 
 bbh <= ich ; 
 DIH <= ILH ; 
 OLH <= ILH ; 
 ogk <=  ick & tub  |  bek & tpb  |  tpb & tub  ; 
 ohk <=  ick & tub  |  bek & tpb  |  tpb & tub  ; 
 agk <=  ico & TNB  |  agk & TJB  |  eck & TGF  ; 
 ahk <=  ico & TNB  |  agk & TJB  |  eck & TGF  ; 
 aik <=  ico & TNB  |  agk & TJB  |  eck & TGF  ; 
 agc <=  icg & TNB  |  agc & TJB  |  ecc & TGF  ; 
 ahc <=  icg & TNB  |  agc & TJB  |  ecc & TGF  ; 
 aic <=  icg & TNB  |  agc & TJB  |  ecc & TGF  ; 
 agg <=  ick & TNB  |  agg & TJB  |  ecg & TGF  ; 
 ahg <=  ick & TNB  |  agg & TJB  |  ecg & TGF  ; 
 aig <=  ick & TNB  |  agg & TJB  |  ecg & TGF  ; 
 agd <=  ich & TNB  |  agd & TJB  |  ecd & TGF  ; 
 ahd <=  ich & TNB  |  agd & TJB  |  ecd & TGF  ; 
 aid <=  ich & TNB  |  agd & TJB  |  ecd & TGF  ; 
 agh <=  icl & TNB  |  agh & TJB  |  ech & TGF  ; 
 ahh <=  icl & TNB  |  agh & TJB  |  ech & TGF  ; 
 aih <=  icl & TNB  |  agh & TJB  |  ech & TGF  ; 
 ogh <=  ich & tub  |  beh & tpb  |  tpb & tub  ; 
 ohh <=  ich & tub  |  beh & tpb  |  tpb & tub  ; 
 agl <=  qra & TNB  |  agl & TJB  |  ecl & TGF  ; 
 ahl <=  qra & TNB  |  agl & TJB  |  ecl & TGF  ; 
 ail <=  qra & TNB  |  agl & TJB  |  ecl & TGF  ; 
 dcd <= did ; 
 dch <= dih ; 
 OIB <= NBH ; 
 TEA <= QMA ; 
 OCV <=  NBB  |  IAL & TBF  |  CAL  ; 
 ODV <=  NBB  |  IAL & TBF  |  CAL  ; 
 ogb <=  icb & tub  |  beb & tpb  |  tpb & tub  ; 
 ohb <=  icb & tub  |  beb & tpb  |  tpb & tub  ; 
 QNA <= IRB & QMA ; 
 QNB <= IRB & QMB ; 
 QNC <= IRB & QMC ; 
 QND <= IRB & QMD ; 
 TEC <=  QNC  |  QNE  ; 
 TED <=  QND  |  QNF  ; 
 OCL <=  NAL  |  IAB & TBF  |  CAB  ; 
 ODL <=  NAL  |  IAB & TBF  |  CAB  ; 
 OKB <=  BFB & TEA  |  BFA & TEB  ; 
 OKC <=  BFC & TEA  |  BFB & TEB  |  BFA & TEC  ; 
 PEB <=  PDA & pdb & pdc  |  pda & PDB & pdc  |  pda & pdb & PDC  |  PDA & PDB & PDC  ;
 PCK <=  PBQ & pba & pae  |  pbq & PBA & pae  |  pbq & pba & PAE  |  PBQ & PBA & PAE  ;
 tqq <= qhg ; 
 trq <= qhk ; 
 tsq <= qho ; 
 ttq <= qhs ; 
 TQN <= QHG ; 
 TRN <= QHK ; 
 TSN <= QHO ; 
 TTN <= QHS ; 
 BDC <= BCC ; 
 BDI <= BCI ; 
 BCC <= BBC ; 
 BCI <= BBI ; 
 BEC <= BDC ; 
 BEI <= BDI ; 
 pae <= nae ; 
 pba <= nba ; 
 pbq <= nbq ; 
 qhk <=  qge  |  QGF  |  qjb  ; 
 qhl <=  qge  |  QGF  |  qjb  ; 
 qhg <=  QGE  |  QGF  |  qjb  ; 
 qhh <=  QGE  |  QGF  |  qjb  ; 
 tqi <= qhg ; 
 trii <= qhk ; 
 tsi <= qho ; 
 tti <= qhs ; 
 AMF <=  ICF & TPC  |  BEF & TUC  ; 
 TQF <= QHG ; 
 TRF <= QHK ; 
 TSF <= QHO ; 
 TTF <= QHS ; 
 pan <= nan ; 
 pbj <= nbj ; 
 OLI <= ILI ; 
 qmc <=  bbm  |  BBM  |  BBO  ; 
 qmd <=  BBM  |  BBN  |  BBO  ; 
 BDF <= BCF ; 
 BDN <= BCN ; 
 BCF <= BBF ; 
 BCN <= BBN ; 
 BEF <= BDF ; 
 BEN <= BDN ; 
 OAE <= NAE ; 
 OBE <= NAE ; 
 OCE <= NAE ; 
 ODE <= NAE ; 
 BAK <=  NAK  |  IAA & TBG  |  CAA  ; 
 OAK <=  NAK  |  IAA & TBG  |  CAA  ; 
 OBK <=  NAK  |  IAA & TBG  |  CAA  ; 
 toc <=  qhd  |  QFB  |  ira  ; 
 tod <=  qhd  |  QFB  |  IRA  ; 
 dda <= dia ; 
 dde <= die ; 
 OIK <= NBQ ; 
 BAU <=  NBA  |  IAK & TBG  |  CAK  ; 
 OAU <=  NBA  |  IAK & TBG  |  CAK  ; 
 OBU <=  NBA  |  IAK & TBG  |  CAK  ; 
 bbc <= icc ; 
 bbi <= ici ; 
 oja <= iga ; 
 QRA <= IRA ; 
 ogc <=  icc & tuc  |  bec & tpc  |  tpc & tuc  ; 
 ohc <=  icc & tuc  |  bec & tpc  |  tpc & tuc  ; 
 OBN <=  NAN  |  IAD & TBG  |  CAD  ; 
 ogi <=  ici & tuc  |  bei & tpc  |  tpc & tuc  ; 
 ohi <=  ici & tuc  |  bei & tpc  |  tpc & tuc  ; 
 aji <=  icm & TOA  |  aji & TKA  |  eci & TGG  ; 
 aki <=  icm & TOA  |  aji & TKA  |  eci & TGG  ; 
 ali <=  icm & TOA  |  aji & TKA  |  eci & TGG  ; 
 aka <=  ice & TOC  |  iga & TOD  |  aka & TKA  |  eca & TGG  ; 
 ala <=  ice & TOC  |  iga & TOD  |  aka & TKA  |  eca & TGG  ; 
 aje <=  ici & TOA  |  aje & TKA  |  ece & TGG  ; 
 ake <=  ici & TOA  |  aje & TKA  |  ece & TGG  ; 
 ale <=  ici & TOA  |  aje & TKA  |  ece & TGG  ; 
 ajb <=  icf & TOA  |  ajb & TKA  |  ecb & TGG  ; 
 akb <=  icf & TOA  |  ajb & TKA  |  ecb & TGG  ; 
 alb <=  icf & TOA  |  ajb & TKA  |  ecb & TGG  ; 
 ajf <=  icj & TOA  |  ajf & TKA  |  ecf & TGG  ; 
 akf <=  icj & TOA  |  ajf & TKA  |  ecf & TGG  ; 
 alf <=  icj & TOA  |  ajf & TKA  |  ecf & TGG  ; 
 tqa <= qhg ; 
 tra <= qhk ; 
 tsa <= qho ; 
 tta <= qhs ; 
 bbf <= icf ; 
 bbn <= icn ; 
 TEB <= QNB ; 
 TEE <= QNG ; 
 ogf <=  icf & tuc  |  bef & tpc  |  tpc & tuc  ; 
 ohf <=  icf & tuc  |  bef & tpc  |  tpc & tuc  ; 
 ajj <=  icn & TOA  |  ajj & TKA  |  ecj & TGG  ; 
 akj <=  icn & TOA  |  ajj & TKA  |  ecj & TGG  ; 
 alj <=  icn & TOA  |  ajj & TKA  |  ecj & TGG  ; 
 ddb <= dib ; 
 ddf <= dif ; 
 OID <= NBJ ; 
 BAT <=  NAT  |  IAJ & TBG  |  CAJ  ; 
 OAT <=  NAT  |  IAJ & TBG  |  CAJ  ; 
 OBT <=  NAT  |  IAJ & TBG  |  CAJ  ; 
 ogn <=  icn & tuc  |  ben & tpc  |  tpc & tuc  ; 
 ohn <=  icn & tuc  |  ben & tpc  |  tpc & tuc  ; 
 QNE <=  QME & ISA  ; 
 QNG <=  QMF & ISA  ; 
 BAN <=  NAN  |  IAD & TBG  |  CAD  ; 
 OAN <=  NAN  |  IAD & TBG  |  CAD  ; 
 OKD <=  TEB & BFC  |  TEC & BFB  |  TED & BFA  ; 
 OKE <=  TEC & BFC  |  TED & BFB  |  TEE & BFA  ; 
 TQP <= QHH ; 
 TSP <= QHP ; 
 TTP <= QHT ; 
 PCL <=  PBP & pat & pad  |  pbp & PAT & pad  |  pbp & pat & PAD  |  PBP & PAT & PAD  ;
 PDA <=  PCM & pcn & pcl  |  pcm & PCN & pcl  |  pcm & pcn & PCL  |  PCM & PCN & PCL  ;
 PCM <=  PBG & pak & pbj  |  pbg & PAK & pbj  |  pbg & pak & PBJ  |  PBG & PAK & PBJ  ;
 PCN <= PAN ; 
 tqs <= qhh ; 
 trs <= qhl ; 
 tss <= qhp ; 
 tts <= qht ; 
 TRP <= QHL ; 
 BDA <= BCA ; 
 BDG <= BCG ; 
 BCA <= BBA ; 
 BCG <= BBG ; 
 BEA <= BDA ; 
 BEG <= BDG ; 
 pak <= nak ; 
 pbg <= nbg ; 
 tqk <= qhh ; 
 qhs <=  qge  |  qgf  |  qjb  ; 
 qht <=  qge  |  qgf  |  qjb  ; 
 qho <=  QGE  |  qgf  |  qjb  ; 
 qhp <=  QGE  |  qgf  |  qjb  ; 
 trk <= qhl ; 
 tsk <= qhp ; 
 ttk <= qht ; 
 tqg <= qhh ; 
 trg <= qhl ; 
 tsg <= qhp ; 
 ttg <= qht ; 
 WBE <= QEB & QBH ; 
 WBF <= QEB & QBH ; 
 WBG <= QEB & QBH ; 
 WBH <= QEB & QBH ; 
 WCA <= QEB & QBF ; 
 WCB <= QEB & QBF ; 
 WCC <= QEB & QBF ; 
 WCD <= QEB & QBF ; 
 WCE <= QEB & QBF ; 
 WCF <= QEB & QBF ; 
 WCG <= QEB & QBF ; 
 WCH <= QEB & QBF ; 
 WBA <= QEB & QBH ; 
 WBB <= QEB & QBH ; 
 WBC <= QEB & QBH ; 
 WBD <= QEB & QBH ; 
 pad <= nad ; 
 pat <= nat ; 
 pbp <= nbp ; 
 QME <=  BBN & BBO  ; 
 BDL <= BCL ; 
 BDP <= BCP ; 
 QMF <=  bbn & bbo  ; 
 BCL <= BBL ; 
 BCP <= BBP ; 
 BEL <= BDL ; 
 BEP <= BDP ; 
 OCK <=  NAK  |  IAA & TBH  |  CAA  ; 
 ODK <=  NAK  |  IAA & TBH  |  CAA  ; 
 TKA <= qfb & qhd ; 
 TKB <= qfb & qhd ; 
 TOA <= qfb & QHD ; 
 TOB <= qfb & QHD ; 
 ddc <= dic ; 
 ddg <= dig ; 
 OIA <= NBG ; 
 OCU <=  NBA  |  IAK & TBH  |  CAK  ; 
 ODU <=  NBA  |  IAK & TBH  |  CAK  ; 
 bba <= ica ; 
 bbg <= icg ; 
 oga <=  ica & tud  |  bea & tpd  |  tpd & tud  ; 
 oha <=  ica & tud  |  bea & tpd  |  tpd & tud  ; 
 bbl <= icl ; 
 bbp <= icp ; 
 tge <= qfa ; 
 ogg <=  icg & tud  |  beg & tpd  |  tpd & tud  ; 
 ohg <=  icg & tud  |  beg & tpd  |  tpd & tud  ; 
 ajk <=  ico & TOB  |  ajk & TKB  |  eck & TGH  ; 
 akk <=  ico & TOB  |  ajk & TKB  |  eck & TGH  ; 
 alk <=  ico & TOB  |  ajk & TKB  |  eck & TGH  ; 
 ogl <=  icl & tud  |  bel & tpd  |  tpd & tud  ; 
 ajc <=  icg & TOB  |  ajc & TKB  |  ecc & TGH  ; 
 akc <=  icg & TOB  |  ajc & TKB  |  ecc & TGH  ; 
 alc <=  icg & TOB  |  ajc & TKB  |  ecc & TGH  ; 
 ajg <=  ick & TOB  |  ajg & TKB  |  ecg & TGH  ; 
 akg <=  ick & TOB  |  ajg & TKB  |  ecg & TGH  ; 
 alg <=  ick & TOB  |  ajg & TKB  |  ecg & TGH  ; 
 tgf <= qfa ; 
 tgg <= qfa ; 
 tgh <= qfa ; 
 ajd <=  ich & TOB  |  ajd & TKB  |  ecd & TGH  ; 
 akd <=  ich & TOB  |  ajd & TKB  |  ecd & TGH  ; 
 ald <=  ich & TOB  |  ajd & TKB  |  ecd & TGH  ; 
 ajh <=  icl & TOB  |  ajh & TKB  |  ech & TGH  ; 
 akh <=  icl & TOB  |  ajh & TKB  |  ech & TGH  ; 
 alh <=  icl & TOB  |  ajh & TKB  |  ech & TGH  ; 
 TQD <= QHH ; 
 TRD <= QHL ; 
 TSD <= QHP ; 
 TTD <= QHT ; 
 ohl <=  icl & tud  |  bel & tpd  |  tpd & tud  ; 
 ajl <=  qra & TOB  |  ajl & TKB  |  ecl & TGH  ; 
 akl <=  qra & TOB  |  ajl & TKB  |  ecl & TGH  ; 
 all <=  qra & TOB  |  ajl & TKB  |  ecl & TGH  ; 
 ddd <= did ; 
 ddh <= dih ; 
 OIJ <= NBP ; 
 OCT <=  NAT  |  IAJ & TBH  |  CAJ  ; 
 ODT <=  NAT  |  IAJ & TBH  |  CAJ  ; 
 ogp <=  icp & tud  |  bep & tpd  |  tpd & tud  ; 
 ohp <=  icp & tud  |  bep & tpd  |  tpd & tud  ; 
 QNF <=  qme & qmf & ISA  ; 
 OAD <= NAD ; 
 OBD <= NAD ; 
 OCD <= NAD ; 
 ODD <= NAD ; 
 OCN <=  NAN  |  IAD & TBH  |  CAD  ; 
 ODN <=  NAN  |  IAD & TBH  |  CAD  ; 
 OKF <=  TED & BFC  |  BFB & TEE  ; 
 OKG <=  TEE & BFC  ; 
end 
ram_4096x1 sinst_000(MAA,DAA,{AAA,AAB,AAC,AAD,AAE,AAF,AAG,AAH,AAI,AAJ,AAK,AAL}, ZZI, WAA, IZZ); 
ram_4096x1 sinst_001(MCA,DBA,{AEA,AEB,AEC,AED,AEE,AEF,AEG,AEH,AEI,AEJ,AEK,AEL}, ZZI, WAA, IZZ); 
ram_4096x1 sinst_002(MEA,DCA,{AHA,AHB,AHC,AHD,AHE,AHF,AHG,AHH,AHI,AHJ,AHK,AHL}, ZZI, WAA, IZZ); 
ram_4096x1 sinst_003(MGA,DDA,{AKA,AKB,AKC,AKD,AKE,AKF,AKG,AKH,AKI,AKJ,AKK,AKL}, ZZI, WAA, IZZ); 
ram_4096x1 sinst_004(MAB,DAB,{aaa,aab,aac,aad,aae,aaf,aag,aah,aai,aaj,aak,aal}, ZZI, WAB, IZZ); 
ram_4096x1 sinst_005(MCB,DBB,{aea,aeb,aec,aed,aee,aef,aeg,aeh,aei,aej,aek,ael}, ZZI, WAB, IZZ); 
ram_4096x1 sinst_006(MEB,DCB,{aha,ahb,ahc,ahd,ahe,ahf,ahg,ahh,ahi,ahj,ahk,ahl}, ZZI, WAB, IZZ); 
ram_4096x1 sinst_007(MGB,DDB,{aka,akb,akc,akd,ake,akf,akg,akh,aki,akj,akk,akl}, ZZI, WAB, IZZ); 
ram_4096x1 sinst_008(MAC,DAC,{ABA,ABB,ABC,ABD,ABE,ABF,ABG,ABH,ABI,ABJ,ABK,ABL}, ZZI, WAC, IZZ); 
ram_4096x1 sinst_009(MCC,DBC,{AFA,AFB,AFC,AFD,AFE,AFF,AFG,AFH,AFI,AFJ,AFK,AFL}, ZZI, WAC, IZZ); 
ram_4096x1 sinst_010(MEC,DCC,{AIA,AIB,AIC,AID,AIE,AIF,AIG,AIH,AII,AIJ,AIK,AIL}, ZZI, WAC, IZZ); 
ram_4096x1 sinst_011(MGC,DDC,{ALA,ALB,ALC,ALD,ALE,ALF,ALG,ALH,ALI,ALJ,ALK,ALL}, ZZI, WAC, IZZ); 
ram_4096x1 sinst_012(MAD,DAD,{aba,abb,abc,abd,abe,abf,abg,abh,abi,abj,abk,abl}, ZZI, WAD, IZZ); 
ram_4096x1 sinst_013(MCD,DBD,{afa,afb,afc,afd,afe,aff,afg,afh,afi,afj,afk,afl}, ZZI, WAD, IZZ); 
ram_4096x1 sinst_014(MED,DCD,{aia,aib,aic,aid,aie,aif,aig,aih,aii,aij,aik,ail}, ZZI, WAD, IZZ); 
ram_4096x1 sinst_015(MGD,DDD,{ala,alb,alc,ald,ale,alf,alg,alh,ali,alj,alk,all}, ZZI, WAD, IZZ); 
ram_4096x1 sinst_016(MAE,DAE,{AAA,AAB,AAC,AAD,AAE,AAF,AAG,AAH,AAI,AAJ,AAK,AAL}, ZZI, WAE, IZZ); 
ram_4096x1 sinst_017(MCE,DBE,{AEA,AEB,AEC,AED,AEE,AEF,AEG,AEH,AEI,AEJ,AEK,AEL}, ZZI, WAE, IZZ); 
ram_4096x1 sinst_018(MEE,DCE,{AHA,AHB,AHC,AHD,AHE,AHF,AHG,AHH,AHI,AHJ,AHK,AHL}, ZZI, WAE, IZZ); 
ram_4096x1 sinst_019(MGE,DDE,{AKA,AKB,AKC,AKD,AKE,AKF,AKG,AKH,AKI,AKJ,AKK,AKL}, ZZI, WAE, IZZ); 
ram_4096x1 sinst_020(MAF,DAF,{aaa,aab,aac,aad,aae,aaf,aag,aah,aai,aaj,aak,aal}, ZZI, WAF, IZZ); 
ram_4096x1 sinst_021(MCF,DBF,{aea,aeb,aec,aed,aee,aef,aeg,aeh,aei,aej,aek,ael}, ZZI, WAF, IZZ); 
ram_4096x1 sinst_022(MEF,DCF,{aha,ahb,ahc,ahd,ahe,ahf,ahg,ahh,ahi,ahj,ahk,ahl}, ZZI, WAF, IZZ); 
ram_4096x1 sinst_023(MGF,DDF,{aka,akb,akc,akd,ake,akf,akg,akh,aki,akj,akk,akl}, ZZI, WAF, IZZ); 
ram_4096x1 sinst_024(MAG,DAG,{ABA,ABB,ABC,ABD,ABE,ABF,ABG,ABH,ABI,ABJ,ABK,ABL}, ZZI, WAG, IZZ); 
ram_4096x1 sinst_025(MCG,DBG,{AFA,AFB,AFC,AFD,AFE,AFF,AFG,AFH,AFI,AFJ,AFK,AFL}, ZZI, WAG, IZZ); 
ram_4096x1 sinst_026(MEG,DCG,{AIA,AIB,AIC,AID,AIE,AIF,AIG,AIH,AII,AIJ,AIK,AIL}, ZZI, WAG, IZZ); 
ram_4096x1 sinst_027(MGG,DDG,{ALA,ALB,ALC,ALD,ALE,ALF,ALG,ALH,ALI,ALJ,ALK,ALL}, ZZI, WAG, IZZ); 
ram_4096x1 sinst_028(MAH,DAH,{aba,abb,abc,abd,abe,abf,abg,abh,abi,abj,abk,abl}, ZZI, WAH, IZZ); 
ram_4096x1 sinst_029(MCH,DBH,{afa,afb,afc,afd,afe,aff,afg,afh,afi,afj,afk,afl}, ZZI, WAH, IZZ); 
ram_4096x1 sinst_030(MEH,DCH,{aia,aib,aic,aid,aie,aif,aig,aih,aii,aij,aik,ail}, ZZI, WAH, IZZ); 
ram_4096x1 sinst_031(MGH,DDH,{ala,alb,alc,ald,ale,alf,alg,alh,ali,alj,alk,all}, ZZI, WAH, IZZ); 
ram_4096x1 sinst_032(MAI,DAA,{AAA,AAB,AAC,AAD,AAE,AAF,AAG,AAH,AAI,AAJ,AAK,AAL}, ZZI, WBA, IZZ); 
ram_4096x1 sinst_033(MCI,DBA,{AEA,AEB,AEC,AED,AEE,AEF,AEG,AEH,AEI,AEJ,AEK,AEL}, ZZI, WBA, IZZ); 
ram_4096x1 sinst_034(MEI,DCA,{AHA,AHB,AHC,AHD,AHE,AHF,AHG,AHH,AHI,AHJ,AHK,AHL}, ZZI, WBA, IZZ); 
ram_4096x1 sinst_035(MGI,DDA,{AKA,AKB,AKC,AKD,AKE,AKF,AKG,AKH,AKI,AKJ,AKK,AKL}, ZZI, WBA, IZZ); 
ram_4096x1 sinst_036(MAJ,DAB,{aaa,aab,aac,aad,aae,aaf,aag,aah,aai,aaj,aak,aal}, ZZI, WBB, IZZ); 
ram_4096x1 sinst_037(MCJ,DBB,{aea,aeb,aec,aed,aee,aef,aeg,aeh,aei,aej,aek,ael}, ZZI, WBB, IZZ); 
ram_4096x1 sinst_038(MEJ,DCB,{aha,ahb,ahc,ahd,ahe,ahf,ahg,ahh,ahi,ahj,ahk,ahl}, ZZI, WBB, IZZ); 
ram_4096x1 sinst_039(MGJ,DDB,{aka,akb,akc,akd,ake,akf,akg,akh,aki,akj,akk,akl}, ZZI, WBB, IZZ); 
ram_4096x1 sinst_040(MAK,DAC,{ABA,ABB,ABC,ABD,ABE,ABF,ABG,ABH,ABI,ABJ,ABK,ABL}, ZZI, WBC, IZZ); 
ram_4096x1 sinst_041(MCK,DBC,{AFA,AFB,AFC,AFD,AFE,AFF,AFG,AFH,AFI,AFJ,AFK,AFL}, ZZI, WBC, IZZ); 
ram_4096x1 sinst_042(MEK,DCC,{AIA,AIB,AIC,AID,AIE,AIF,AIG,AIH,AII,AIJ,AIK,AIL}, ZZI, WBC, IZZ); 
ram_4096x1 sinst_043(MGK,DDC,{ALA,ALB,ALC,ALD,ALE,ALF,ALG,ALH,ALI,ALJ,ALK,ALL}, ZZI, WBC, IZZ); 
ram_4096x1 sinst_044(MAL,DAD,{aba,abb,abc,abd,abe,abf,abg,abh,abi,abj,abk,abl}, ZZI, WBD, IZZ); 
ram_4096x1 sinst_045(MCL,DBD,{afa,afb,afc,afd,afe,aff,afg,afh,afi,afj,afk,afl}, ZZI, WBD, IZZ); 
ram_4096x1 sinst_046(MEL,DCD,{aia,aib,aic,aid,aie,aif,aig,aih,aii,aij,aik,ail}, ZZI, WBD, IZZ); 
ram_4096x1 sinst_047(MGL,DDD,{ala,alb,alc,ald,ale,alf,alg,alh,ali,alj,alk,all}, ZZI, WBD, IZZ); 
ram_4096x1 sinst_048(MAM,DAE,{AAA,AAB,AAC,AAD,AAE,AAF,AAG,AAH,AAI,AAJ,AAK,AAL}, ZZI, WBE, IZZ); 
ram_4096x1 sinst_049(MCM,DBE,{AEA,AEB,AEC,AED,AEE,AEF,AEG,AEH,AEI,AEJ,AEK,AEL}, ZZI, WBE, IZZ); 
ram_4096x1 sinst_050(MEM,DCE,{AHA,AHB,AHC,AHD,AHE,AHF,AHG,AHH,AHI,AHJ,AHK,AHL}, ZZI, WBE, IZZ); 
ram_4096x1 sinst_051(MGM,DDE,{AKA,AKB,AKC,AKD,AKE,AKF,AKG,AKH,AKI,AKJ,AKK,AKL}, ZZI, WBE, IZZ); 
ram_4096x1 sinst_052(MAN,DAF,{aaa,aab,aac,aad,aae,aaf,aag,aah,aai,aaj,aak,aal}, ZZI, WBF, IZZ); 
ram_4096x1 sinst_053(MCN,DBF,{aea,aeb,aec,aed,aee,aef,aeg,aeh,aei,aej,aek,ael}, ZZI, WBF, IZZ); 
ram_4096x1 sinst_054(MEN,DCF,{aha,ahb,ahc,ahd,ahe,ahf,ahg,ahh,ahi,ahj,ahk,ahl}, ZZI, WBF, IZZ); 
ram_4096x1 sinst_055(MGN,DDF,{aka,akb,akc,akd,ake,akf,akg,akh,aki,akj,akk,akl}, ZZI, WBF, IZZ); 
ram_4096x1 sinst_056(MAO,DAG,{ABA,ABB,ABC,ABD,ABE,ABF,ABG,ABH,ABI,ABJ,ABK,ABL}, ZZI, WBG, IZZ); 
ram_4096x1 sinst_057(MCO,DBG,{AFA,AFB,AFC,AFD,AFE,AFF,AFG,AFH,AFI,AFJ,AFK,AFL}, ZZI, WBG, IZZ); 
ram_4096x1 sinst_058(MEO,DCG,{AIA,AIB,AIC,AID,AIE,AIF,AIG,AIH,AII,AIJ,AIK,AIL}, ZZI, WBG, IZZ); 
ram_4096x1 sinst_059(MGO,DDG,{ALA,ALB,ALC,ALD,ALE,ALF,ALG,ALH,ALI,ALJ,ALK,ALL}, ZZI, WBG, IZZ); 
ram_4096x1 sinst_060(MAP,DAH,{aba,abb,abc,abd,abe,abf,abg,abh,abi,abj,abk,abl}, ZZI, WBH, IZZ); 
ram_4096x1 sinst_061(MCP,DBH,{afa,afb,afc,afd,afe,aff,afg,afh,afi,afj,afk,afl}, ZZI, WBH, IZZ); 
ram_4096x1 sinst_062(MEP,DCH,{aia,aib,aic,aid,aie,aif,aig,aih,aii,aij,aik,ail}, ZZI, WBH, IZZ); 
ram_4096x1 sinst_063(MGP,DDH,{ala,alb,alc,ald,ale,alf,alg,alh,ali,alj,alk,all}, ZZI, WBH, IZZ); 
ram_4096x1 sinst_064(MAQ,DAA,{AAA,AAB,AAC,AAD,AAE,AAF,AAG,AAH,AAI,AAJ,AAK,AAL}, ZZI, WCA, IZZ); 
ram_4096x1 sinst_065(MCQ,DBA,{AEA,AEB,AEC,AED,AEE,AEF,AEG,AEH,AEI,AEJ,AEK,AEL}, ZZI, WCA, IZZ); 
ram_4096x1 sinst_066(MEQ,DCA,{AHA,AHB,AHC,AHD,AHE,AHF,AHG,AHH,AHI,AHJ,AHK,AHL}, ZZI, WCA, IZZ); 
ram_4096x1 sinst_067(MGQ,DDA,{AKA,AKB,AKC,AKD,AKE,AKF,AKG,AKH,AKI,AKJ,AKK,AKL}, ZZI, WCA, IZZ); 
ram_4096x1 sinst_068(MAR,DAB,{aaa,aab,aac,aad,aae,aaf,aag,aah,aai,aaj,aak,aal}, ZZI, WCB, IZZ); 
ram_4096x1 sinst_069(MCR,DBB,{aea,aeb,aec,aed,aee,aef,aeg,aeh,aei,aej,aek,ael}, ZZI, WCB, IZZ); 
ram_4096x1 sinst_070(MER,DCB,{aha,ahb,ahc,ahd,ahe,ahf,ahg,ahh,ahi,ahj,ahk,ahl}, ZZI, WCB, IZZ); 
ram_4096x1 sinst_071(MGR,DDB,{aka,akb,akc,akd,ake,akf,akg,akh,aki,akj,akk,akl}, ZZI, WCB, IZZ); 
ram_4096x1 sinst_072(MAS,DAC,{ABA,ABB,ABC,ABD,ABE,ABF,ABG,ABH,ABI,ABJ,ABK,ABL}, ZZI, WCC, IZZ); 
ram_4096x1 sinst_073(MCS,DBC,{AFA,AFB,AFC,AFD,AFE,AFF,AFG,AFH,AFI,AFJ,AFK,AFL}, ZZI, WCC, IZZ); 
ram_4096x1 sinst_074(MES,DCC,{AIA,AIB,AIC,AID,AIE,AIF,AIG,AIH,AII,AIJ,AIK,AIL}, ZZI, WCC, IZZ); 
ram_4096x1 sinst_075(MGS,DDC,{ALA,ALB,ALC,ALD,ALE,ALF,ALG,ALH,ALI,ALJ,ALK,ALL}, ZZI, WCC, IZZ); 
ram_4096x1 sinst_076(MAT,DAD,{aba,abb,abc,abd,abe,abf,abg,abh,abi,abj,abk,abl}, ZZI, WCD, IZZ); 
ram_4096x1 sinst_077(MCT,DBD,{afa,afb,afc,afd,afe,aff,afg,afh,afi,afj,afk,afl}, ZZI, WCD, IZZ); 
ram_4096x1 sinst_078(MET,DCD,{aia,aib,aic,aid,aie,aif,aig,aih,aii,aij,aik,ail}, ZZI, WCD, IZZ); 
ram_4096x1 sinst_079(MGT,DDD,{ala,alb,alc,ald,ale,alf,alg,alh,ali,alj,alk,all}, ZZI, WCD, IZZ); 
ram_4096x1 sinst_080(MBA,DAE,{AAA,AAB,AAC,AAD,AAE,AAF,AAG,AAH,AAI,AAJ,AAK,AAL}, ZZI, WCE, IZZ); 
ram_4096x1 sinst_081(MDA,DBE,{AEA,AEB,AEC,AED,AEE,AEF,AEG,AEH,AEI,AEJ,AEK,AEL}, ZZI, WCE, IZZ); 
ram_4096x1 sinst_082(MFA,DCE,{AHA,AHB,AHC,AHD,AHE,AHF,AHG,AHH,AHI,AHJ,AHK,AHL}, ZZI, WCE, IZZ); 
ram_4096x1 sinst_083(MHA,DDE,{AKA,AKB,AKC,AKD,AKE,AKF,AKG,AKH,AKI,AKJ,AKK,AKL}, ZZI, WCE, IZZ); 
ram_4096x1 sinst_084(MBB,DAF,{aaa,aab,aac,aad,aae,aaf,aag,aah,aai,aaj,aak,aal}, ZZI, WCF, IZZ); 
ram_4096x1 sinst_085(MDB,DBF,{aea,aeb,aec,aed,aee,aef,aeg,aeh,aei,aej,aek,ael}, ZZI, WCF, IZZ); 
ram_4096x1 sinst_086(MFB,DCF,{aha,ahb,ahc,ahd,ahe,ahf,ahg,ahh,ahi,ahj,ahk,ahl}, ZZI, WCF, IZZ); 
ram_4096x1 sinst_087(MHB,DDF,{aka,akb,akc,akd,ake,akf,akg,akh,aki,akj,akk,akl}, ZZI, WCF, IZZ); 
ram_4096x1 sinst_088(MBC,DAG,{ABA,ABB,ABC,ABD,ABE,ABF,ABG,ABH,ABI,ABJ,ABK,ABL}, ZZI, WCG, IZZ); 
ram_4096x1 sinst_089(MDC,DBG,{AFA,AFB,AFC,AFD,AFE,AFF,AFG,AFH,AFI,AFJ,AFK,AFL}, ZZI, WCG, IZZ); 
ram_4096x1 sinst_090(MFC,DCG,{AIA,AIB,AIC,AID,AIE,AIF,AIG,AIH,AII,AIJ,AIK,AIL}, ZZI, WCG, IZZ); 
ram_4096x1 sinst_091(MHC,DDG,{ALA,ALB,ALC,ALD,ALE,ALF,ALG,ALH,ALI,ALJ,ALK,ALL}, ZZI, WCG, IZZ); 
ram_4096x1 sinst_092(MBD,DAH,{aba,abb,abc,abd,abe,abf,abg,abh,abi,abj,abk,abl}, ZZI, WCH, IZZ); 
ram_4096x1 sinst_093(MDD,DBH,{afa,afb,afc,afd,afe,aff,afg,afh,afi,afj,afk,afl}, ZZI, WCH, IZZ); 
ram_4096x1 sinst_094(MFD,DCH,{aia,aib,aic,aid,aie,aif,aig,aih,aii,aij,aik,ail}, ZZI, WCH, IZZ); 
ram_4096x1 sinst_095(MHD,DDH,{ala,alb,alc,ald,ale,alf,alg,alh,ali,alj,alk,all}, ZZI, WCH, IZZ); 
ram_4096x1 sinst_096(MBE,DAA,{AAA,AAB,AAC,AAD,AAE,AAF,AAG,AAH,AAI,AAJ,AAK,AAL}, ZZI, WDA, IZZ); 
ram_4096x1 sinst_097(MDE,DBA,{AEA,AEB,AEC,AED,AEE,AEF,AEG,AEH,AEI,AEJ,AEK,AEL}, ZZI, WDA, IZZ); 
ram_4096x1 sinst_098(MFE,DCA,{AHA,AHB,AHC,AHD,AHE,AHF,AHG,AHH,AHI,AHJ,AHK,AHL}, ZZI, WDA, IZZ); 
ram_4096x1 sinst_099(MHE,DDA,{AKA,AKB,AKC,AKD,AKE,AKF,AKG,AKH,AKI,AKJ,AKK,AKL}, ZZI, WDA, IZZ); 
ram_4096x1 sinst_100(MBF,DAB,{aaa,aab,aac,aad,aae,aaf,aag,aah,aai,aaj,aak,aal}, ZZI, WDB, IZZ); 
ram_4096x1 sinst_101(MDF,DBB,{aea,aeb,aec,aed,aee,aef,aeg,aeh,aei,aej,aek,ael}, ZZI, WDB, IZZ); 
ram_4096x1 sinst_102(MFF,DCB,{aha,ahb,ahc,ahd,ahe,ahf,ahg,ahh,ahi,ahj,ahk,ahl}, ZZI, WDB, IZZ); 
ram_4096x1 sinst_103(MHF,DDB,{aka,akb,akc,akd,ake,akf,akg,akh,aki,akj,akk,akl}, ZZI, WDB, IZZ); 
ram_4096x1 sinst_104(MBG,DAC,{ABA,ABB,ABC,ABD,ABE,ABF,ABG,ABH,ABI,ABJ,ABK,ABL}, ZZI, WDC, IZZ); 
ram_4096x1 sinst_105(MDG,DBC,{AFA,AFB,AFC,AFD,AFE,AFF,AFG,AFH,AFI,AFJ,AFK,AFL}, ZZI, WDC, IZZ); 
ram_4096x1 sinst_106(MFG,DCC,{AIA,AIB,AIC,AID,AIE,AIF,AIG,AIH,AII,AIJ,AIK,AIL}, ZZI, WDC, IZZ); 
ram_4096x1 sinst_107(MHG,DDC,{ALA,ALB,ALC,ALD,ALE,ALF,ALG,ALH,ALI,ALJ,ALK,ALL}, ZZI, WDC, IZZ); 
ram_4096x1 sinst_108(MBH,DAD,{aba,abb,abc,abd,abe,abf,abg,abh,abi,abj,abk,abl}, ZZI, WDD, IZZ); 
ram_4096x1 sinst_109(MDH,DBD,{afa,afb,afc,afd,afe,aff,afg,afh,afi,afj,afk,afl}, ZZI, WDD, IZZ); 
ram_4096x1 sinst_110(MFH,DCD,{aia,aib,aic,aid,aie,aif,aig,aih,aii,aij,aik,ail}, ZZI, WDD, IZZ); 
ram_4096x1 sinst_111(MHH,DDD,{ala,alb,alc,ald,ale,alf,alg,alh,ali,alj,alk,all}, ZZI, WDD, IZZ); 
ram_4096x1 sinst_112(MBI,DAE,{AAA,AAB,AAC,AAD,AAE,AAF,AAG,AAH,AAI,AAJ,AAK,AAL}, ZZI, WDE, IZZ); 
ram_4096x1 sinst_113(MDI,DBE,{AEA,AEB,AEC,AED,AEE,AEF,AEG,AEH,AEI,AEJ,AEK,AEL}, ZZI, WDE, IZZ); 
ram_4096x1 sinst_114(MFI,DCE,{AHA,AHB,AHC,AHD,AHE,AHF,AHG,AHH,AHI,AHJ,AHK,AHL}, ZZI, WDE, IZZ); 
ram_4096x1 sinst_115(MHI,DDE,{AKA,AKB,AKC,AKD,AKE,AKF,AKG,AKH,AKI,AKJ,AKK,AKL}, ZZI, WDE, IZZ); 
ram_4096x1 sinst_116(MBJ,DAF,{aaa,aab,aac,aad,aae,aaf,aag,aah,aai,aaj,aak,aal}, ZZI, WDF, IZZ); 
ram_4096x1 sinst_117(MDJ,DBF,{aea,aeb,aec,aed,aee,aef,aeg,aeh,aei,aej,aek,ael}, ZZI, WDF, IZZ); 
ram_4096x1 sinst_118(MFJ,DCF,{aha,ahb,ahc,ahd,ahe,ahf,ahg,ahh,ahi,ahj,ahk,ahl}, ZZI, WDF, IZZ); 
ram_4096x1 sinst_119(MHJ,DDF,{aka,akb,akc,akd,ake,akf,akg,akh,aki,akj,akk,akl}, ZZI, WDF, IZZ); 
ram_4096x1 sinst_120(MBK,DAG,{ABA,ABB,ABC,ABD,ABE,ABF,ABG,ABH,ABI,ABJ,ABK,ABL}, ZZI, WDG, IZZ); 
ram_4096x1 sinst_121(MDK,DBG,{AFA,AFB,AFC,AFD,AFE,AFF,AFG,AFH,AFI,AFJ,AFK,AFL}, ZZI, WDG, IZZ); 
ram_4096x1 sinst_122(MFK,DCG,{AIA,AIB,AIC,AID,AIE,AIF,AIG,AIH,AII,AIJ,AIK,AIL}, ZZI, WDG, IZZ); 
ram_4096x1 sinst_123(MHK,DDG,{ALA,ALB,ALC,ALD,ALE,ALF,ALG,ALH,ALI,ALJ,ALK,ALL}, ZZI, WDG, IZZ); 
ram_4096x1 sinst_124(MBL,DAH,{aba,abb,abc,abd,abe,abf,abg,abh,abi,abj,abk,abl}, ZZI, WDH, IZZ); 
ram_4096x1 sinst_125(MDL,DBH,{afa,afb,afc,afd,afe,aff,afg,afh,afi,afj,afk,afl}, ZZI, WDH, IZZ); 
ram_4096x1 sinst_126(MFL,DCH,{aia,aib,aic,aid,aie,aif,aig,aih,aii,aij,aik,ail}, ZZI, WDH, IZZ); 
ram_4096x1 sinst_127(MHL,DDH,{ala,alb,alc,ald,ale,alf,alg,alh,ali,alj,alk,all}, ZZI, WDH, IZZ); 
ram_4096x1 sinst_128(MBM,DAA,{AAA,AAB,AAC,AAD,AAE,AAF,AAG,AAH,AAI,AAJ,AAK,AAL}, ZZI, WEA, IZZ); 
ram_4096x1 sinst_129(MDM,DBA,{AEA,AEB,AEC,AED,AEE,AEF,AEG,AEH,AEI,AEJ,AEK,AEL}, ZZI, WEA, IZZ); 
ram_4096x1 sinst_130(MFM,DCA,{AHA,AHB,AHC,AHD,AHE,AHF,AHG,AHH,AHI,AHJ,AHK,AHL}, ZZI, WEA, IZZ); 
ram_4096x1 sinst_131(MHM,DDA,{AKA,AKB,AKC,AKD,AKE,AKF,AKG,AKH,AKI,AKJ,AKK,AKL}, ZZI, WEA, IZZ); 
ram_4096x1 sinst_132(MBN,DAB,{aaa,aab,aac,aad,aae,aaf,aag,aah,aai,aaj,aak,aal}, ZZI, WEB, IZZ); 
ram_4096x1 sinst_133(MDN,DBB,{aea,aeb,aec,aed,aee,aef,aeg,aeh,aei,aej,aek,ael}, ZZI, WEB, IZZ); 
ram_4096x1 sinst_134(MFN,DCB,{aha,ahb,ahc,ahd,ahe,ahf,ahg,ahh,ahi,ahj,ahk,ahl}, ZZI, WEB, IZZ); 
ram_4096x1 sinst_135(MHN,DDB,{aka,akb,akc,akd,ake,akf,akg,akh,aki,akj,akk,akl}, ZZI, WEB, IZZ); 
ram_4096x1 sinst_136(MBO,DAC,{ABA,ABB,ABC,ABD,ABE,ABF,ABG,ABH,ABI,ABJ,ABK,ABL}, ZZI, WEC, IZZ); 
ram_4096x1 sinst_137(MDO,DBC,{AFA,AFB,AFC,AFD,AFE,AFF,AFG,AFH,AFI,AFJ,AFK,AFL}, ZZI, WEC, IZZ); 
ram_4096x1 sinst_138(MFO,DCC,{AIA,AIB,AIC,AID,AIE,AIF,AIG,AIH,AII,AIJ,AIK,AIL}, ZZI, WEC, IZZ); 
ram_4096x1 sinst_139(MHO,DDC,{ALA,ALB,ALC,ALD,ALE,ALF,ALG,ALH,ALI,ALJ,ALK,ALL}, ZZI, WEC, IZZ); 
ram_4096x1 sinst_140(MBP,DAD,{aba,abb,abc,abd,abe,abf,abg,abh,abi,abj,abk,abl}, ZZI, WED, IZZ); 
ram_4096x1 sinst_141(MDP,DBD,{afa,afb,afc,afd,afe,aff,afg,afh,afi,afj,afk,afl}, ZZI, WED, IZZ); 
ram_4096x1 sinst_142(MFP,DCD,{aia,aib,aic,aid,aie,aif,aig,aih,aii,aij,aik,ail}, ZZI, WED, IZZ); 
ram_4096x1 sinst_143(MHP,DDD,{ala,alb,alc,ald,ale,alf,alg,alh,ali,alj,alk,all}, ZZI, WED, IZZ); 
ram_4096x1 sinst_144(MBQ,DAE,{AAA,AAB,AAC,AAD,AAE,AAF,AAG,AAH,AAI,AAJ,AAK,AAL}, ZZI, WEE, IZZ); 
ram_4096x1 sinst_145(MDQ,DBE,{AEA,AEB,AEC,AED,AEE,AEF,AEG,AEH,AEI,AEJ,AEK,AEL}, ZZI, WEE, IZZ); 
ram_4096x1 sinst_146(MFQ,DCE,{AHA,AHB,AHC,AHD,AHE,AHF,AHG,AHH,AHI,AHJ,AHK,AHL}, ZZI, WEE, IZZ); 
ram_4096x1 sinst_147(MHQ,DDE,{AKA,AKB,AKC,AKD,AKE,AKF,AKG,AKH,AKI,AKJ,AKK,AKL}, ZZI, WEE, IZZ); 
ram_4096x1 sinst_148(MBR,DAF,{aaa,aab,aac,aad,aae,aaf,aag,aah,aai,aaj,aak,aal}, ZZI, WEF, IZZ); 
ram_4096x1 sinst_149(MDR,DBF,{aea,aeb,aec,aed,aee,aef,aeg,aeh,aei,aej,aek,ael}, ZZI, WEF, IZZ); 
ram_4096x1 sinst_150(MFR,DCF,{aha,ahb,ahc,ahd,ahe,ahf,ahg,ahh,ahi,ahj,ahk,ahl}, ZZI, WEF, IZZ); 
ram_4096x1 sinst_151(MHR,DDF,{aka,akb,akc,akd,ake,akf,akg,akh,aki,akj,akk,akl}, ZZI, WEF, IZZ); 
ram_4096x1 sinst_152(MBS,DAG,{ABA,ABB,ABC,ABD,ABE,ABF,ABG,ABH,ABI,ABJ,ABK,ABL}, ZZI, WEG, IZZ); 
ram_4096x1 sinst_153(MDS,DBG,{AFA,AFB,AFC,AFD,AFE,AFF,AFG,AFH,AFI,AFJ,AFK,AFL}, ZZI, WEG, IZZ); 
ram_4096x1 sinst_154(MFS,DCG,{AIA,AIB,AIC,AID,AIE,AIF,AIG,AIH,AII,AIJ,AIK,AIL}, ZZI, WEG, IZZ); 
ram_4096x1 sinst_155(MHS,DDG,{ALA,ALB,ALC,ALD,ALE,ALF,ALG,ALH,ALI,ALJ,ALK,ALL}, ZZI, WEG, IZZ); 
ram_4096x1 sinst_156(MBT,DAH,{aba,abb,abc,abd,abe,abf,abg,abh,abi,abj,abk,abl}, ZZI, WEH, IZZ); 
ram_4096x1 sinst_157(MDT,DBH,{afa,afb,afc,afd,afe,aff,afg,afh,afi,afj,afk,afl}, ZZI, WEH, IZZ); 
ram_4096x1 sinst_158(MFT,DCH,{aia,aib,aic,aid,aie,aif,aig,aih,aii,aij,aik,ail}, ZZI, WEH, IZZ); 
ram_4096x1 sinst_159(MHT,DDH,{ala,alb,alc,ald,ale,alf,alg,alh,ali,alj,alk,all}, ZZI, WEH, IZZ); 
endmodule;
