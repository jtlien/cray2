module md( IZZ,
 IAA, 
 IAB, 
 IAC, 
 IAD, 
 IAE, 
 IAF, 
 IAG, 
 IAH, 
 IAI, 
 IAJ, 
 IAK, 
 IAL, 
 IAM, 
 IAN, 
 IAO, 
 IAP, 
 IAQ, 
 IAR, 
 IAS, 
 IAT, 
 IAU, 
 IAV, 
 IAW, 
 IAX, 
 IAY, 
 IAZ, 
 IBA, 
 IBB, 
 IBC, 
 IBD, 
 IBE, 
 IBF, 
 IBG, 
 IBH, 
 IBI, 
 IBJ, 
 IBK, 
 IBL, 
 IBM, 
 IBN, 
 IBO, 
 IBP, 
 IBQ, 
 IBR, 
 IBS, 
 IBT, 
 IBU, 
 IBV, 
 IBW, 
 IBX, 
 IBY, 
 IBZ, 
 ICA, 
 ICB, 
 ICC, 
 ICD, 
 ICE, 
 ICF, 
 ICG, 
 ICH, 
 ICI, 
 ICJ, 
 IIA, 
 IKA, 
 IKB, 
 IKC, 
 IKD, 
 IKE, 
 IKF, 
 IKG, 
 IKH, 
 IKI, 
 IKJ, 
 IKK, 
 IKL, 
 IKM, 
 ILA, 
 ILB, 
 ILC, 
 ILD, 
 ILE, 
 ILF, 
 ILG, 
 ILH, 
 ILI, 
 IMA, 
 IMB, 
 IMC, 
 IMD, 
 IME, 
 IMF, 
 IMG, 
 IMH, 
 INA, 
 INB, 
 INC, 
 IND, 
 IOA, 
 IOB, 
 IRA, 
 ISA, 
 ISB, 
 ISC, 
 ITA, 
 OAA, 
 OAM, 
 OBA, 
 OBM, 
 OCA, 
 OCM, 
 ODA, 
 OEA, 
 OEB, 
 OFA, 
 OFB, 
 OGA, 
 OGB, 
 OHA, 
 OHB, 
 OIA, 
 OIB, 
 OJA, 
 OJB, 
 OKA, 
 OKB, 
 OLA, 
 OLB, 
 OMA, 
 OMB, 
 ONA, 
 ONB, 
 OOA, 
 OOB, 
 OPA, 
 OPB, 
 OQA, 
 OQB, 
 ORA, 
 ORB, 
 OSA, 
 OSB, 
 OTA, 
 OTB, 
 OUA, 
 OUB, 
 OVA, 
 OVB, 
 OWA, 
 OWB, 
 OXA, 
 OXB, 
 OYA, 
 OYB, 
 OZA, 
 OZB, 
 OZM, 
OZN ); 
    
 input IZZ; 
 input IAA; 
 input IAB; 
 input IAC; 
 input IAD; 
 input IAE; 
 input IAF; 
 input IAG; 
 input IAH; 
 input IAI; 
 input IAJ; 
 input IAK; 
 input IAL; 
 input IAM; 
 input IAN; 
 input IAO; 
 input IAP; 
 input IAQ; 
 input IAR; 
 input IAS; 
 input IAT; 
 input IAU; 
 input IAV; 
 input IAW; 
 input IAX; 
 input IAY; 
 input IAZ; 
 input IBA; 
 input IBB; 
 input IBC; 
 input IBD; 
 input IBE; 
 input IBF; 
 input IBG; 
 input IBH; 
 input IBI; 
 input IBJ; 
 input IBK; 
 input IBL; 
 input IBM; 
 input IBN; 
 input IBO; 
 input IBP; 
 input IBQ; 
 input IBR; 
 input IBS; 
 input IBT; 
 input IBU; 
 input IBV; 
 input IBW; 
 input IBX; 
 input IBY; 
 input IBZ; 
 input ICA; 
 input ICB; 
 input ICC; 
 input ICD; 
 input ICE; 
 input ICF; 
 input ICG; 
 input ICH; 
 input ICI; 
 input ICJ; 
 input IIA; 
 input IKA; 
 input IKB; 
 input IKC; 
 input IKD; 
 input IKE; 
 input IKF; 
 input IKG; 
 input IKH; 
 input IKI; 
 input IKJ; 
 input IKK; 
 input IKL; 
 input IKM; 
 input ILA; 
 input ILB; 
 input ILC; 
 input ILD; 
 input ILE; 
 input ILF; 
 input ILG; 
 input ILH; 
 input ILI; 
 input IMA; 
 input IMB; 
 input IMC; 
 input IMD; 
 input IME; 
 input IMF; 
 input IMG; 
 input IMH; 
 input INA; 
 input INB; 
 input INC; 
 input IND; 
 input IOA; 
 input IOB; 
 input IRA; 
 input ISA; 
 input ISB; 
 input ISC; 
 input ITA; 
 output OAA; 
 output OAM; 
 output OBA; 
 output OBM; 
 output OCA; 
 output OCM; 
 output ODA; 
 output OEA; 
 output OEB; 
 output OFA; 
 output OFB; 
 output OGA; 
 output OGB; 
 output OHA; 
 output OHB; 
 output OIA; 
 output OIB; 
 output OJA; 
 output OJB; 
 output OKA; 
 output OKB; 
 output OLA; 
 output OLB; 
 output OMA; 
 output OMB; 
 output ONA; 
 output ONB; 
 output OOA; 
 output OOB; 
 output OPA; 
 output OPB; 
 output OQA; 
 output OQB; 
 output ORA; 
 output ORB; 
 output OSA; 
 output OSB; 
 output OTA; 
 output OTB; 
 output OUA; 
 output OUB; 
 output OVA; 
 output OVB; 
 output OWA; 
 output OWB; 
 output OXA; 
 output OXB; 
 output OYA; 
 output OYB; 
 output OZA; 
 output OZB; 
 output OZM; 
 output OZN; 
  
  
reg  CAD ;
reg  CAE ;
reg  CAF ;
reg  CAG ;
reg  CAH ;
reg  CAI ;
reg  CAJ ;
reg  CAK ;
reg  CAL ;
reg  CAM ;
reg  CAN ;
reg  CAO ;
reg  CAP ;
reg  CAQ ;
reg  CAR ;
reg  CAS ;
reg  CAT ;
reg  CAU ;
reg  CAV ;
reg  CAW ;
reg  CAX ;
reg  CAY ;
reg  CAZ ;
reg  CBC ;
reg  CBD ;
reg  CBE ;
reg  CBF ;
reg  CBG ;
reg  CBH ;
reg  CBI ;
reg  CBJ ;
reg  CBK ;
reg  CBL ;
reg  CBM ;
reg  CBN ;
reg  CBO ;
reg  CBP ;
reg  CBQ ;
reg  CBR ;
reg  CBS ;
reg  CBT ;
reg  CBU ;
reg  CBV ;
reg  CBW ;
reg  CBX ;
reg  CBY ;
reg  CBZ ;
reg  CCA ;
reg  CCB ;
reg  CCC ;
reg  CCD ;
reg  CCE ;
reg  CCF ;
reg  CCG ;
reg  CCH ;
reg  CCI ;
reg  CCJ ;
reg  CCK ;
reg  CCL ;
reg  CCM ;
reg  CCN ;
reg  CCO ;
reg  CCP ;
reg  CCQ ;
reg  CCR ;
reg  CCS ;
reg  CCT ;
reg  CCU ;
reg  CCV ;
reg  CCW ;
reg  CCX ;
reg  CCY ;
reg  CCZ ;
reg  CDB ;
reg  CDC ;
reg  cdd ;
reg  cde ;
reg  cdf ;
reg  cdg ;
reg  cdh ;
reg  cdi ;
reg  cdj ;
reg  CDK ;
reg  CDL ;
reg  CDM ;
reg  CDN ;
reg  CDO ;
reg  CDP ;
reg  CDQ ;
reg  CDR ;
reg  CDS ;
reg  CDT ;
reg  CDU ;
reg  CDV ;
reg  CDW ;
reg  CDX ;
reg  CDY ;
reg  CDZ ;
reg  DAA ;
reg  DAB ;
reg  DAC ;
reg  DAE ;
reg  DAF ;
reg  DAG ;
reg  DAI ;
reg  DAJ ;
reg  DAK ;
reg  DAM ;
reg  DAN ;
reg  DAO ;
reg  DAQ ;
reg  DAR ;
reg  DAS ;
reg  DAU ;
reg  DAV ;
reg  DAW ;
reg  DAY ;
reg  DAZ ;
reg  DBB ;
reg  DBC ;
reg  DBD ;
reg  DBF ;
reg  DBG ;
reg  DBH ;
reg  DBJ ;
reg  DBK ;
reg  DBL ;
reg  DBN ;
reg  DBO ;
reg  DBP ;
reg  DBR ;
reg  DBS ;
reg  DBT ;
reg  DBV ;
reg  DBW ;
reg  DBX ;
reg  DBZ ;
reg  DCC ;
reg  DCD ;
reg  DCE ;
reg  DCG ;
reg  DCH ;
reg  DCI ;
reg  DCK ;
reg  DCL ;
reg  DCM ;
reg  DCO ;
reg  DCP ;
reg  DCQ ;
reg  DCS ;
reg  DCT ;
reg  DCU ;
reg  DCW ;
reg  DCX ;
reg  DCY ;
reg  DCZ ;
reg  DDD ;
reg  DDE ;
reg  DDF ;
reg  DDH ;
reg  DDI ;
reg  DDJ ;
reg  DDL ;
reg  DDM ;
reg  DDN ;
reg  DDP ;
reg  DDQ ;
reg  DDR ;
reg  DDT ;
reg  DDU ;
reg  DDV ;
reg  DDX ;
reg  DDY ;
reg  DDZ ;
reg  DEM ;
reg  DEN ;
reg  DEO ;
reg  DEQ ;
reg  DER ;
reg  DES ;
reg  DEU ;
reg  DEV ;
reg  DEW ;
reg  DEY ;
reg  dez ;
reg  DFJ ;
reg  DFK ;
reg  DFL ;
reg  dfn ;
reg  dfo ;
reg  DFP ;
reg  dfr ;
reg  dfs ;
reg  DFT ;
reg  dfv ;
reg  dfw ;
reg  DFX ;
reg  dfz ;
reg  dgk ;
reg  dgl ;
reg  dgm ;
reg  dgo ;
reg  dgp ;
reg  dgq ;
reg  dgs ;
reg  dgt ;
reg  dgu ;
reg  dgw ;
reg  dgx ;
reg  dgy ;
reg  dgz ;
reg  dhl ;
reg  dhm ;
reg  dhn ;
reg  dhp ;
reg  dhq ;
reg  dhr ;
reg  dht ;
reg  dhu ;
reg  dhv ;
reg  dhx ;
reg  dhy ;
reg  dhz ;
reg  dky ;
reg  FAA ;
reg  FAB ;
reg  FAC ;
reg  FAD ;
reg  FAE ;
reg  FAF ;
reg  FAG ;
reg  FAH ;
reg  FAI ;
reg  fam ;
reg  fan ;
reg  fao ;
reg  fap ;
reg  faq ;
reg  far ;
reg  fas ;
reg  fat ;
reg  fau ;
reg  FBA ;
reg  FBB ;
reg  FBC ;
reg  FBD ;
reg  FBE ;
reg  FBF ;
reg  FBG ;
reg  FBH ;
reg  FBI ;
reg  FBJ ;
reg  fbm ;
reg  fbn ;
reg  fbo ;
reg  fbp ;
reg  fbq ;
reg  fbr ;
reg  fbs ;
reg  fbt ;
reg  FCA ;
reg  FCB ;
reg  FCC ;
reg  FCD ;
reg  FCE ;
reg  FCF ;
reg  FCG ;
reg  FCH ;
reg  FCI ;
reg  fcm ;
reg  fcn ;
reg  fco ;
reg  fcp ;
reg  fcq ;
reg  fcr ;
reg  fcs ;
reg  fct ;
reg  FDA ;
reg  FDB ;
reg  FDC ;
reg  FDD ;
reg  FDE ;
reg  FDF ;
reg  FDG ;
reg  FDH ;
reg  fdm ;
reg  fdn ;
reg  fdo ;
reg  fdp ;
reg  fdq ;
reg  fdr ;
reg  fds ;
reg  fdt ;
reg  FEA ;
reg  FEB ;
reg  FEC ;
reg  FED ;
reg  FEE ;
reg  FEF ;
reg  FEG ;
reg  FEH ;
reg  FEI ;
reg  fem ;
reg  fen ;
reg  feo ;
reg  fep ;
reg  feq ;
reg  fer ;
reg  fes ;
reg  FFA ;
reg  FFB ;
reg  FFC ;
reg  FFD ;
reg  FFE ;
reg  FFF ;
reg  FFG ;
reg  FFH ;
reg  ffm ;
reg  ffn ;
reg  ffo ;
reg  ffp ;
reg  ffq ;
reg  ffr ;
reg  ffs ;
reg  FGA ;
reg  FGB ;
reg  FGC ;
reg  FGD ;
reg  FGE ;
reg  FGF ;
reg  FGG ;
reg  fgm ;
reg  fgn ;
reg  fgo ;
reg  fgp ;
reg  fgq ;
reg  fgr ;
reg  fgs ;
reg  FHA ;
reg  FHB ;
reg  FHC ;
reg  FHD ;
reg  FHE ;
reg  FHF ;
reg  FHG ;
reg  FHH ;
reg  fhm ;
reg  fhn ;
reg  fho ;
reg  fhp ;
reg  fhq ;
reg  fhr ;
reg  FIA ;
reg  FIB ;
reg  FIC ;
reg  FID ;
reg  FIE ;
reg  FIF ;
reg  FIG ;
reg  fim ;
reg  fin ;
reg  fio ;
reg  fip ;
reg  fiq ;
reg  fir ;
reg  FJA ;
reg  FJB ;
reg  FJC ;
reg  FJD ;
reg  FJE ;
reg  FJF ;
reg  fjm ;
reg  fjn ;
reg  fjo ;
reg  fjp ;
reg  fjq ;
reg  fjr ;
reg  FKA ;
reg  FKB ;
reg  FKC ;
reg  FKD ;
reg  FKE ;
reg  FKF ;
reg  FKG ;
reg  fkm ;
reg  fkn ;
reg  fko ;
reg  fkp ;
reg  fkq ;
reg  FLA ;
reg  FLB ;
reg  FLC ;
reg  FLD ;
reg  FLE ;
reg  FLF ;
reg  flm ;
reg  fln ;
reg  flo ;
reg  flp ;
reg  flq ;
reg  FMA ;
reg  FMB ;
reg  FMC ;
reg  FMD ;
reg  FME ;
reg  fmm ;
reg  fmn ;
reg  fmo ;
reg  fmp ;
reg  fmq ;
reg  FNA ;
reg  FNB ;
reg  FNC ;
reg  FND ;
reg  FNE ;
reg  FNF ;
reg  fnm ;
reg  fnn ;
reg  fno ;
reg  fnp ;
reg  FOA ;
reg  FOB ;
reg  FOC ;
reg  FOD ;
reg  FOE ;
reg  fom ;
reg  fon ;
reg  foo ;
reg  fop ;
reg  FPA ;
reg  FPB ;
reg  FPC ;
reg  FPD ;
reg  fpm ;
reg  fpn ;
reg  fpo ;
reg  fpp ;
reg  FQA ;
reg  FQB ;
reg  FQC ;
reg  FQD ;
reg  FQE ;
reg  fqm ;
reg  fqn ;
reg  fqo ;
reg  FRA ;
reg  FRB ;
reg  FRC ;
reg  FRD ;
reg  frm ;
reg  frn ;
reg  fro ;
reg  FSA ;
reg  FSB ;
reg  FSC ;
reg  fsm ;
reg  fsn ;
reg  fso ;
reg  FTA ;
reg  FTB ;
reg  FTC ;
reg  FTD ;
reg  ftm ;
reg  ftn ;
reg  FUA ;
reg  FUB ;
reg  FUC ;
reg  fum ;
reg  fun ;
reg  FVA ;
reg  FVB ;
reg  fvm ;
reg  fvn ;
reg  FWA ;
reg  FWB ;
reg  FWC ;
reg  fwm ;
reg  FXA ;
reg  FXB ;
reg  fxm ;
reg  FYA ;
reg  fym ;
reg  FZA ;
reg  FZB ;
reg  HAA ;
reg  HAB ;
reg  HAC ;
reg  HAD ;
reg  ham ;
reg  han ;
reg  hao ;
reg  hap ;
reg  HBA ;
reg  HBB ;
reg  HBC ;
reg  HBD ;
reg  hbm ;
reg  hbn ;
reg  hbo ;
reg  HCA ;
reg  HCB ;
reg  HCC ;
reg  HCD ;
reg  HCE ;
reg  hcm ;
reg  hcn ;
reg  hco ;
reg  hcp ;
reg  HDA ;
reg  HDB ;
reg  HDC ;
reg  HDD ;
reg  HDE ;
reg  hdm ;
reg  hdn ;
reg  hdo ;
reg  HEA ;
reg  HEB ;
reg  HEC ;
reg  HED ;
reg  hem ;
reg  hen ;
reg  heo ;
reg  hep ;
reg  HFA ;
reg  HFB ;
reg  HFC ;
reg  HFD ;
reg  hfm ;
reg  hfn ;
reg  hfo ;
reg  HGA ;
reg  HGB ;
reg  HGC ;
reg  HGD ;
reg  HGE ;
reg  hgm ;
reg  hgn ;
reg  hgo ;
reg  HHA ;
reg  HHB ;
reg  HHC ;
reg  hhm ;
reg  hhn ;
reg  hho ;
reg  HIA ;
reg  HIB ;
reg  HIC ;
reg  HID ;
reg  him ;
reg  hin ;
reg  hio ;
reg  HJA ;
reg  HJB ;
reg  HJC ;
reg  HJD ;
reg  hjm ;
reg  hjn ;
reg  HKA ;
reg  HKB ;
reg  HKC ;
reg  hkm ;
reg  hkn ;
reg  hko ;
reg  HLA ;
reg  HLB ;
reg  HLC ;
reg  hlm ;
reg  hln ;
reg  hlo ;
reg  HMA ;
reg  HMB ;
reg  HMC ;
reg  hmm ;
reg  hmn ;
reg  HNA ;
reg  HNB ;
reg  HNC ;
reg  HND ;
reg  hnm ;
reg  hnn ;
reg  HOA ;
reg  HOB ;
reg  hom ;
reg  hon ;
reg  HPA ;
reg  HPB ;
reg  HPC ;
reg  hpm ;
reg  hpn ;
reg  HQA ;
reg  HQB ;
reg  HQC ;
reg  hqm ;
reg  HRA ;
reg  HRB ;
reg  hrm ;
reg  hrn ;
reg  HSA ;
reg  HSB ;
reg  hsm ;
reg  HTA ;
reg  HTB ;
reg  HTC ;
reg  htm ;
reg  HUA ;
reg  HUB ;
reg  HUC ;
reg  hum ;
reg  HVA ;
reg  hvm ;
reg  HWA ;
reg  HWB ;
reg  hwm ;
reg  HXA ;
reg  HXB ;
reg  HYA ;
reg  hym ;
reg  HZA ;
reg  HZM ;
reg  KAA ;
reg  KAB ;
reg  KAC ;
reg  KAD ;
reg  kam ;
reg  kan ;
reg  KBA ;
reg  KBB ;
reg  KBC ;
reg  kbm ;
reg  kbn ;
reg  KCA ;
reg  KCB ;
reg  kcm ;
reg  kcn ;
reg  KDA ;
reg  KDB ;
reg  KDC ;
reg  kdm ;
reg  KEA ;
reg  KEB ;
reg  kem ;
reg  ken ;
reg  KFA ;
reg  KFB ;
reg  kfm ;
reg  kfn ;
reg  KGA ;
reg  KGB ;
reg  kgm ;
reg  kgn ;
reg  KHA ;
reg  KHB ;
reg  khm ;
reg  KIA ;
reg  KIB ;
reg  KIC ;
reg  kim ;
reg  KJA ;
reg  KJB ;
reg  KJC ;
reg  kjm ;
reg  KKA ;
reg  KKB ;
reg  KKC ;
reg  kkm ;
reg  KLA ;
reg  klm ;
reg  KMA ;
reg  KMB ;
reg  kmm ;
reg  KNA ;
reg  KNB ;
reg  knm ;
reg  KOA ;
reg  KOB ;
reg  kom ;
reg  KPA ;
reg  KPB ;
reg  kpm ;
reg  KQA ;
reg  KQB ;
reg  kqm ;
reg  KRA ;
reg  KRB ;
reg  KSA ;
reg  ksm ;
reg  KTA ;
reg  ktm ;
reg  KUA ;
reg  kum ;
reg  KVA ;
reg  kvm ;
reg  KWA ;
reg  KXA ;
reg  KXB ;
reg  KYA ;
reg  KYB ;
reg  KZA ;
reg  KZB ;
reg  KZM ;
reg  MAA ;
reg  MAB ;
reg  MAC ;
reg  mam ;
reg  MBA ;
reg  MBB ;
reg  MBC ;
reg  mbm ;
reg  MCA ;
reg  mcm ;
reg  MDA ;
reg  MDB ;
reg  mdm ;
reg  MEA ;
reg  MEB ;
reg  MFA ;
reg  mfm ;
reg  MGA ;
reg  mgm ;
reg  MHA ;
reg  mhm ;
reg  MIA ;
reg  mim ;
reg  MJA ;
reg  mjm ;
reg  MKA ;
reg  mkm ;
reg  MLA ;
reg  mlm ;
reg  MMA ;
reg  MNA ;
reg  MNB ;
reg  MOA ;
reg  MOB ;
reg  MPA ;
reg  MPB ;
reg  MQA ;
reg  MQB ;
reg  MRA ;
reg  MRB ;
reg  MSA ;
reg  MSB ;
reg  MTA ;
reg  MTB ;
reg  MUA ;
reg  MUB ;
reg  MVA ;
reg  MVB ;
reg  MWA ;
reg  MWB ;
reg  MXA ;
reg  MXB ;
reg  MYA ;
reg  MYB ;
reg  MZA ;
reg  MZB ;
reg  MZM ;
reg  OAA ;
reg  oam ;
reg  OBA ;
reg  obm ;
reg  OCA ;
reg  ocm ;
reg  ODA ;
reg  OEA ;
reg  OEB ;
reg  OFA ;
reg  OFB ;
reg  OGA ;
reg  OGB ;
reg  OHA ;
reg  OHB ;
reg  OIA ;
reg  OIB ;
reg  OJA ;
reg  OJB ;
reg  OKA ;
reg  OKB ;
reg  OLA ;
reg  OLB ;
reg  OMA ;
reg  OMB ;
reg  ONA ;
reg  ONB ;
reg  OOA ;
reg  OOB ;
reg  OPA ;
reg  OPB ;
reg  OQA ;
reg  OQB ;
reg  ORA ;
reg  ORB ;
reg  OSA ;
reg  OSB ;
reg  OTA ;
reg  OTB ;
reg  OUA ;
reg  OUB ;
reg  OVA ;
reg  OVB ;
reg  OWA ;
reg  OWB ;
reg  OXA ;
reg  OXB ;
reg  OYA ;
reg  OYB ;
reg  OZA ;
reg  OZB ;
reg  OZM ;
reg  OZN ;
reg  qaa ;
reg  qab ;
reg  qac ;
reg  qad ;
reg  qae ;
reg  qaf ;
reg  qag ;
reg  qah ;
reg  qai ;
reg  qaj ;
reg  qak ;
reg  qal ;
reg  qam ;
reg  QAN ;
reg  QAO ;
reg  QAP ;
reg  QAQ ;
reg  QAR ;
reg  QAS ;
reg  QAT ;
reg  QAU ;
reg  QAV ;
reg  QAW ;
reg  QAX ;
reg  QAY ;
reg  QAZ ;
reg  QBA ;
reg  QBB ;
reg  QBC ;
reg  QBD ;
reg  QBE ;
reg  QIA ;
reg  QIB ;
reg  QIC ;
reg  QID ;
reg  QIE ;
reg  QRA ;
reg  QTA ;
reg  TRA ;
reg  TRB ;
reg  TRC ;
reg  TRD ;
reg  TRE ;
reg  TRF ;
reg  TRG ;
reg  TRH ;
reg  TTA ;
reg  TTB ;
wire  cad ;
wire  cae ;
wire  caf ;
wire  cag ;
wire  cah ;
wire  cai ;
wire  caj ;
wire  cak ;
wire  cal ;
wire  cam ;
wire  can ;
wire  cao ;
wire  cap ;
wire  caq ;
wire  car ;
wire  cas ;
wire  cat ;
wire  cau ;
wire  cav ;
wire  caw ;
wire  cax ;
wire  cay ;
wire  caz ;
wire  cbc ;
wire  cbd ;
wire  cbe ;
wire  cbf ;
wire  cbg ;
wire  cbh ;
wire  cbi ;
wire  cbj ;
wire  cbk ;
wire  cbl ;
wire  cbm ;
wire  cbn ;
wire  cbo ;
wire  cbp ;
wire  cbq ;
wire  cbr ;
wire  cbs ;
wire  cbt ;
wire  cbu ;
wire  cbv ;
wire  cbw ;
wire  cbx ;
wire  cby ;
wire  cbz ;
wire  cca ;
wire  ccb ;
wire  ccc ;
wire  ccd ;
wire  cce ;
wire  ccf ;
wire  ccg ;
wire  cch ;
wire  cci ;
wire  ccj ;
wire  cck ;
wire  ccl ;
wire  ccm ;
wire  ccn ;
wire  cco ;
wire  ccp ;
wire  ccq ;
wire  ccr ;
wire  ccs ;
wire  cct ;
wire  ccu ;
wire  ccv ;
wire  ccw ;
wire  ccx ;
wire  ccy ;
wire  ccz ;
wire  cdb ;
wire  cdc ;
wire  CDD ;
wire  CDE ;
wire  CDF ;
wire  CDG ;
wire  CDH ;
wire  CDI ;
wire  CDJ ;
wire  cdk ;
wire  cdl ;
wire  cdm ;
wire  cdn ;
wire  cdo ;
wire  cdp ;
wire  cdq ;
wire  cdr ;
wire  cds ;
wire  cdt ;
wire  cdu ;
wire  cdv ;
wire  cdw ;
wire  cdx ;
wire  cdy ;
wire  cdz ;
wire  daa ;
wire  dab ;
wire  dac ;
wire  dae ;
wire  daf ;
wire  dag ;
wire  dai ;
wire  daj ;
wire  dak ;
wire  dam ;
wire  dan ;
wire  dao ;
wire  daq ;
wire  dar ;
wire  das ;
wire  dau ;
wire  dav ;
wire  daw ;
wire  day ;
wire  daz ;
wire  dbb ;
wire  dbc ;
wire  dbd ;
wire  dbf ;
wire  dbg ;
wire  dbh ;
wire  dbj ;
wire  dbk ;
wire  dbl ;
wire  dbn ;
wire  dbo ;
wire  dbp ;
wire  dbr ;
wire  dbs ;
wire  dbt ;
wire  dbv ;
wire  dbw ;
wire  dbx ;
wire  dbz ;
wire  dcc ;
wire  dcd ;
wire  dce ;
wire  dcg ;
wire  dch ;
wire  dci ;
wire  dck ;
wire  dcl ;
wire  dcm ;
wire  dco ;
wire  dcp ;
wire  dcq ;
wire  dcs ;
wire  dct ;
wire  dcu ;
wire  dcw ;
wire  dcx ;
wire  dcy ;
wire  dcz ;
wire  ddd ;
wire  dde ;
wire  ddf ;
wire  ddh ;
wire  ddi ;
wire  ddj ;
wire  ddl ;
wire  ddm ;
wire  ddn ;
wire  ddp ;
wire  ddq ;
wire  ddr ;
wire  ddt ;
wire  ddu ;
wire  ddv ;
wire  ddx ;
wire  ddy ;
wire  ddz ;
wire  dem ;
wire  den ;
wire  deo ;
wire  deq ;
wire  der ;
wire  des ;
wire  deu ;
wire  dev ;
wire  dew ;
wire  dey ;
wire  DEZ ;
wire  dfj ;
wire  dfk ;
wire  dfl ;
wire  DFN ;
wire  DFO ;
wire  dfp ;
wire  DFR ;
wire  DFS ;
wire  dft ;
wire  DFV ;
wire  DFW ;
wire  dfx ;
wire  DFZ ;
wire  DGK ;
wire  DGL ;
wire  DGM ;
wire  DGO ;
wire  DGP ;
wire  DGQ ;
wire  DGS ;
wire  DGT ;
wire  DGU ;
wire  DGW ;
wire  DGX ;
wire  DGY ;
wire  DGZ ;
wire  DHL ;
wire  DHM ;
wire  DHN ;
wire  DHP ;
wire  DHQ ;
wire  DHR ;
wire  DHT ;
wire  DHU ;
wire  DHV ;
wire  DHX ;
wire  DHY ;
wire  DHZ ;
wire  DKY ;
wire  eaa ;
wire  EAA ;
wire  eab ;
wire  EAB ;
wire  eac ;
wire  EAC ;
wire  ead ;
wire  EAD ;
wire  eae ;
wire  EAE ;
wire  eaf ;
wire  EAF ;
wire  eag ;
wire  EAG ;
wire  eah ;
wire  EAH ;
wire  eai ;
wire  EAI ;
wire  eaj ;
wire  EAJ ;
wire  eak ;
wire  EAK ;
wire  eal ;
wire  EAL ;
wire  eam ;
wire  EAM ;
wire  ean ;
wire  EAN ;
wire  eao ;
wire  EAO ;
wire  eap ;
wire  EAP ;
wire  eaq ;
wire  EAQ ;
wire  ear ;
wire  EAR ;
wire  eas ;
wire  EAS ;
wire  eat ;
wire  EAT ;
wire  eau ;
wire  EAU ;
wire  eav ;
wire  EAV ;
wire  eaw ;
wire  EAW ;
wire  eax ;
wire  EAX ;
wire  eay ;
wire  EAY ;
wire  eaz ;
wire  EAZ ;
wire  ebb ;
wire  EBB ;
wire  ebc ;
wire  EBC ;
wire  ebd ;
wire  EBD ;
wire  ebe ;
wire  EBE ;
wire  ebf ;
wire  EBF ;
wire  ebg ;
wire  EBG ;
wire  ebh ;
wire  EBH ;
wire  ebi ;
wire  EBI ;
wire  ebj ;
wire  EBJ ;
wire  ebk ;
wire  EBK ;
wire  ebl ;
wire  EBL ;
wire  ebm ;
wire  EBM ;
wire  ebn ;
wire  EBN ;
wire  ebo ;
wire  EBO ;
wire  ebp ;
wire  EBP ;
wire  ebq ;
wire  EBQ ;
wire  ebr ;
wire  EBR ;
wire  ebs ;
wire  EBS ;
wire  ebt ;
wire  EBT ;
wire  ebu ;
wire  EBU ;
wire  ebv ;
wire  EBV ;
wire  ebw ;
wire  EBW ;
wire  ebx ;
wire  EBX ;
wire  eby ;
wire  EBY ;
wire  ebz ;
wire  EBZ ;
wire  ecc ;
wire  ECC ;
wire  ecd ;
wire  ECD ;
wire  ece ;
wire  ECE ;
wire  ecf ;
wire  ECF ;
wire  ecg ;
wire  ECG ;
wire  ech ;
wire  ECH ;
wire  eci ;
wire  ECI ;
wire  ecj ;
wire  ECJ ;
wire  eck ;
wire  ECK ;
wire  ecl ;
wire  ECL ;
wire  ecm ;
wire  ECM ;
wire  ecn ;
wire  ECN ;
wire  eco ;
wire  ECO ;
wire  ecp ;
wire  ECP ;
wire  ecq ;
wire  ECQ ;
wire  ecr ;
wire  ECR ;
wire  ecs ;
wire  ECS ;
wire  ect ;
wire  ECT ;
wire  ecu ;
wire  ECU ;
wire  ecv ;
wire  ECV ;
wire  ecw ;
wire  ECW ;
wire  ecx ;
wire  ECX ;
wire  ecy ;
wire  ECY ;
wire  ecz ;
wire  ECZ ;
wire  edd ;
wire  EDD ;
wire  ede ;
wire  EDE ;
wire  edf ;
wire  EDF ;
wire  edg ;
wire  EDG ;
wire  edh ;
wire  EDH ;
wire  edi ;
wire  EDI ;
wire  edj ;
wire  EDJ ;
wire  edk ;
wire  EDK ;
wire  edl ;
wire  EDL ;
wire  edm ;
wire  EDM ;
wire  edn ;
wire  EDN ;
wire  edo ;
wire  EDO ;
wire  edp ;
wire  EDP ;
wire  edq ;
wire  EDQ ;
wire  edr ;
wire  EDR ;
wire  eds ;
wire  EDS ;
wire  edt ;
wire  EDT ;
wire  edu ;
wire  EDU ;
wire  edv ;
wire  EDV ;
wire  edw ;
wire  EDW ;
wire  edx ;
wire  EDX ;
wire  edy ;
wire  EDY ;
wire  edz ;
wire  EDZ ;
wire  eee ;
wire  EEE ;
wire  eef ;
wire  EEF ;
wire  eeg ;
wire  EEG ;
wire  eeh ;
wire  EEH ;
wire  eei ;
wire  EEI ;
wire  eej ;
wire  EEJ ;
wire  eek ;
wire  EEK ;
wire  eel ;
wire  EEL ;
wire  eem ;
wire  EEM ;
wire  een ;
wire  EEN ;
wire  eeo ;
wire  EEO ;
wire  eep ;
wire  EEP ;
wire  eeq ;
wire  EEQ ;
wire  eer ;
wire  EER ;
wire  ees ;
wire  EES ;
wire  eet ;
wire  EET ;
wire  eeu ;
wire  EEU ;
wire  eev ;
wire  EEV ;
wire  eew ;
wire  EEW ;
wire  eex ;
wire  EEX ;
wire  eey ;
wire  EEY ;
wire  eez ;
wire  EEZ ;
wire  eff ;
wire  EFF ;
wire  efg ;
wire  EFG ;
wire  efh ;
wire  EFH ;
wire  efi ;
wire  EFI ;
wire  efj ;
wire  EFJ ;
wire  efk ;
wire  EFK ;
wire  efl ;
wire  EFL ;
wire  efm ;
wire  EFM ;
wire  efn ;
wire  EFN ;
wire  efo ;
wire  EFO ;
wire  efp ;
wire  EFP ;
wire  efq ;
wire  EFQ ;
wire  efr ;
wire  EFR ;
wire  efs ;
wire  EFS ;
wire  eft ;
wire  EFT ;
wire  efu ;
wire  EFU ;
wire  efv ;
wire  EFV ;
wire  efw ;
wire  EFW ;
wire  efx ;
wire  EFX ;
wire  efy ;
wire  EFY ;
wire  efz ;
wire  EFZ ;
wire  egg ;
wire  EGG ;
wire  egh ;
wire  EGH ;
wire  egi ;
wire  EGI ;
wire  egj ;
wire  EGJ ;
wire  egk ;
wire  EGK ;
wire  egl ;
wire  EGL ;
wire  egm ;
wire  EGM ;
wire  egn ;
wire  EGN ;
wire  ego ;
wire  EGO ;
wire  egp ;
wire  EGP ;
wire  egq ;
wire  EGQ ;
wire  egr ;
wire  EGR ;
wire  egs ;
wire  EGS ;
wire  egt ;
wire  EGT ;
wire  egu ;
wire  EGU ;
wire  egv ;
wire  EGV ;
wire  egw ;
wire  EGW ;
wire  egx ;
wire  EGX ;
wire  egy ;
wire  EGY ;
wire  egz ;
wire  EGZ ;
wire  ehh ;
wire  EHH ;
wire  ehi ;
wire  EHI ;
wire  ehj ;
wire  EHJ ;
wire  ehk ;
wire  EHK ;
wire  ehl ;
wire  EHL ;
wire  ehm ;
wire  EHM ;
wire  ehn ;
wire  EHN ;
wire  eho ;
wire  EHO ;
wire  ehp ;
wire  EHP ;
wire  ehq ;
wire  EHQ ;
wire  ehr ;
wire  EHR ;
wire  ehs ;
wire  EHS ;
wire  eht ;
wire  EHT ;
wire  ehu ;
wire  EHU ;
wire  ehv ;
wire  EHV ;
wire  ehw ;
wire  EHW ;
wire  ehx ;
wire  EHX ;
wire  ehy ;
wire  EHY ;
wire  ehz ;
wire  EHZ ;
wire  eii ;
wire  EII ;
wire  eij ;
wire  EIJ ;
wire  eik ;
wire  EIK ;
wire  eil ;
wire  EIL ;
wire  eim ;
wire  EIM ;
wire  ein ;
wire  EIN ;
wire  eio ;
wire  EIO ;
wire  eip ;
wire  EIP ;
wire  eiq ;
wire  EIQ ;
wire  eir ;
wire  EIR ;
wire  eis ;
wire  EIS ;
wire  eit ;
wire  EIT ;
wire  eiu ;
wire  EIU ;
wire  eiv ;
wire  EIV ;
wire  eiw ;
wire  EIW ;
wire  eix ;
wire  EIX ;
wire  eiy ;
wire  EIY ;
wire  eiz ;
wire  EIZ ;
wire  ejj ;
wire  EJJ ;
wire  ejk ;
wire  EJK ;
wire  ejl ;
wire  EJL ;
wire  ejm ;
wire  EJM ;
wire  ejn ;
wire  EJN ;
wire  ejo ;
wire  EJO ;
wire  ejp ;
wire  EJP ;
wire  ejq ;
wire  EJQ ;
wire  ejr ;
wire  EJR ;
wire  ejs ;
wire  EJS ;
wire  ejt ;
wire  EJT ;
wire  eju ;
wire  EJU ;
wire  ejv ;
wire  EJV ;
wire  ejw ;
wire  EJW ;
wire  ejx ;
wire  EJX ;
wire  ejy ;
wire  EJY ;
wire  ejz ;
wire  EJZ ;
wire  ekk ;
wire  EKK ;
wire  ekl ;
wire  EKL ;
wire  ekm ;
wire  EKM ;
wire  ekn ;
wire  EKN ;
wire  eko ;
wire  EKO ;
wire  ekp ;
wire  EKP ;
wire  ekq ;
wire  EKQ ;
wire  ekr ;
wire  EKR ;
wire  eks ;
wire  EKS ;
wire  ekt ;
wire  EKT ;
wire  eku ;
wire  EKU ;
wire  ekv ;
wire  EKV ;
wire  ekw ;
wire  EKW ;
wire  ekx ;
wire  EKX ;
wire  eky ;
wire  EKY ;
wire  ekz ;
wire  EKZ ;
wire  ell ;
wire  ELL ;
wire  elm ;
wire  ELM ;
wire  eln ;
wire  ELN ;
wire  elo ;
wire  ELO ;
wire  elp ;
wire  ELP ;
wire  elq ;
wire  ELQ ;
wire  elr ;
wire  ELR ;
wire  els ;
wire  ELS ;
wire  elt ;
wire  ELT ;
wire  elu ;
wire  ELU ;
wire  elv ;
wire  ELV ;
wire  elw ;
wire  ELW ;
wire  elx ;
wire  ELX ;
wire  ely ;
wire  ELY ;
wire  elz ;
wire  ELZ ;
wire  emm ;
wire  EMM ;
wire  emn ;
wire  EMN ;
wire  emo ;
wire  EMO ;
wire  emp ;
wire  EMP ;
wire  emq ;
wire  EMQ ;
wire  emr ;
wire  EMR ;
wire  ems ;
wire  EMS ;
wire  emt ;
wire  EMT ;
wire  emu ;
wire  EMU ;
wire  emv ;
wire  EMV ;
wire  emw ;
wire  EMW ;
wire  emx ;
wire  EMX ;
wire  emy ;
wire  EMY ;
wire  emz ;
wire  EMZ ;
wire  enn ;
wire  ENN ;
wire  eno ;
wire  ENO ;
wire  enp ;
wire  ENP ;
wire  enq ;
wire  ENQ ;
wire  enr ;
wire  ENR ;
wire  ens ;
wire  ENS ;
wire  ent ;
wire  ENT ;
wire  enu ;
wire  ENU ;
wire  env ;
wire  ENV ;
wire  enw ;
wire  ENW ;
wire  enx ;
wire  ENX ;
wire  eny ;
wire  ENY ;
wire  enz ;
wire  ENZ ;
wire  eoo ;
wire  EOO ;
wire  eop ;
wire  EOP ;
wire  eoq ;
wire  EOQ ;
wire  eor ;
wire  EOR ;
wire  eos ;
wire  EOS ;
wire  eot ;
wire  EOT ;
wire  eou ;
wire  EOU ;
wire  eov ;
wire  EOV ;
wire  eow ;
wire  EOW ;
wire  eox ;
wire  EOX ;
wire  eoy ;
wire  EOY ;
wire  eoz ;
wire  EOZ ;
wire  epp ;
wire  EPP ;
wire  epq ;
wire  EPQ ;
wire  epr ;
wire  EPR ;
wire  eps ;
wire  EPS ;
wire  ept ;
wire  EPT ;
wire  epu ;
wire  EPU ;
wire  epv ;
wire  EPV ;
wire  epw ;
wire  EPW ;
wire  epx ;
wire  EPX ;
wire  epy ;
wire  EPY ;
wire  epz ;
wire  EPZ ;
wire  eqq ;
wire  EQQ ;
wire  eqr ;
wire  EQR ;
wire  eqs ;
wire  EQS ;
wire  eqt ;
wire  EQT ;
wire  equ ;
wire  EQU ;
wire  eqv ;
wire  EQV ;
wire  eqw ;
wire  EQW ;
wire  eqx ;
wire  EQX ;
wire  eqy ;
wire  EQY ;
wire  eqz ;
wire  EQZ ;
wire  err ;
wire  ERR ;
wire  ers ;
wire  ERS ;
wire  ert ;
wire  ERT ;
wire  eru ;
wire  ERU ;
wire  erv ;
wire  ERV ;
wire  erw ;
wire  ERW ;
wire  erx ;
wire  ERX ;
wire  ery ;
wire  ERY ;
wire  erz ;
wire  ERZ ;
wire  ess ;
wire  ESS ;
wire  est ;
wire  EST ;
wire  esu ;
wire  ESU ;
wire  esv ;
wire  ESV ;
wire  esw ;
wire  ESW ;
wire  esx ;
wire  ESX ;
wire  esy ;
wire  ESY ;
wire  esz ;
wire  ESZ ;
wire  ett ;
wire  ETT ;
wire  etu ;
wire  ETU ;
wire  etv ;
wire  ETV ;
wire  etw ;
wire  ETW ;
wire  etx ;
wire  ETX ;
wire  ety ;
wire  ETY ;
wire  etz ;
wire  ETZ ;
wire  euu ;
wire  EUU ;
wire  euv ;
wire  EUV ;
wire  euw ;
wire  EUW ;
wire  eux ;
wire  EUX ;
wire  euy ;
wire  EUY ;
wire  euz ;
wire  EUZ ;
wire  evv ;
wire  EVV ;
wire  evw ;
wire  EVW ;
wire  evx ;
wire  EVX ;
wire  evy ;
wire  EVY ;
wire  evz ;
wire  EVZ ;
wire  eww ;
wire  EWW ;
wire  ewx ;
wire  EWX ;
wire  ewy ;
wire  EWY ;
wire  ewz ;
wire  EWZ ;
wire  exx ;
wire  EXX ;
wire  exy ;
wire  EXY ;
wire  exz ;
wire  EXZ ;
wire  eyy ;
wire  EYY ;
wire  eyz ;
wire  EYZ ;
wire  ezz ;
wire  EZZ ;
wire  faa ;
wire  fab ;
wire  fac ;
wire  fad ;
wire  fae ;
wire  faf ;
wire  fag ;
wire  fah ;
wire  fai ;
wire  FAM ;
wire  FAN ;
wire  FAO ;
wire  FAP ;
wire  FAQ ;
wire  FAR ;
wire  FAS ;
wire  FAT ;
wire  FAU ;
wire  fba ;
wire  fbb ;
wire  fbc ;
wire  fbd ;
wire  fbe ;
wire  fbf ;
wire  fbg ;
wire  fbh ;
wire  fbi ;
wire  fbj ;
wire  FBM ;
wire  FBN ;
wire  FBO ;
wire  FBP ;
wire  FBQ ;
wire  FBR ;
wire  FBS ;
wire  FBT ;
wire  fca ;
wire  fcb ;
wire  fcc ;
wire  fcd ;
wire  fce ;
wire  fcf ;
wire  fcg ;
wire  fch ;
wire  fci ;
wire  FCM ;
wire  FCN ;
wire  FCO ;
wire  FCP ;
wire  FCQ ;
wire  FCR ;
wire  FCS ;
wire  FCT ;
wire  fda ;
wire  fdb ;
wire  fdc ;
wire  fdd ;
wire  fde ;
wire  fdf ;
wire  fdg ;
wire  fdh ;
wire  FDM ;
wire  FDN ;
wire  FDO ;
wire  FDP ;
wire  FDQ ;
wire  FDR ;
wire  FDS ;
wire  FDT ;
wire  fea ;
wire  feb ;
wire  fec ;
wire  fed ;
wire  fee ;
wire  fef ;
wire  feg ;
wire  feh ;
wire  fei ;
wire  FEM ;
wire  FEN ;
wire  FEO ;
wire  FEP ;
wire  FEQ ;
wire  FER ;
wire  FES ;
wire  ffa ;
wire  ffb ;
wire  ffc ;
wire  ffd ;
wire  ffe ;
wire  fff ;
wire  ffg ;
wire  ffh ;
wire  FFM ;
wire  FFN ;
wire  FFO ;
wire  FFP ;
wire  FFQ ;
wire  FFR ;
wire  FFS ;
wire  fga ;
wire  fgb ;
wire  fgc ;
wire  fgd ;
wire  fge ;
wire  fgf ;
wire  fgg ;
wire  FGM ;
wire  FGN ;
wire  FGO ;
wire  FGP ;
wire  FGQ ;
wire  FGR ;
wire  FGS ;
wire  fha ;
wire  fhb ;
wire  fhc ;
wire  fhd ;
wire  fhe ;
wire  fhf ;
wire  fhg ;
wire  fhh ;
wire  FHM ;
wire  FHN ;
wire  FHO ;
wire  FHP ;
wire  FHQ ;
wire  FHR ;
wire  fia ;
wire  fib ;
wire  fic ;
wire  fid ;
wire  fie ;
wire  fif ;
wire  fig ;
wire  FIM ;
wire  FIN ;
wire  FIO ;
wire  FIP ;
wire  FIQ ;
wire  FIR ;
wire  fja ;
wire  fjb ;
wire  fjc ;
wire  fjd ;
wire  fje ;
wire  fjf ;
wire  FJM ;
wire  FJN ;
wire  FJO ;
wire  FJP ;
wire  FJQ ;
wire  FJR ;
wire  fka ;
wire  fkb ;
wire  fkc ;
wire  fkd ;
wire  fke ;
wire  fkf ;
wire  fkg ;
wire  FKM ;
wire  FKN ;
wire  FKO ;
wire  FKP ;
wire  FKQ ;
wire  fla ;
wire  flb ;
wire  flc ;
wire  fld ;
wire  fle ;
wire  flf ;
wire  FLM ;
wire  FLN ;
wire  FLO ;
wire  FLP ;
wire  FLQ ;
wire  fma ;
wire  fmb ;
wire  fmc ;
wire  fmd ;
wire  fme ;
wire  FMM ;
wire  FMN ;
wire  FMO ;
wire  FMP ;
wire  FMQ ;
wire  fna ;
wire  fnb ;
wire  fnc ;
wire  fnd ;
wire  fne ;
wire  fnf ;
wire  FNM ;
wire  FNN ;
wire  FNO ;
wire  FNP ;
wire  foa ;
wire  fob ;
wire  foc ;
wire  fod ;
wire  foe ;
wire  FOM ;
wire  FON ;
wire  FOO ;
wire  FOP ;
wire  fpa ;
wire  fpb ;
wire  fpc ;
wire  fpd ;
wire  FPM ;
wire  FPN ;
wire  FPO ;
wire  FPP ;
wire  fqa ;
wire  fqb ;
wire  fqc ;
wire  fqd ;
wire  fqe ;
wire  FQM ;
wire  FQN ;
wire  FQO ;
wire  fra ;
wire  frb ;
wire  frc ;
wire  frd ;
wire  FRM ;
wire  FRN ;
wire  FRO ;
wire  fsa ;
wire  fsb ;
wire  fsc ;
wire  FSM ;
wire  FSN ;
wire  FSO ;
wire  fta ;
wire  ftb ;
wire  ftc ;
wire  ftd ;
wire  FTM ;
wire  FTN ;
wire  fua ;
wire  fub ;
wire  fuc ;
wire  FUM ;
wire  FUN ;
wire  fva ;
wire  fvb ;
wire  FVM ;
wire  FVN ;
wire  fwa ;
wire  fwb ;
wire  fwc ;
wire  FWM ;
wire  fxa ;
wire  fxb ;
wire  FXM ;
wire  fya ;
wire  FYM ;
wire  fza ;
wire  fzb ;
wire  gaa ;
wire  GAA ;
wire  gab ;
wire  GAB ;
wire  gac ;
wire  GAC ;
wire  gam ;
wire  GAM ;
wire  gan ;
wire  GAN ;
wire  gao ;
wire  GAO ;
wire  gba ;
wire  GBA ;
wire  gbb ;
wire  GBB ;
wire  gbc ;
wire  GBC ;
wire  gbd ;
wire  GBD ;
wire  gbe ;
wire  GBE ;
wire  gbf ;
wire  GBF ;
wire  gbm ;
wire  GBM ;
wire  gbn ;
wire  GBN ;
wire  gbo ;
wire  GBO ;
wire  gbp ;
wire  GBP ;
wire  gbq ;
wire  GBQ ;
wire  gbr ;
wire  GBR ;
wire  gca ;
wire  GCA ;
wire  gcb ;
wire  GCB ;
wire  gcc ;
wire  GCC ;
wire  gcd ;
wire  GCD ;
wire  gce ;
wire  GCE ;
wire  gcm ;
wire  GCM ;
wire  gcn ;
wire  GCN ;
wire  gco ;
wire  GCO ;
wire  gcp ;
wire  GCP ;
wire  gcq ;
wire  GCQ ;
wire  gda ;
wire  GDA ;
wire  gdb ;
wire  GDB ;
wire  gdc ;
wire  GDC ;
wire  gdd ;
wire  GDD ;
wire  gde ;
wire  GDE ;
wire  gdm ;
wire  GDM ;
wire  gdn ;
wire  GDN ;
wire  gdo ;
wire  GDO ;
wire  gdp ;
wire  GDP ;
wire  gdq ;
wire  GDQ ;
wire  gea ;
wire  GEA ;
wire  geb ;
wire  GEB ;
wire  gec ;
wire  GEC ;
wire  ged ;
wire  GED ;
wire  gee ;
wire  GEE ;
wire  gem ;
wire  GEM ;
wire  gen ;
wire  GEN ;
wire  geo ;
wire  GEO ;
wire  gep ;
wire  GEP ;
wire  geq ;
wire  GEQ ;
wire  gfa ;
wire  GFA ;
wire  gfb ;
wire  GFB ;
wire  gfc ;
wire  GFC ;
wire  gfd ;
wire  GFD ;
wire  gfe ;
wire  GFE ;
wire  gfm ;
wire  GFM ;
wire  gfn ;
wire  GFN ;
wire  gfo ;
wire  GFO ;
wire  gfp ;
wire  GFP ;
wire  gfq ;
wire  GFQ ;
wire  gga ;
wire  GGA ;
wire  ggb ;
wire  GGB ;
wire  ggc ;
wire  GGC ;
wire  ggd ;
wire  GGD ;
wire  ggm ;
wire  GGM ;
wire  ggn ;
wire  GGN ;
wire  ggo ;
wire  GGO ;
wire  ggp ;
wire  GGP ;
wire  gha ;
wire  GHA ;
wire  ghb ;
wire  GHB ;
wire  ghc ;
wire  GHC ;
wire  ghd ;
wire  GHD ;
wire  ghe ;
wire  GHE ;
wire  ghm ;
wire  GHM ;
wire  ghn ;
wire  GHN ;
wire  gho ;
wire  GHO ;
wire  ghp ;
wire  GHP ;
wire  ghq ;
wire  GHQ ;
wire  gia ;
wire  GIA ;
wire  gib ;
wire  GIB ;
wire  gic ;
wire  GIC ;
wire  gid ;
wire  GID ;
wire  gim ;
wire  GIM ;
wire  gin ;
wire  GIN ;
wire  gio ;
wire  GIO ;
wire  gip ;
wire  GIP ;
wire  gja ;
wire  GJA ;
wire  gjb ;
wire  GJB ;
wire  gjc ;
wire  GJC ;
wire  gjd ;
wire  GJD ;
wire  gjm ;
wire  GJM ;
wire  gjn ;
wire  GJN ;
wire  gjo ;
wire  GJO ;
wire  gjp ;
wire  GJP ;
wire  gka ;
wire  GKA ;
wire  gkb ;
wire  GKB ;
wire  gkc ;
wire  GKC ;
wire  gkd ;
wire  GKD ;
wire  gkm ;
wire  GKM ;
wire  gkn ;
wire  GKN ;
wire  gko ;
wire  GKO ;
wire  gkp ;
wire  GKP ;
wire  gla ;
wire  GLA ;
wire  glb ;
wire  GLB ;
wire  glc ;
wire  GLC ;
wire  glm ;
wire  GLM ;
wire  gln ;
wire  GLN ;
wire  glo ;
wire  GLO ;
wire  gma ;
wire  GMA ;
wire  gmb ;
wire  GMB ;
wire  gmc ;
wire  GMC ;
wire  gmm ;
wire  GMM ;
wire  gmn ;
wire  GMN ;
wire  gmo ;
wire  GMO ;
wire  gna ;
wire  GNA ;
wire  gnb ;
wire  GNB ;
wire  gnc ;
wire  GNC ;
wire  gnm ;
wire  GNM ;
wire  gnn ;
wire  GNN ;
wire  gno ;
wire  GNO ;
wire  goa ;
wire  GOA ;
wire  gob ;
wire  GOB ;
wire  goc ;
wire  GOC ;
wire  gom ;
wire  GOM ;
wire  gon ;
wire  GON ;
wire  goo ;
wire  GOO ;
wire  gpa ;
wire  GPA ;
wire  gpb ;
wire  GPB ;
wire  gpm ;
wire  GPM ;
wire  gpn ;
wire  GPN ;
wire  gqa ;
wire  GQA ;
wire  gqb ;
wire  GQB ;
wire  gqc ;
wire  GQC ;
wire  gqm ;
wire  GQM ;
wire  gqn ;
wire  GQN ;
wire  gqo ;
wire  GQO ;
wire  gra ;
wire  GRA ;
wire  grb ;
wire  GRB ;
wire  grm ;
wire  GRM ;
wire  grn ;
wire  GRN ;
wire  gsa ;
wire  GSA ;
wire  gsb ;
wire  GSB ;
wire  gsm ;
wire  GSM ;
wire  gsn ;
wire  GSN ;
wire  gta ;
wire  GTA ;
wire  gtb ;
wire  GTB ;
wire  gtm ;
wire  GTM ;
wire  gtn ;
wire  GTN ;
wire  gua ;
wire  GUA ;
wire  gum ;
wire  GUM ;
wire  gva ;
wire  GVA ;
wire  gvm ;
wire  GVM ;
wire  gwa ;
wire  GWA ;
wire  gwm ;
wire  GWM ;
wire  gxa ;
wire  GXA ;
wire  gxm ;
wire  GXM ;
wire  gza ;
wire  GZA ;
wire  gzm ;
wire  GZM ;
wire  haa ;
wire  hab ;
wire  hac ;
wire  had ;
wire  HAM ;
wire  HAN ;
wire  HAO ;
wire  HAP ;
wire  hba ;
wire  hbb ;
wire  hbc ;
wire  hbd ;
wire  HBM ;
wire  HBN ;
wire  HBO ;
wire  hca ;
wire  hcb ;
wire  hcc ;
wire  hcd ;
wire  hce ;
wire  HCM ;
wire  HCN ;
wire  HCO ;
wire  HCP ;
wire  hda ;
wire  hdb ;
wire  hdc ;
wire  hdd ;
wire  hde ;
wire  HDM ;
wire  HDN ;
wire  HDO ;
wire  hea ;
wire  heb ;
wire  hec ;
wire  hed ;
wire  HEM ;
wire  HEN ;
wire  HEO ;
wire  HEP ;
wire  hfa ;
wire  hfb ;
wire  hfc ;
wire  hfd ;
wire  HFM ;
wire  HFN ;
wire  HFO ;
wire  hga ;
wire  hgb ;
wire  hgc ;
wire  hgd ;
wire  hge ;
wire  HGM ;
wire  HGN ;
wire  HGO ;
wire  hha ;
wire  hhb ;
wire  hhc ;
wire  HHM ;
wire  HHN ;
wire  HHO ;
wire  hia ;
wire  hib ;
wire  hic ;
wire  hid ;
wire  HIM ;
wire  HIN ;
wire  HIO ;
wire  hja ;
wire  hjb ;
wire  hjc ;
wire  hjd ;
wire  HJM ;
wire  HJN ;
wire  hka ;
wire  hkb ;
wire  hkc ;
wire  HKM ;
wire  HKN ;
wire  HKO ;
wire  hla ;
wire  hlb ;
wire  hlc ;
wire  HLM ;
wire  HLN ;
wire  HLO ;
wire  hma ;
wire  hmb ;
wire  hmc ;
wire  HMM ;
wire  HMN ;
wire  hna ;
wire  hnb ;
wire  hnc ;
wire  hnd ;
wire  HNM ;
wire  HNN ;
wire  hoa ;
wire  hob ;
wire  HOM ;
wire  HON ;
wire  hpa ;
wire  hpb ;
wire  hpc ;
wire  HPM ;
wire  HPN ;
wire  hqa ;
wire  hqb ;
wire  hqc ;
wire  HQM ;
wire  hra ;
wire  hrb ;
wire  HRM ;
wire  HRN ;
wire  hsa ;
wire  hsb ;
wire  HSM ;
wire  hta ;
wire  htb ;
wire  htc ;
wire  HTM ;
wire  hua ;
wire  hub ;
wire  huc ;
wire  HUM ;
wire  hva ;
wire  HVM ;
wire  hwa ;
wire  hwb ;
wire  HWM ;
wire  hxa ;
wire  hxb ;
wire  hya ;
wire  HYM ;
wire  hza ;
wire  hzm ;
wire  iaa ;
wire  iab ;
wire  iac ;
wire  iad ;
wire  iae ;
wire  iaf ;
wire  iag ;
wire  iah ;
wire  iai ;
wire  iaj ;
wire  iak ;
wire  ial ;
wire  iam ;
wire  ian ;
wire  iao ;
wire  iap ;
wire  iaq ;
wire  iar ;
wire  ias ;
wire  iat ;
wire  iau ;
wire  iav ;
wire  iaw ;
wire  iax ;
wire  iay ;
wire  iaz ;
wire  iba ;
wire  ibb ;
wire  ibc ;
wire  ibd ;
wire  ibe ;
wire  ibf ;
wire  ibg ;
wire  ibh ;
wire  ibi ;
wire  ibj ;
wire  ibk ;
wire  ibl ;
wire  ibm ;
wire  ibn ;
wire  ibo ;
wire  ibp ;
wire  ibq ;
wire  ibr ;
wire  ibs ;
wire  ibt ;
wire  ibu ;
wire  ibv ;
wire  ibw ;
wire  ibx ;
wire  iby ;
wire  ibz ;
wire  ica ;
wire  icb ;
wire  icc ;
wire  icd ;
wire  ice ;
wire  icf ;
wire  icg ;
wire  ich ;
wire  ici ;
wire  icj ;
wire  iia ;
wire  ika ;
wire  ikb ;
wire  ikc ;
wire  ikd ;
wire  ike ;
wire  ikf ;
wire  ikg ;
wire  ikh ;
wire  iki ;
wire  ikj ;
wire  ikk ;
wire  ikl ;
wire  ikm ;
wire  ila ;
wire  ilb ;
wire  ilc ;
wire  ild ;
wire  ile ;
wire  ilf ;
wire  ilg ;
wire  ilh ;
wire  ili ;
wire  ima ;
wire  imb ;
wire  imc ;
wire  imd ;
wire  ime ;
wire  imf ;
wire  img ;
wire  imh ;
wire  ina ;
wire  inb ;
wire  inc ;
wire  ind ;
wire  ioa ;
wire  iob ;
wire  ira ;
wire  isa ;
wire  isb ;
wire  isc ;
wire  ita ;
wire  jaa ;
wire  JAA ;
wire  jam ;
wire  JAM ;
wire  jba ;
wire  JBA ;
wire  jbb ;
wire  JBB ;
wire  jbm ;
wire  JBM ;
wire  jbn ;
wire  JBN ;
wire  jca ;
wire  JCA ;
wire  jcb ;
wire  JCB ;
wire  jcm ;
wire  JCM ;
wire  jcn ;
wire  JCN ;
wire  jda ;
wire  JDA ;
wire  jdb ;
wire  JDB ;
wire  jdc ;
wire  JDC ;
wire  jdm ;
wire  JDM ;
wire  jdn ;
wire  JDN ;
wire  jdo ;
wire  JDO ;
wire  jea ;
wire  JEA ;
wire  jeb ;
wire  JEB ;
wire  jem ;
wire  JEM ;
wire  jen ;
wire  JEN ;
wire  jfa ;
wire  JFA ;
wire  jfb ;
wire  JFB ;
wire  jfm ;
wire  JFM ;
wire  jfn ;
wire  JFN ;
wire  jga ;
wire  JGA ;
wire  jgb ;
wire  JGB ;
wire  jgm ;
wire  JGM ;
wire  jgn ;
wire  JGN ;
wire  jha ;
wire  JHA ;
wire  jhb ;
wire  JHB ;
wire  jhm ;
wire  JHM ;
wire  jhn ;
wire  JHN ;
wire  jia ;
wire  JIA ;
wire  jib ;
wire  JIB ;
wire  jim ;
wire  JIM ;
wire  jin ;
wire  JIN ;
wire  jja ;
wire  JJA ;
wire  jjb ;
wire  JJB ;
wire  jjm ;
wire  JJM ;
wire  jjn ;
wire  JJN ;
wire  jka ;
wire  JKA ;
wire  jkm ;
wire  JKM ;
wire  jla ;
wire  JLA ;
wire  jlb ;
wire  JLB ;
wire  jlm ;
wire  JLM ;
wire  jln ;
wire  JLN ;
wire  jma ;
wire  JMA ;
wire  jmb ;
wire  JMB ;
wire  jmm ;
wire  JMM ;
wire  jmn ;
wire  JMN ;
wire  jna ;
wire  JNA ;
wire  jnb ;
wire  JNB ;
wire  jnm ;
wire  JNM ;
wire  jnn ;
wire  JNN ;
wire  joa ;
wire  JOA ;
wire  jom ;
wire  JOM ;
wire  jpa ;
wire  JPA ;
wire  jpm ;
wire  JPM ;
wire  jqa ;
wire  JQA ;
wire  jqm ;
wire  JQM ;
wire  jra ;
wire  JRA ;
wire  jrm ;
wire  JRM ;
wire  jsa ;
wire  JSA ;
wire  jsm ;
wire  JSM ;
wire  jta ;
wire  JTA ;
wire  jtm ;
wire  JTM ;
wire  jua ;
wire  JUA ;
wire  jum ;
wire  JUM ;
wire  jwa ;
wire  JWA ;
wire  jwm ;
wire  JWM ;
wire  jxa ;
wire  JXA ;
wire  jxm ;
wire  JXM ;
wire  kaa ;
wire  kab ;
wire  kac ;
wire  kad ;
wire  KAM ;
wire  KAN ;
wire  kba ;
wire  kbb ;
wire  kbc ;
wire  KBM ;
wire  KBN ;
wire  kca ;
wire  kcb ;
wire  KCM ;
wire  KCN ;
wire  kda ;
wire  kdb ;
wire  kdc ;
wire  KDM ;
wire  kea ;
wire  keb ;
wire  KEM ;
wire  KEN ;
wire  kfa ;
wire  kfb ;
wire  KFM ;
wire  KFN ;
wire  kga ;
wire  kgb ;
wire  KGM ;
wire  KGN ;
wire  kha ;
wire  khb ;
wire  KHM ;
wire  kia ;
wire  kib ;
wire  kic ;
wire  KIM ;
wire  kja ;
wire  kjb ;
wire  kjc ;
wire  KJM ;
wire  kka ;
wire  kkb ;
wire  kkc ;
wire  KKM ;
wire  kla ;
wire  KLM ;
wire  kma ;
wire  kmb ;
wire  KMM ;
wire  kna ;
wire  knb ;
wire  KNM ;
wire  koa ;
wire  kob ;
wire  KOM ;
wire  kpa ;
wire  kpb ;
wire  KPM ;
wire  kqa ;
wire  kqb ;
wire  KQM ;
wire  kra ;
wire  krb ;
wire  ksa ;
wire  KSM ;
wire  kta ;
wire  KTM ;
wire  kua ;
wire  KUM ;
wire  kva ;
wire  KVM ;
wire  kwa ;
wire  kxa ;
wire  kxb ;
wire  kya ;
wire  kyb ;
wire  kza ;
wire  kzb ;
wire  kzm ;
wire  laa ;
wire  LAA ;
wire  lam ;
wire  LAM ;
wire  lba ;
wire  LBA ;
wire  lbm ;
wire  LBM ;
wire  lca ;
wire  LCA ;
wire  lcm ;
wire  LCM ;
wire  lda ;
wire  LDA ;
wire  ldm ;
wire  LDM ;
wire  lea ;
wire  LEA ;
wire  lem ;
wire  LEM ;
wire  lfa ;
wire  LFA ;
wire  lfm ;
wire  LFM ;
wire  lga ;
wire  LGA ;
wire  lgm ;
wire  LGM ;
wire  lha ;
wire  LHA ;
wire  lhm ;
wire  LHM ;
wire  lia ;
wire  LIA ;
wire  lim ;
wire  LIM ;
wire  lja ;
wire  LJA ;
wire  ljm ;
wire  LJM ;
wire  lka ;
wire  LKA ;
wire  lkm ;
wire  LKM ;
wire  lma ;
wire  LMA ;
wire  lmm ;
wire  LMM ;
wire  lna ;
wire  LNA ;
wire  lnm ;
wire  LNM ;
wire  loa ;
wire  LOA ;
wire  lom ;
wire  LOM ;
wire  lpa ;
wire  LPA ;
wire  lpm ;
wire  LPM ;
wire  lqa ;
wire  LQA ;
wire  lqm ;
wire  LQM ;
wire  lra ;
wire  LRA ;
wire  lrm ;
wire  LRM ;
wire  maa ;
wire  mab ;
wire  mac ;
wire  MAM ;
wire  mba ;
wire  mbb ;
wire  mbc ;
wire  MBM ;
wire  mca ;
wire  MCM ;
wire  mda ;
wire  mdb ;
wire  MDM ;
wire  mea ;
wire  meb ;
wire  mfa ;
wire  MFM ;
wire  mga ;
wire  MGM ;
wire  mha ;
wire  MHM ;
wire  mia ;
wire  MIM ;
wire  mja ;
wire  MJM ;
wire  mka ;
wire  MKM ;
wire  mla ;
wire  MLM ;
wire  mma ;
wire  mna ;
wire  mnb ;
wire  moa ;
wire  mob ;
wire  mpa ;
wire  mpb ;
wire  mqa ;
wire  mqb ;
wire  mra ;
wire  mrb ;
wire  msa ;
wire  msb ;
wire  mta ;
wire  mtb ;
wire  mua ;
wire  mub ;
wire  mva ;
wire  mvb ;
wire  mwa ;
wire  mwb ;
wire  mxa ;
wire  mxb ;
wire  mya ;
wire  myb ;
wire  mza ;
wire  mzb ;
wire  mzm ;
wire  naa ;
wire  NAA ;
wire  nam ;
wire  NAM ;
wire  nba ;
wire  NBA ;
wire  nbm ;
wire  NBM ;
wire  nda ;
wire  NDA ;
wire  ndm ;
wire  NDM ;
wire  nea ;
wire  NEA ;
wire  nem ;
wire  NEM ;
wire  oaa ;
wire  OAM ;
wire  oba ;
wire  OBM ;
wire  oca ;
wire  OCM ;
wire  oda ;
wire  oea ;
wire  oeb ;
wire  ofa ;
wire  ofb ;
wire  oga ;
wire  ogb ;
wire  oha ;
wire  ohb ;
wire  oia ;
wire  oib ;
wire  oja ;
wire  ojb ;
wire  oka ;
wire  okb ;
wire  ola ;
wire  olb ;
wire  oma ;
wire  omb ;
wire  ona ;
wire  onb ;
wire  ooa ;
wire  oob ;
wire  opa ;
wire  opb ;
wire  oqa ;
wire  oqb ;
wire  ora ;
wire  orb ;
wire  osa ;
wire  osb ;
wire  ota ;
wire  otb ;
wire  oua ;
wire  oub ;
wire  ova ;
wire  ovb ;
wire  owa ;
wire  owb ;
wire  oxa ;
wire  oxb ;
wire  oya ;
wire  oyb ;
wire  oza ;
wire  ozb ;
wire  ozm ;
wire  ozn ;
wire  QAA ;
wire  QAB ;
wire  QAC ;
wire  QAD ;
wire  QAE ;
wire  QAF ;
wire  QAG ;
wire  QAH ;
wire  QAI ;
wire  QAJ ;
wire  QAK ;
wire  QAL ;
wire  QAM ;
wire  qan ;
wire  qao ;
wire  qap ;
wire  qaq ;
wire  qar ;
wire  qas ;
wire  qat ;
wire  qau ;
wire  qav ;
wire  qaw ;
wire  qax ;
wire  qay ;
wire  qaz ;
wire  qba ;
wire  qbb ;
wire  qbc ;
wire  qbd ;
wire  qbe ;
wire  qia ;
wire  qib ;
wire  qic ;
wire  qid ;
wire  qie ;
wire  qra ;
wire  qta ;
wire  tra ;
wire  trb ;
wire  trc ;
wire  trd ;
wire  tre ;
wire  trf ;
wire  trg ;
wire  trh ;
wire  tta ;
wire  ttb ;
wire  ZZI ;
wire  ZZO ;
assign ZZI = 1'b1;
assign ZZO = 1'b0;
assign EAA =  CAZ & DAA  ; 
assign eaa = ~EAA;  //complement 
assign EAB =  CAY & DAB  ; 
assign eab = ~EAB;  //complement 
assign EAC =  CAX & DAC  ; 
assign eac = ~EAC;  //complement 
assign EDY =  CAE & DEY  ; 
assign edy = ~EDY;  //complement 
assign EDZ =  CAD & DEZ  ; 
assign edz = ~EDZ;  //complement 
assign EEE =  CAZ & DAE  ; 
assign eee = ~EEE;  //complement 
assign EEF =  CAY & DAF  ; 
assign eef = ~EEF;  //complement 
assign EEG =  CAX & DAG  ; 
assign eeg = ~EEG;  //complement 
assign EII =  CAZ & DAI  ; 
assign eii = ~EII;  //complement 
assign EIJ =  CAY & DAJ  ; 
assign eij = ~EIJ;  //complement 
assign EIK =  CAX & DAK  ; 
assign eik = ~EIK;  //complement 
assign faa = ~FAA;  //complement 
assign FAM = ~fam;  //complement 
assign fda = ~FDA;  //complement 
assign FDM = ~fdm;  //complement 
assign fea = ~FEA;  //complement 
assign FEM = ~fem;  //complement 
assign fia = ~FIA;  //complement 
assign FIM = ~fim;  //complement 
assign EBE =  CAW & DAE  ; 
assign ebe = ~EBE;  //complement 
assign EBF =  CAV & DAF  ; 
assign ebf = ~EBF;  //complement 
assign EBG =  CAU & DAG  ; 
assign ebg = ~EBG;  //complement 
assign EEQ =  CAN & DEQ  ; 
assign eeq = ~EEQ;  //complement 
assign EER =  CAM & DER  ; 
assign eer = ~EER;  //complement 
assign EES =  CAL & DES  ; 
assign ees = ~EES;  //complement 
assign EFI =  CAW & DAI  ; 
assign efi = ~EFI;  //complement 
assign EFJ =  CAV & DAJ  ; 
assign efj = ~EFJ;  //complement 
assign EFK =  CAU & DAK  ; 
assign efk = ~EFK;  //complement 
assign EGY =  CAH & DEY  ; 
assign egy = ~EGY;  //complement 
assign EGZ =  CAG & DEZ  ; 
assign egz = ~EGZ;  //complement 
assign fba = ~FBA;  //complement 
assign FBM = ~fbm;  //complement 
assign fca = ~FCA;  //complement 
assign FCM = ~fcm;  //complement 
assign ffa = ~FFA;  //complement 
assign FFM = ~ffm;  //complement 
assign fga = ~FGA;  //complement 
assign FGM = ~fgm;  //complement 
assign EBQ =  CAK & DEQ  ; 
assign ebq = ~EBQ;  //complement 
assign EBR =  CAJ & DER  ; 
assign ebr = ~EBR;  //complement 
assign EBS =  CAI & DES  ; 
assign ebs = ~EBS;  //complement 
assign ECI =  CAT & DAI  ; 
assign eci = ~ECI;  //complement 
assign ECJ =  CAS & DAJ  ; 
assign ecj = ~ECJ;  //complement 
assign ECK =  CAR & DAK  ; 
assign eck = ~ECK;  //complement 
assign EFV =  CAJ & DEV  ; 
assign efv = ~EFV;  //complement 
assign EFW =  CAI & DEW  ; 
assign efw = ~EFW;  //complement 
assign EFU =  CAK & DEU  ; 
assign efu = ~EFU;  //complement 
assign EGM =  CAT & DAM  ; 
assign egm = ~EGM;  //complement 
assign EGN =  CAS & DAN  ; 
assign egn = ~EGN;  //complement 
assign EGO =  CAR & DAO  ; 
assign ego = ~EGO;  //complement 
assign fbb = ~FBB;  //complement 
assign FBN = ~fbn;  //complement 
assign fcb = ~FCB;  //complement 
assign FCN = ~fcn;  //complement 
assign ffb = ~FFB;  //complement 
assign FFN = ~ffn;  //complement 
assign fgb = ~FGB;  //complement 
assign FGN = ~fgn;  //complement 
assign EAM =  CAN & DEM  ; 
assign eam = ~EAM;  //complement 
assign EAN =  CAM & DEN  ; 
assign ean = ~EAN;  //complement 
assign EAO =  CAL & DEO  ; 
assign eao = ~EAO;  //complement 
assign EDM =  CAQ & DEM  ; 
assign edm = ~EDM;  //complement 
assign EDN =  CAP & DEN  ; 
assign edn = ~EDN;  //complement 
assign EDO =  CAO & DEO  ; 
assign edo = ~EDO;  //complement 
assign ECU =  CAH & DEU  ; 
assign ecu = ~ECU;  //complement 
assign ECV =  CAG & DEV  ; 
assign ecv = ~ECV;  //complement 
assign ECW =  CAF & DEW  ; 
assign ecw = ~ECW;  //complement 
assign EHQ =  CAQ & DEQ  ; 
assign ehq = ~EHQ;  //complement 
assign EHR =  CAP & DER  ; 
assign ehr = ~EHR;  //complement 
assign EHS =  CAO & DES  ; 
assign ehs = ~EHS;  //complement 
assign fab = ~FAB;  //complement 
assign FAN = ~fan;  //complement 
assign fdb = ~FDB;  //complement 
assign FDN = ~fdn;  //complement 
assign feb = ~FEB;  //complement 
assign FEN = ~fen;  //complement 
assign fha = ~FHA;  //complement 
assign FHM = ~fhm;  //complement 
assign EMM =  CAZ & DAM  ; 
assign emm = ~EMM;  //complement 
assign EMN =  CAY & DAN  ; 
assign emn = ~EMN;  //complement 
assign EMO =  CAX & DAO  ; 
assign emo = ~EMO;  //complement 
assign EQQ =  CAZ & DAQ  ; 
assign eqq = ~EQQ;  //complement 
assign EQR =  CAY & DAR  ; 
assign eqr = ~EQR;  //complement 
assign EQS =  CAX & DAS  ; 
assign eqs = ~EQS;  //complement 
assign EUU =  CAZ & DAU  ; 
assign euu = ~EUU;  //complement 
assign EUV =  CAY & DAV  ; 
assign euv = ~EUV;  //complement 
assign EUW =  CAX & DAW  ; 
assign euw = ~EUW;  //complement 
assign fma = ~FMA;  //complement 
assign FMM = ~fmm;  //complement 
assign fqa = ~FQA;  //complement 
assign FQM = ~fqm;  //complement 
assign fua = ~FUA;  //complement 
assign FUM = ~fum;  //complement 
assign EJM =  CAW & DAM  ; 
assign ejm = ~EJM;  //complement 
assign EJN =  CAV & DAN  ; 
assign ejn = ~EJN;  //complement 
assign EJO =  CAU & DAO  ; 
assign ejo = ~EJO;  //complement 
assign ELU =  CAQ & DAU  ; 
assign elu = ~ELU;  //complement 
assign ELV =  CAP & DAV  ; 
assign elv = ~ELV;  //complement 
assign ELW =  CAO & DAW  ; 
assign elw = ~ELW;  //complement 
assign ENQ =  CAW & DAQ  ; 
assign enq = ~ENQ;  //complement 
assign ENR =  CAV & DAR  ; 
assign enr = ~ENR;  //complement 
assign ENS =  CAU & DAS  ; 
assign ens = ~ENS;  //complement 
assign ERU =  CAW & DAU  ; 
assign eru = ~ERU;  //complement 
assign ERV =  CAV & DAV  ; 
assign erv = ~ERV;  //complement 
assign ERW =  CAU & DAW  ; 
assign erw = ~ERW;  //complement 
assign fja = ~FJA;  //complement 
assign FJM = ~fjm;  //complement 
assign fna = ~FNA;  //complement 
assign FNM = ~fnm;  //complement 
assign fra = ~FRA;  //complement 
assign FRM = ~frm;  //complement 
assign EJY =  CAK & DEY  ; 
assign ejy = ~EJY;  //complement 
assign EJZ =  CAJ & DEZ  ; 
assign ejz = ~EJZ;  //complement 
assign EKQ =  CAT & DAQ  ; 
assign ekq = ~EKQ;  //complement 
assign EKR =  CAS & DAR  ; 
assign ekr = ~EKR;  //complement 
assign EKS =  CAR & DAS  ; 
assign eks = ~EKS;  //complement 
assign EOU =  CAT & DAU  ; 
assign eou = ~EOU;  //complement 
assign EOV =  CAS & DAV  ; 
assign eov = ~EOV;  //complement 
assign EOW =  CAR & DAW  ; 
assign eow = ~EOW;  //complement 
assign fjb = ~FJB;  //complement 
assign FJN = ~fjn;  //complement 
assign fka = ~FKA;  //complement 
assign FKM = ~fkm;  //complement 
assign foa = ~FOA;  //complement 
assign FOM = ~fom;  //complement 
assign EIU =  CAN & DEU  ; 
assign eiu = ~EIU;  //complement 
assign EIV =  CAM & DEV  ; 
assign eiv = ~EIV;  //complement 
assign EIW =  CAL & DEW  ; 
assign eiw = ~EIW;  //complement 
assign EMY =  CAN & DAY  ; 
assign emy = ~EMY;  //complement 
assign EMZ =  CAM & DAZ  ; 
assign emz = ~EMZ;  //complement 
assign fib = ~FIB;  //complement 
assign FIN = ~fin;  //complement 
assign fla = ~FLA;  //complement 
assign FLM = ~flm;  //complement 
assign fmb = ~FMB;  //complement 
assign FMN = ~fmn;  //complement 
assign EYY =  CAZ & DAY  ; 
assign eyy = ~EYY;  //complement 
assign EYZ =  CAY & DAZ  ; 
assign eyz = ~EYZ;  //complement 
assign daa = ~DAA;  //complement 
assign dab = ~DAB;  //complement 
assign dbb = ~DBB;  //complement 
assign fya = ~FYA;  //complement 
assign FYM = ~fym;  //complement 
assign EVY =  CAW & DAY  ; 
assign evy = ~EVY;  //complement 
assign EVZ =  CAV & DAZ  ; 
assign evz = ~EVZ;  //complement 
assign fva = ~FVA;  //complement 
assign FVM = ~fvm;  //complement 
assign qra = ~QRA;  //complement 
assign ESY =  CAT & DAY  ; 
assign esy = ~ESY;  //complement 
assign ESZ =  CAS & DAZ  ; 
assign esz = ~ESZ;  //complement 
assign fsa = ~FSA;  //complement 
assign FSM = ~fsm;  //complement 
assign tra = ~TRA;  //complement 
assign EPY =  CAQ & DAY  ; 
assign epy = ~EPY;  //complement 
assign EPZ =  CAP & DAZ  ; 
assign epz = ~EPZ;  //complement 
assign fpa = ~FPA;  //complement 
assign FPM = ~fpm;  //complement 
assign fac = ~FAC;  //complement 
assign FAO = ~fao;  //complement 
assign fbc = ~FBC;  //complement 
assign FBO = ~fbo;  //complement 
assign ffc = ~FFC;  //complement 
assign FFO = ~ffo;  //complement 
assign EAV =  CBE & DFV  ; 
assign eav = ~EAV;  //complement 
assign EAW =  CBD & DFW  ; 
assign eaw = ~EAW;  //complement 
assign EAX =  CBC & DFX  ; 
assign eax = ~EAX;  //complement 
assign EBB =  CBZ & DBB  ; 
assign ebb = ~EBB;  //complement 
assign EBC =  CBY & DBC  ; 
assign ebc = ~EBC;  //complement 
assign EBD =  CBX & DBD  ; 
assign ebd = ~EBD;  //complement 
assign EEZ =  CBE & DFZ  ; 
assign eez = ~EEZ;  //complement 
assign EFF =  CBZ & DBF  ; 
assign eff = ~EFF;  //complement 
assign EFG =  CBY & DBG  ; 
assign efg = ~EFG;  //complement 
assign EFH =  CBX & DBH  ; 
assign efh = ~EFH;  //complement 
assign fcc = ~FCC;  //complement 
assign FCO = ~fco;  //complement 
assign fdc = ~FDC;  //complement 
assign FDO = ~fdo;  //complement 
assign fgc = ~FGC;  //complement 
assign FGO = ~fgo;  //complement 
assign feh = ~FEH;  //complement 
assign fec = ~FEC;  //complement 
assign FEO = ~feo;  //complement 
assign ECF =  CBW & DBF  ; 
assign ecf = ~ECF;  //complement 
assign ECG =  CBV & DBG  ; 
assign ecg = ~ECG;  //complement 
assign ECH =  CBU & DBH  ; 
assign ech = ~ECH;  //complement 
assign EDV =  CBH & DFV  ; 
assign edv = ~EDV;  //complement 
assign EDW =  CBG & DFW  ; 
assign edw = ~EDW;  //complement 
assign EDX =  CBF & DFX  ; 
assign edx = ~EDX;  //complement 
assign EGJ =  CBW & DFJ  ; 
assign egj = ~EGJ;  //complement 
assign EGK =  CBV & DBK  ; 
assign egk = ~EGK;  //complement 
assign EGL =  CBU & DBL  ; 
assign egl = ~EGL;  //complement 
assign EHZ =  CBH & DFZ  ; 
assign ehz = ~EHZ;  //complement 
assign fcd = ~FCD;  //complement 
assign FCP = ~fcp;  //complement 
assign fdd = ~FDD;  //complement 
assign FDP = ~fdp;  //complement 
assign fgd = ~FGD;  //complement 
assign FGP = ~fgp;  //complement 
assign fhb = ~FHB;  //complement 
assign FHN = ~fhn;  //complement 
assign fhg = ~FHG;  //complement 
assign ECR =  CBK & DFR  ; 
assign ecr = ~ECR;  //complement 
assign ECS =  CBJ & DFS  ; 
assign ecs = ~ECS;  //complement 
assign ECT =  CBI & DFT  ; 
assign ect = ~ECT;  //complement 
assign EDJ =  CBT & DBJ  ; 
assign edj = ~EDJ;  //complement 
assign EDK =  CBS & DFK  ; 
assign edk = ~EDK;  //complement 
assign EDL =  CBR & DFL  ; 
assign edl = ~EDL;  //complement 
assign EGV =  CBK & DFV  ; 
assign egv = ~EGV;  //complement 
assign EGW =  CBJ & DFW  ; 
assign egw = ~EGW;  //complement 
assign EGX =  CBI & DFX  ; 
assign egx = ~EGX;  //complement 
assign fad = ~FAD;  //complement 
assign FAP = ~fap;  //complement 
assign fbd = ~FBD;  //complement 
assign FBP = ~fbp;  //complement 
assign EHN =  CBT & DFN  ; 
assign ehn = ~EHN;  //complement 
assign EHO =  CBS & DFO  ; 
assign eho = ~EHO;  //complement 
assign EHP =  CBR & DFP  ; 
assign ehp = ~EHP;  //complement 
assign ffd = ~FFD;  //complement 
assign FFP = ~ffp;  //complement 
assign EAJ =  CBQ & DBJ  ; 
assign eaj = ~EAJ;  //complement 
assign EAK =  CBP & DFK  ; 
assign eak = ~EAK;  //complement 
assign EAL =  CBO & DFL  ; 
assign eal = ~EAL;  //complement 
assign EBN =  CBN & DFN  ; 
assign ebn = ~EBN;  //complement 
assign EBO =  CBM & DFO  ; 
assign ebo = ~EBO;  //complement 
assign EBP =  CBL & DFP  ; 
assign ebp = ~EBP;  //complement 
assign EEN =  CBQ & DFN  ; 
assign een = ~EEN;  //complement 
assign EEO =  CBP & DFO  ; 
assign eeo = ~EEO;  //complement 
assign EEP =  CBO & DFP  ; 
assign eep = ~EEP;  //complement 
assign EFS =  CBM & DFS  ; 
assign efs = ~EFS;  //complement 
assign EFT =  CBL & DFT  ; 
assign eft = ~EFT;  //complement 
assign EFR =  CBN & DFR  ; 
assign efr = ~EFR;  //complement 
assign fjc = ~FJC;  //complement 
assign FJO = ~fjo;  //complement 
assign fnb = ~FNB;  //complement 
assign FNN = ~fnn;  //complement 
assign frb = ~FRB;  //complement 
assign FRN = ~frn;  //complement 
assign fwc = ~FWC;  //complement 
assign EJJ =  CBZ & DFJ  ; 
assign ejj = ~EJJ;  //complement 
assign EJK =  CBY & DBK  ; 
assign ejk = ~EJK;  //complement 
assign EJL =  CBX & DBL  ; 
assign ejl = ~EJL;  //complement 
assign ENN =  CBZ & DBN  ; 
assign enn = ~ENN;  //complement 
assign ENO =  CBY & DBO  ; 
assign eno = ~ENO;  //complement 
assign ENP =  CBX & DBP  ; 
assign enp = ~ENP;  //complement 
assign ERR =  CBZ & DBR  ; 
assign err = ~ERR;  //complement 
assign ERS =  CBY & DBS  ; 
assign ers = ~ERS;  //complement 
assign ERT =  CBX & DBT  ; 
assign ert = ~ERT;  //complement 
assign fkb = ~FKB;  //complement 
assign FKN = ~fkn;  //complement 
assign fkf = ~FKF;  //complement 
assign fjd = ~FJD;  //complement 
assign FJP = ~fjp;  //complement 
assign fob = ~FOB;  //complement 
assign FON = ~fon;  //complement 
assign fsb = ~FSB;  //complement 
assign FSN = ~fsn;  //complement 
assign ftd = ~FTD;  //complement 
assign EKN =  CBW & DBN  ; 
assign ekn = ~EKN;  //complement 
assign EKO =  CBV & DBO  ; 
assign eko = ~EKO;  //complement 
assign EKP =  CBU & DBP  ; 
assign ekp = ~EKP;  //complement 
assign EOR =  CBW & DBR  ; 
assign eor = ~EOR;  //complement 
assign EOS =  CBV & DBS  ; 
assign eos = ~EOS;  //complement 
assign EOT =  CBU & DBT  ; 
assign eot = ~EOT;  //complement 
assign ESV =  CBW & DBV  ; 
assign esv = ~ESV;  //complement 
assign ESW =  CBV & DBW  ; 
assign esw = ~ESW;  //complement 
assign ESX =  CBU & DBX  ; 
assign esx = ~ESX;  //complement 
assign flb = ~FLB;  //complement 
assign FLN = ~fln;  //complement 
assign fpb = ~FPB;  //complement 
assign FPN = ~fpn;  //complement 
assign fqe = ~FQE;  //complement 
assign EKZ =  CBK & DFZ  ; 
assign ekz = ~EKZ;  //complement 
assign ELR =  CBT & DBR  ; 
assign elr = ~ELR;  //complement 
assign ELS =  CBS & DBS  ; 
assign els = ~ELS;  //complement 
assign ELT =  CBR & DBT  ; 
assign elt = ~ELT;  //complement 
assign EPV =  CBT & DBV  ; 
assign epv = ~EPV;  //complement 
assign EPW =  CBS & DBW  ; 
assign epw = ~EPW;  //complement 
assign EPX =  CBR & DBX  ; 
assign epx = ~EPX;  //complement 
assign fic = ~FIC;  //complement 
assign FIO = ~fio;  //complement 
assign EIR =  CBQ & DFR  ; 
assign eir = ~EIR;  //complement 
assign EIS =  CBP & DFS  ; 
assign eis = ~EIS;  //complement 
assign EIT =  CBO & DFT  ; 
assign eit = ~EIT;  //complement 
assign fmc = ~FMC;  //complement 
assign FMO = ~fmo;  //complement 
assign fnf = ~FNF;  //complement 
assign EJV =  CBN & DBV  ; 
assign ejv = ~EJV;  //complement 
assign EJX =  CBL & DBX  ; 
assign ejx = ~EJX;  //complement 
assign EJW =  CBM & DBW  ; 
assign ejw = ~EJW;  //complement 
assign EMV =  CBQ & DBV  ; 
assign emv = ~EMV;  //complement 
assign EMW =  CBP & DBW  ; 
assign emw = ~EMW;  //complement 
assign EMX =  CBO & DBX  ; 
assign emx = ~EMX;  //complement 
assign fvb = ~FVB;  //complement 
assign FVN = ~fvn;  //complement 
assign daf = ~DAF;  //complement 
assign dbf = ~DBF;  //complement 
assign ddf = ~DDF;  //complement 
assign EVV =  CBZ & DBV  ; 
assign evv = ~EVV;  //complement 
assign EVW =  CBY & DBW  ; 
assign evw = ~EVW;  //complement 
assign EVX =  CBX & DBX  ; 
assign evx = ~EVX;  //complement 
assign daj = ~DAJ;  //complement 
assign dbj = ~DBJ;  //complement 
assign ddj = ~DDJ;  //complement 
assign dfj = ~DFJ;  //complement 
assign dag = ~DAG;  //complement 
assign dbg = ~DBG;  //complement 
assign dcg = ~DCG;  //complement 
assign ddr = ~DDR;  //complement 
assign ddv = ~DDV;  //complement 
assign DGK = ~dgk;  //complement 
assign dak = ~DAK;  //complement 
assign dbk = ~DBK;  //complement 
assign dck = ~DCK;  //complement 
assign dfk = ~DFK;  //complement 
assign CDF = ~cdf;  //complement 
assign CDG = ~cdg;  //complement 
assign EWZ =  CBW & DBZ  ; 
assign ewz = ~EWZ;  //complement 
assign dao = ~DAO;  //complement 
assign dbo = ~DBO;  //complement 
assign dco = ~DCO;  //complement 
assign deo = ~DEO;  //complement 
assign cag = ~CAG;  //complement 
assign cbg = ~CBG;  //complement 
assign ccg = ~CCG;  //complement 
assign caf = ~CAF;  //complement 
assign cbf = ~CBF;  //complement 
assign ccf = ~CCF;  //complement 
assign ftc = ~FTC;  //complement 
assign fuc = ~FUC;  //complement 
assign fwb = ~FWB;  //complement 
assign DFN = ~dfn;  //complement 
assign DFO = ~dfo;  //complement 
assign DGO = ~dgo;  //complement 
assign DHN = ~dhn;  //complement 
assign CDI = ~cdi;  //complement 
assign cai = ~CAI;  //complement 
assign cbi = ~CBI;  //complement 
assign cci = ~CCI;  //complement 
assign ETZ =  CBT & DBZ  ; 
assign etz = ~ETZ;  //complement 
assign DFV = ~dfv;  //complement 
assign DFW = ~dfw;  //complement 
assign DGW = ~dgw;  //complement 
assign DHV = ~dhv;  //complement 
assign dan = ~DAN;  //complement 
assign dbn = ~DBN;  //complement 
assign ddn = ~DDN;  //complement 
assign den = ~DEN;  //complement 
assign trb = ~TRB;  //complement 
assign fqd = ~FQD;  //complement 
assign daw = ~DAW;  //complement 
assign dbw = ~DBW;  //complement 
assign dcw = ~DCW;  //complement 
assign dew = ~DEW;  //complement 
assign dav = ~DAV;  //complement 
assign dbv = ~DBV;  //complement 
assign dev = ~DEV;  //complement 
assign EQZ =  CBQ & DBZ  ; 
assign eqz = ~EQZ;  //complement 
assign DFR = ~dfr;  //complement 
assign DFS = ~dfs;  //complement 
assign DGS = ~dgs;  //complement 
assign DHR = ~dhr;  //complement 
assign dar = ~DAR;  //complement 
assign dbr = ~DBR;  //complement 
assign der = ~DER;  //complement 
assign das = ~DAS;  //complement 
assign dbs = ~DBS;  //complement 
assign dcs = ~DCS;  //complement 
assign des = ~DES;  //complement 
assign haa = ~HAA;  //complement 
assign HAM = ~ham;  //complement 
assign GBA =  FBC & fao & fbi  |  fbc & FAO & fbi  |  fbc & fao & FBI  |  FBC & FAO & FBI  ; 
assign gba = ~GBA; //complement 
assign gbm =  FBC & fao & fbi  |  fbc & FAO & fbi  |  fbc & fao & FBI  |  fbc & fao & fbi  ; 
assign GBM = ~gbm;  //complement 
assign hea = ~HEA;  //complement 
assign HEM = ~hem;  //complement 
assign hgd = ~HGD;  //complement 
assign GFA =  FEM & ffc & fff  |  fem & FFC & fff  |  fem & ffc & FFF  |  FEM & FFC & FFF  ; 
assign gfa = ~GFA; //complement 
assign gfm =  FEM & ffc & fff  |  fem & FFC & fff  |  fem & ffc & FFF  |  fem & ffc & fff  ; 
assign GFM = ~gfm;  //complement 
assign GAA =  FAH & faa & fac  |  fah & FAA & fac  |  fah & faa & FAC  |  FAH & FAA & FAC  ; 
assign gaa = ~GAA; //complement 
assign gam =  FAH & faa & fac  |  fah & FAA & fac  |  fah & faa & FAC  |  fah & faa & fac  ; 
assign GAM = ~gam;  //complement 
assign hba = ~HBA;  //complement 
assign HBM = ~hbm;  //complement 
assign GEA =  FDS & fea & fdm  |  fds & FEA & fdm  |  fds & fea & FDM  |  FDS & FEA & FDM  ; 
assign gea = ~GEA; //complement 
assign gem =  FDS & fea & fdm  |  fds & FEA & fdm  |  fds & fea & FDM  |  fds & fea & fdm  ; 
assign GEM = ~gem;  //complement 
assign hha = ~HHA;  //complement 
assign HHM = ~hhm;  //complement 
assign had = ~HAD;  //complement 
assign HAP = ~hap;  //complement 
assign hed = ~HED;  //complement 
assign HEP = ~hep;  //complement 
assign GEB =  FEH & fdo & fef  |  feh & FDO & fef  |  feh & fdo & FEF  |  FEH & FDO & FEF  ; 
assign geb = ~GEB; //complement 
assign gen =  FEH & fdo & fef  |  feh & FDO & fef  |  feh & fdo & FEF  |  feh & fdo & fef  ; 
assign GEN = ~gen;  //complement 
assign hfa = ~HFA;  //complement 
assign HFM = ~hfm;  //complement 
assign hfd = ~HFD;  //complement 
assign GCC =  FCA & fbm & fbt  |  fca & FBM & fbt  |  fca & fbm & FBT  |  FCA & FBM & FBT  ; 
assign gcc = ~GCC; //complement 
assign gco =  FCA & fbm & fbt  |  fca & FBM & fbt  |  fca & fbm & FBT  |  fca & fbm & fbt  ; 
assign GCO = ~gco;  //complement 
assign GFB =  FFA & fep & fer  |  ffa & FEP & fer  |  ffa & fep & FER  |  FFA & FEP & FER  ; 
assign gfb = ~GFB; //complement 
assign gfn =  FFA & fep & fer  |  ffa & FEP & fer  |  ffa & fep & FER  |  ffa & fep & fer  ; 
assign GFN = ~gfn;  //complement 
assign GGB =  FGA & ffm & fgc  |  fga & FFM & fgc  |  fga & ffm & FGC  |  FGA & FFM & FGC  ; 
assign ggb = ~GGB; //complement 
assign ggn =  FGA & ffm & fgc  |  fga & FFM & fgc  |  fga & ffm & FGC  |  fga & ffm & fgc  ; 
assign GGN = ~ggn;  //complement 
assign hac = ~HAC;  //complement 
assign HAO = ~hao;  //complement 
assign hcb = ~HCB;  //complement 
assign HCN = ~hcn;  //complement 
assign hde = ~HDE;  //complement 
assign hec = ~HEC;  //complement 
assign HEO = ~heo;  //complement 
assign hga = ~HGA;  //complement 
assign HGM = ~hgm;  //complement 
assign GCD =  FBN & fcb & fch  |  fbn & FCB & fch  |  fbn & fcb & FCH  |  FBN & FCB & FCH  ; 
assign gcd = ~GCD; //complement 
assign gcp =  FBN & fcb & fch  |  fbn & FCB & fch  |  fbn & fcb & FCH  |  fbn & fcb & fch  ; 
assign GCP = ~gcp;  //complement 
assign GDD =  FDF & fcn & fcp  |  fdf & FCN & fcp  |  fdf & fcn & FCP  |  FDF & FCN & FCP  ; 
assign gdd = ~GDD; //complement 
assign gdp =  FDF & fcn & fcp  |  fdf & FCN & fcp  |  fdf & fcn & FCP  |  fdf & fcn & fcp  ; 
assign GDP = ~gdp;  //complement 
assign hdb = ~HDB;  //complement 
assign HDN = ~hdn;  //complement 
assign GGC =  FGB & ffn & ffs  |  fgb & FFN & ffs  |  fgb & ffn & FFS  |  FGB & FFN & FFS  ; 
assign ggc = ~GGC; //complement 
assign ggo =  FGB & ffn & ffs  |  fgb & FFN & ffs  |  fgb & ffn & FFS  |  fgb & ffn & ffs  ; 
assign GGO = ~ggo;  //complement 
assign GBF =  FBF & fbd & fap  |  fbf & FBD & fap  |  fbf & fbd & FAP  |  FBF & FBD & FAP  ; 
assign gbf = ~GBF; //complement 
assign gbr =  FBF & fbd & fap  |  fbf & FBD & fap  |  fbf & fbd & FAP  |  fbf & fbd & fap  ; 
assign GBR = ~gbr;  //complement 
assign GDB =  FDA & fdc & fco  |  fda & FDC & fco  |  fda & fdc & FCO  |  FDA & FDC & FCO  ; 
assign gdb = ~GDB; //complement 
assign gdn =  FDA & fdc & fco  |  fda & FDC & fco  |  fda & fdc & FCO  |  fda & fdc & fco  ; 
assign GDN = ~gdn;  //complement 
assign GFD =  FFB & ffd & feo  |  ffb & FFD & feo  |  ffb & ffd & FEO  |  FFB & FFD & FEO  ; 
assign gfd = ~GFD; //complement 
assign gfp =  FFB & ffd & feo  |  ffb & FFD & feo  |  ffb & ffd & FEO  |  ffb & ffd & feo  ; 
assign GFP = ~gfp;  //complement 
assign GAC =  FAG & fad & fab  |  fag & FAD & fab  |  fag & fad & FAB  |  FAG & FAD & FAB  ; 
assign gac = ~GAC; //complement 
assign gao =  FAG & fad & fab  |  fag & FAD & fab  |  fag & fad & FAB  |  fag & fad & fab  ; 
assign GAO = ~gao;  //complement 
assign hbc = ~HBC;  //complement 
assign HBO = ~hbo;  //complement 
assign GEE =  FEC & feb & fdn  |  fec & FEB & fdn  |  fec & feb & FDN  |  FEC & FEB & FDN  ; 
assign gee = ~GEE; //complement 
assign geq =  FEC & feb & fdn  |  fec & FEB & fdn  |  fec & feb & FDN  |  fec & feb & fdn  ; 
assign GEQ = ~geq;  //complement 
assign hfc = ~HFC;  //complement 
assign HFO = ~hfo;  //complement 
assign hka = ~HKA;  //complement 
assign HKM = ~hkm;  //complement 
assign GOA =  FOC & fnn & fob  |  foc & FNN & fob  |  foc & fnn & FOB  |  FOC & FNN & FOB  ; 
assign goa = ~GOA; //complement 
assign gom =  FOC & fnn & fob  |  foc & FNN & fob  |  foc & fnn & FOB  |  foc & fnn & fob  ; 
assign GOM = ~gom;  //complement 
assign fxb = ~FXB;  //complement 
assign GJA =  FIM & fjc & fiq  |  fim & FJC & fiq  |  fim & fjc & FIQ  |  FIM & FJC & FIQ  ; 
assign gja = ~GJA; //complement 
assign gjm =  FIM & fjc & fiq  |  fim & FJC & fiq  |  fim & fjc & FIQ  |  fim & fjc & fiq  ; 
assign GJM = ~gjm;  //complement 
assign GNA =  FNB & fmm & fmq  |  fnb & FMM & fmq  |  fnb & fmm & FMQ  |  FNB & FMM & FMQ  ; 
assign gna = ~GNA; //complement 
assign gnm =  FNB & fmm & fmq  |  fnb & FMM & fmq  |  fnb & fmm & FMQ  |  fnb & fmm & fmq  ; 
assign GNM = ~gnm;  //complement 
assign GRA =  FQO & fqm & frb  |  fqo & FQM & frb  |  fqo & fqm & FRB  |  FQO & FQM & FRB  ; 
assign gra = ~GRA; //complement 
assign grm =  FQO & fqm & frb  |  fqo & FQM & frb  |  fqo & fqm & FRB  |  fqo & fqm & frb  ; 
assign GRM = ~grm;  //complement 
assign hja = ~HJA;  //complement 
assign HJM = ~hjm;  //complement 
assign GJC =  FJD & fip & fjb  |  fjd & FIP & fjb  |  fjd & fip & FJB  |  FJD & FIP & FJB  ; 
assign gjc = ~GJC; //complement 
assign gjo =  FJD & fip & fjb  |  fjd & FIP & fjb  |  fjd & fip & FJB  |  fjd & fip & fjb  ; 
assign GJO = ~gjo;  //complement 
assign hoa = ~HOA;  //complement 
assign HOM = ~hom;  //complement 
assign hqb = ~HQB;  //complement 
assign hpa = ~HPA;  //complement 
assign HPM = ~hpm;  //complement 
assign GJB =  FJA & fir & fjf  |  fja & FIR & fjf  |  fja & fir & FJF  |  FJA & FIR & FJF  ; 
assign gjb = ~GJB; //complement 
assign gjn =  FJA & fir & fjf  |  fja & FIR & fjf  |  fja & fir & FJF  |  fja & fir & fjf  ; 
assign GJN = ~gjn;  //complement 
assign GKB =  FJM & fjn & fkb  |  fjm & FJN & fkb  |  fjm & fjn & FKB  |  FJM & FJN & FKB  ; 
assign gkb = ~GKB; //complement 
assign gkn =  FJM & fjn & fkb  |  fjm & FJN & fkb  |  fjm & fjn & FKB  |  fjm & fjn & fkb  ; 
assign GKN = ~gkn;  //complement 
assign GPA =  FON & fpb & fpc  |  fon & FPB & fpc  |  fon & fpb & FPC  |  FON & FPB & FPC  ; 
assign gpa = ~GPA; //complement 
assign gpm =  FON & fpb & fpc  |  fon & FPB & fpc  |  fon & fpb & FPC  |  fon & fpb & fpc  ; 
assign GPM = ~gpm;  //complement 
assign hra = ~HRA;  //complement 
assign HRM = ~hrm;  //complement 
assign GHC =  FGP & fhb & fhg  |  fgp & FHB & fhg  |  fgp & fhb & FHG  |  FGP & FHB & FHG  ; 
assign ghc = ~GHC; //complement 
assign gho =  FGP & fhb & fhg  |  fgp & FHB & fhg  |  fgp & fhb & FHG  |  fgp & fhb & fhg  ; 
assign GHO = ~gho;  //complement 
assign ELN =  CDX & DDN  ; 
assign eln = ~ELN;  //complement 
assign hlb = ~HLB;  //complement 
assign HLN = ~hln;  //complement 
assign GOB =  FNM & foa & fnp  |  fnm & FOA & fnp  |  fnm & foa & FNP  |  FNM & FOA & FNP  ; 
assign gob = ~GOB; //complement 
assign gon =  FNM & foa & fnp  |  fnm & FOA & fnp  |  fnm & foa & FNP  |  fnm & foa & fnp  ; 
assign GON = ~gon;  //complement 
assign hgb = ~HGB;  //complement 
assign HGN = ~hgn;  //complement 
assign hid = ~HID;  //complement 
assign hkc = ~HKC;  //complement 
assign HKO = ~hko;  //complement 
assign hnb = ~HNB;  //complement 
assign HNN = ~hnn;  //complement 
assign GID =  FIC & fib & fhm  |  fic & FIB & fhm  |  fic & fib & FHM  |  FIC & FIB & FHM  ; 
assign gid = ~GID; //complement 
assign gip =  FIC & fib & fhm  |  fic & FIB & fhm  |  fic & fib & FHM  |  fic & fib & fhm  ; 
assign GIP = ~gip;  //complement 
assign GNC =  FMO & fmn & fnf  |  fmo & FMN & fnf  |  fmo & fmn & FNF  |  FMO & FMN & FNF  ; 
assign gnc = ~GNC; //complement 
assign gno =  FMO & fmn & fnf  |  fmo & FMN & fnf  |  fmo & fmn & FNF  |  fmo & fmn & fnf  ; 
assign GNO = ~gno;  //complement 
assign GHE =  FHA & fgr & fhf  |  fha & FGR & fhf  |  fha & fgr & FHF  |  FHA & FGR & FHF  ; 
assign ghe = ~GHE; //complement 
assign ghq =  FHA & fgr & fhf  |  fha & FGR & fhf  |  fha & fgr & FHF  |  fha & fgr & fhf  ; 
assign GHQ = ~ghq;  //complement 
assign GSA =  FSC & frn & fsb  |  fsc & FRN & fsb  |  fsc & frn & FSB  |  FSC & FRN & FSB  ; 
assign gsa = ~GSA; //complement 
assign gsm =  FSC & frn & fsb  |  fsc & FRN & fsb  |  fsc & frn & FSB  |  fsc & frn & fsb  ; 
assign GSM = ~gsm;  //complement 
assign GKD =  FKF & fjq & fkd  |  fkf & FJQ & fkd  |  fkf & fjq & FKD  |  FKF & FJQ & FKD  ; 
assign gkd = ~GKD; //complement 
assign gkp =  FKF & fjq & fkd  |  fkf & FJQ & fkd  |  fkf & fjq & FKD  |  fkf & fjq & fkd  ; 
assign GKP = ~gkp;  //complement 
assign GMC =  FMC & fmb & flm  |  fmc & FMB & flm  |  fmc & fmb & FLM  |  FMC & FMB & FLM  ; 
assign gmc = ~GMC; //complement 
assign gmo =  FMC & fmb & flm  |  fmc & FMB & flm  |  fmc & fmb & FLM  |  fmc & fmb & flm  ; 
assign GMO = ~gmo;  //complement 
assign GWA =  FVN & fwc & fwa  |  fvn & FWC & fwa  |  fvn & fwc & FWA  |  FVN & FWC & FWA  ; 
assign gwa = ~GWA; //complement 
assign gwm =  FVN & fwc & fwa  |  fvn & FWC & fwa  |  fvn & fwc & FWA  |  fvn & fwc & fwa  ; 
assign GWM = ~gwm;  //complement 
assign hwa = ~HWA;  //complement 
assign HWM = ~hwm;  //complement 
assign qaw = ~QAW;  //complement 
assign dac = ~DAC;  //complement 
assign dbc = ~DBC;  //complement 
assign dcc = ~DCC;  //complement 
assign GVA =  FUN & fvb & fum  |  fun & FVB & fum  |  fun & fvb & FUM  |  FUN & FVB & FUM  ; 
assign gva = ~GVA; //complement 
assign gvm =  FUN & fvb & fum  |  fun & FVB & fum  |  fun & fvb & FUM  |  fun & fvb & fum  ; 
assign GVM = ~gvm;  //complement 
assign hva = ~HVA;  //complement 
assign HVM = ~hvm;  //complement 
assign qay = ~QAY;  //complement 
assign cad = ~CAD;  //complement 
assign cbd = ~CBD;  //complement 
assign ccd = ~CCD;  //complement 
assign hsa = ~HSA;  //complement 
assign HSM = ~hsm;  //complement 
assign htb = ~HTB;  //complement 
assign QAJ = ~qaj;  //complement 
assign QAM = ~qam;  //complement 
assign qbc = ~QBC;  //complement 
assign qbe = ~QBE;  //complement 
assign QAD = ~qad;  //complement 
assign QAG = ~qag;  //complement 
assign ozn = ~OZN;  //complement 
assign qbb = ~QBB;  //complement 
assign qbd = ~QBD;  //complement 
assign GSB =  FRM & fsa & fro  |  frm & FSA & fro  |  frm & fsa & FRO  |  FRM & FSA & FRO  ; 
assign gsb = ~GSB; //complement 
assign gsn =  FRM & fsa & fro  |  frm & FSA & fro  |  frm & fsa & FRO  |  frm & fsa & fro  ; 
assign GSN = ~gsn;  //complement 
assign hta = ~HTA;  //complement 
assign HTM = ~htm;  //complement 
assign qat = ~QAT;  //complement 
assign qav = ~QAV;  //complement 
assign CDD = ~cdd;  //complement 
assign GQB =  FPN & fqe & fpo  |  fpn & FQE & fpo  |  fpn & fqe & FPO  |  FPN & FQE & FPO  ; 
assign gqb = ~GQB; //complement 
assign gqn =  FPN & fqe & fpo  |  fpn & FQE & fpo  |  fpn & fqe & FPO  |  fpn & fqe & fpo  ; 
assign GQN = ~gqn;  //complement 
assign hpb = ~HPB;  //complement 
assign HPN = ~hpn;  //complement 
assign hwb = ~HWB;  //complement 
assign qba = ~QBA;  //complement 
assign hob = ~HOB;  //complement 
assign HON = ~hon;  //complement 
assign trf = ~TRF;  //complement 
assign qaq = ~QAQ;  //complement 
assign qas = ~QAS;  //complement 
assign tre = ~TRE;  //complement 
assign GPB =  FOP & fom & fpa  |  fop & FOM & fpa  |  fop & fom & FPA  |  FOP & FOM & FPA  ; 
assign gpb = ~GPB; //complement 
assign gpn =  FOP & fom & fpa  |  fop & FOM & fpa  |  fop & fom & FPA  |  fop & fom & fpa  ; 
assign GPN = ~gpn;  //complement 
assign hqa = ~HQA;  //complement 
assign HQM = ~hqm;  //complement 
assign caq = ~CAQ;  //complement 
assign cbq = ~CBQ;  //complement 
assign ccq = ~CCQ;  //complement 
assign cdq = ~CDQ;  //complement 
assign GQC =  FQD & fqb & fpm  |  fqd & FQB & fpm  |  fqd & fqb & FPM  |  FQD & FQB & FPM  ; 
assign gqc = ~GQC; //complement 
assign gqo =  FQD & fqb & fpm  |  fqd & FQB & fpm  |  fqd & fqb & FPM  |  fqd & fqb & fpm  ; 
assign GQO = ~gqo;  //complement 
assign qan = ~QAN;  //complement 
assign qap = ~QAP;  //complement 
assign cap = ~CAP;  //complement 
assign cbp = ~CBP;  //complement 
assign ccp = ~CCP;  //complement 
assign cdp = ~CDP;  //complement 
assign JEB =  HEC & hdn & hed  |  hec & HDN & hed  |  hec & hdn & HED  |  HEC & HDN & HED  ; 
assign jeb = ~JEB; //complement 
assign jen =  HEC & hdn & hed  |  hec & HDN & hed  |  hec & hdn & HED  |  hec & hdn & hed  ; 
assign JEN = ~jen;  //complement 
assign kfa = ~KFA;  //complement 
assign KFM = ~kfm;  //complement 
assign mab = ~MAB;  //complement 
assign LGA =  KFM & kga & kgb  |  kfm & KGA & kgb  |  kfm & kga & KGB  |  KFM & KGA & KGB  ; 
assign lga = ~LGA; //complement 
assign lgm =  KFM & kga & kgb  |  kfm & KGA & kgb  |  kfm & kga & KGB  |  kfm & kga & kgb  ; 
assign LGM = ~lgm;  //complement 
assign JBA =  HAM & hba & han  |  ham & HBA & han  |  ham & hba & HAN  |  HAM & HBA & HAN  ; 
assign jba = ~JBA; //complement 
assign jbm =  HAM & hba & han  |  ham & HBA & han  |  ham & hba & HAN  |  ham & hba & han  ; 
assign JBM = ~jbm;  //complement 
assign mga = ~MGA;  //complement 
assign MGM = ~mgm;  //complement 
assign kga = ~KGA;  //complement 
assign KGM = ~kgm;  //complement 
assign kib = ~KIB;  //complement 
assign JAA =  HAA & hac & hab  |  haa & HAC & hab  |  haa & hac & HAB  |  HAA & HAC & HAB  ; 
assign jaa = ~JAA; //complement 
assign jam =  HAA & hac & hab  |  haa & HAC & hab  |  haa & hac & HAB  |  haa & hac & hab  ; 
assign JAM = ~jam;  //complement 
assign keb = ~KEB;  //complement 
assign KEN = ~ken;  //complement 
assign mbc = ~MBC;  //complement 
assign LFA =  KFA & kem & ken  |  kfa & KEM & ken  |  kfa & kem & KEN  |  KFA & KEM & KEN  ; 
assign lfa = ~LFA; //complement 
assign lfm =  KFA & kem & ken  |  kfa & KEM & ken  |  kfa & kem & KEN  |  kfa & kem & ken  ; 
assign LFM = ~lfm;  //complement 
assign JFA =  HFA & hfd & hen  |  hfa & HFD & hen  |  hfa & hfd & HEN  |  HFA & HFD & HEN  ; 
assign jfa = ~JFA; //complement 
assign jfm =  HFA & hfd & hen  |  hfa & HFD & hen  |  hfa & hfd & HEN  |  hfa & hfd & hen  ; 
assign JFM = ~jfm;  //complement 
assign mba = ~MBA;  //complement 
assign MBM = ~mbm;  //complement 
assign mbb = ~MBB;  //complement 
assign LCA =  KCA & kbm & kbn  |  kca & KBM & kbn  |  kca & kbm & KBN  |  KCA & KBM & KBN  ; 
assign lca = ~LCA; //complement 
assign lcm =  KCA & kbm & kbn  |  kca & KBM & kbn  |  kca & kbm & KBN  |  kca & kbm & kbn  ; 
assign LCM = ~lcm;  //complement 
assign mfa = ~MFA;  //complement 
assign MFM = ~mfm;  //complement 
assign JHA =  HHA & hgm & hhb  |  hha & HGM & hhb  |  hha & hgm & HHB  |  HHA & HGM & HHB  ; 
assign jha = ~JHA; //complement 
assign jhm =  HHA & hgm & hhb  |  hha & HGM & hhb  |  hha & hgm & HHB  |  hha & hgm & hhb  ; 
assign JHM = ~jhm;  //complement 
assign LAA =  KAB & kad & kac  |  kab & KAD & kac  |  kab & kad & KAC  |  KAB & KAD & KAC  ; 
assign laa = ~LAA; //complement 
assign lam =  KAB & kad & kac  |  kab & KAD & kac  |  kab & kad & KAC  |  kab & kad & kac  ; 
assign LAM = ~lam;  //complement 
assign JDB =  HDE & hcn & hdb  |  hde & HCN & hdb  |  hde & hcn & HDB  |  HDE & HCN & HDB  ; 
assign jdb = ~JDB; //complement 
assign jdn =  HDE & hcn & hdb  |  hde & HCN & hdb  |  hde & hcn & HDB  |  hde & hcn & hdb  ; 
assign JDN = ~jdn;  //complement 
assign JFB =  HEO & hfb & hep  |  heo & HFB & hep  |  heo & hfb & HEP  |  HEO & HFB & HEP  ; 
assign jfb = ~JFB; //complement 
assign jfn =  HEO & hfb & hep  |  heo & HFB & hep  |  heo & hfb & HEP  |  heo & hfb & hep  ; 
assign JFN = ~jfn;  //complement 
assign kgb = ~KGB;  //complement 
assign KGN = ~kgn;  //complement 
assign khb = ~KHB;  //complement 
assign kab = ~KAB;  //complement 
assign KAN = ~kan;  //complement 
assign kad = ~KAD;  //complement 
assign LBA =  KAN & kbb & kbc  |  kan & KBB & kbc  |  kan & kbb & KBC  |  KAN & KBB & KBC  ; 
assign lba = ~LBA; //complement 
assign lbm =  KAN & kbb & kbc  |  kan & KBB & kbc  |  kan & kbb & KBC  |  kan & kbb & kbc  ; 
assign LBM = ~lbm;  //complement 
assign LHA =  KHB & kgn & kha  |  khb & KGN & kha  |  khb & kgn & KHA  |  KHB & KGN & KHA  ; 
assign lha = ~LHA; //complement 
assign lhm =  KHB & kgn & kha  |  khb & KGN & kha  |  khb & kgn & KHA  |  khb & kgn & kha  ; 
assign LHM = ~lhm;  //complement 
assign kbb = ~KBB;  //complement 
assign KBN = ~kbn;  //complement 
assign kbc = ~KBC;  //complement 
assign kba = ~KBA;  //complement 
assign KBM = ~kbm;  //complement 
assign JGA =  HGB & hfo & hgc  |  hgb & HFO & hgc  |  hgb & hfo & HGC  |  HGB & HFO & HGC  ; 
assign jga = ~JGA; //complement 
assign jgm =  HGB & hfo & hgc  |  hgb & HFO & hgc  |  hgb & hfo & HGC  |  hgb & hfo & hgc  ; 
assign JGM = ~jgm;  //complement 
assign mca = ~MCA;  //complement 
assign MCM = ~mcm;  //complement 
assign mdb = ~MDB;  //complement 
assign kfb = ~KFB;  //complement 
assign KFN = ~kfn;  //complement 
assign NDA =  MDA & mcm & mdb  |  mda & MCM & mdb  |  mda & mcm & MDB  |  MDA & MCM & MDB  ; 
assign nda = ~NDA; //complement 
assign ndm =  MDA & mcm & mdb  |  mda & MCM & mdb  |  mda & mcm & MDB  |  mda & mcm & mdb  ; 
assign NDM = ~ndm;  //complement 
assign mha = ~MHA;  //complement 
assign MHM = ~mhm;  //complement 
assign JLA =  HKM & hlb & hla  |  hkm & HLB & hla  |  hkm & hlb & HLA  |  HKM & HLB & HLA  ; 
assign jla = ~JLA; //complement 
assign jlm =  HKM & hlb & hla  |  hkm & HLB & hla  |  hkm & hlb & HLA  |  hkm & hlb & hla  ; 
assign JLM = ~jlm;  //complement 
assign kic = ~KIC;  //complement 
assign JJA =  HJA & him & hin  |  hja & HIM & hin  |  hja & him & HIN  |  HJA & HIM & HIN  ; 
assign jja = ~JJA; //complement 
assign jjm =  HJA & him & hin  |  hja & HIM & hin  |  hja & him & HIN  |  hja & him & hin  ; 
assign JJM = ~jjm;  //complement 
assign kka = ~KKA;  //complement 
assign KKM = ~kkm;  //complement 
assign JQA =  HPM & hqb & hqc  |  hpm & HQB & hqc  |  hpm & hqb & HQC  |  HPM & HQB & HQC  ; 
assign jqa = ~JQA; //complement 
assign jqm =  HPM & hqb & hqc  |  hpm & HQB & hqc  |  hpm & hqb & HQC  |  hpm & hqb & hqc  ; 
assign JQM = ~jqm;  //complement 
assign LIA =  KIC & kib & kia  |  kic & KIB & kia  |  kic & kib & KIA  |  KIC & KIB & KIA  ; 
assign lia = ~LIA; //complement 
assign lim =  KIC & kib & kia  |  kic & KIB & kia  |  kic & kib & KIA  |  kic & kib & kia  ; 
assign LIM = ~lim;  //complement 
assign mka = ~MKA;  //complement 
assign MKM = ~mkm;  //complement 
assign mla = ~MLA;  //complement 
assign MLM = ~mlm;  //complement 
assign koa = ~KOA;  //complement 
assign KOM = ~kom;  //complement 
assign kpb = ~KPB;  //complement 
assign kpa = ~KPA;  //complement 
assign KPM = ~kpm;  //complement 
assign kqb = ~KQB;  //complement 
assign mia = ~MIA;  //complement 
assign MIM = ~mim;  //complement 
assign JOA =  HNN & hob & hnm  |  hnn & HOB & hnm  |  hnn & hob & HNM  |  HNN & HOB & HNM  ; 
assign joa = ~JOA; //complement 
assign jom =  HNN & hob & hnm  |  hnn & HOB & hnm  |  hnn & hob & HNM  |  hnn & hob & hnm  ; 
assign JOM = ~jom;  //complement 
assign oda = ~ODA;  //complement 
assign oea = ~OEA;  //complement 
assign cax = ~CAX;  //complement 
assign cbx = ~CBX;  //complement 
assign ccx = ~CCX;  //complement 
assign cdx = ~CDX;  //complement 
assign JXA =  HXB & hwm & hxa  |  hxb & HWM & hxa  |  hxb & hwm & HXA  |  HXB & HWM & HXA  ; 
assign jxa = ~JXA; //complement 
assign jxm =  HXB & hwm & hxa  |  hxb & HWM & hxa  |  hxb & hwm & HXA  |  hxb & hwm & hxa  ; 
assign JXM = ~jxm;  //complement 
assign mwb = ~MWB;  //complement 
assign mxa = ~MXA;  //complement 
assign mxb = ~MXB;  //complement 
assign myb = ~MYB;  //complement 
assign owb = ~OWB;  //complement 
assign oxa = ~OXA;  //complement 
assign oxb = ~OXB;  //complement 
assign oyb = ~OYB;  //complement 
assign JWA =  HWA & hvm & hwb  |  hwa & HVM & hwb  |  hwa & hvm & HWB  |  HWA & HVM & HWB  ; 
assign jwa = ~JWA; //complement 
assign jwm =  HWA & hvm & hwb  |  hwa & HVM & hwb  |  hwa & hvm & HWB  |  hwa & hvm & hwb  ; 
assign JWM = ~jwm;  //complement 
assign kwa = ~KWA;  //complement 
assign kxa = ~KXA;  //complement 
assign kxb = ~KXB;  //complement 
assign kyb = ~KYB;  //complement 
assign ogb = ~OGB;  //complement 
assign oha = ~OHA;  //complement 
assign ohb = ~OHB;  //complement 
assign oia = ~OIA;  //complement 
assign JTA =  HSM & htb & hta  |  hsm & HTB & hta  |  hsm & htb & HTA  |  HSM & HTB & HTA  ; 
assign jta = ~JTA; //complement 
assign jtm =  HSM & htb & hta  |  hsm & HTB & hta  |  hsm & htb & HTA  |  hsm & htb & hta  ; 
assign JTM = ~jtm;  //complement 
assign cau = ~CAU;  //complement 
assign cbu = ~CBU;  //complement 
assign cdu = ~CDU;  //complement 
assign cav = ~CAV;  //complement 
assign cbv = ~CBV;  //complement 
assign ccv = ~CCV;  //complement 
assign cdv = ~CDV;  //complement 
assign krb = ~KRB;  //complement 
assign LPA =  KOM & kpb & kpa  |  kom & KPB & kpa  |  kom & kpb & KPA  |  KOM & KPB & KPA  ; 
assign lpa = ~LPA; //complement 
assign lpm =  KOM & kpb & kpa  |  kom & KPB & kpa  |  kom & kpb & KPA  |  kom & kpb & kpa  ; 
assign LPM = ~lpm;  //complement 
assign mpb = ~MPB;  //complement 
assign mqa = ~MQA;  //complement 
assign mqb = ~MQB;  //complement 
assign mra = ~MRA;  //complement 
assign ofb = ~OFB;  //complement 
assign oga = ~OGA;  //complement 
assign ola = ~OLA;  //complement 
assign olb = ~OLB;  //complement 
assign JRA =  HRA & hqm & hrb  |  hra & HQM & hrb  |  hra & hqm & HRB  |  HRA & HQM & HRB  ; 
assign jra = ~JRA; //complement 
assign jrm =  HRA & hqm & hrb  |  hra & HQM & hrb  |  hra & hqm & HRB  |  hra & hqm & hrb  ; 
assign JRM = ~jrm;  //complement 
assign LQA =  KQA & kpm & kqb  |  kqa & KPM & kqb  |  kqa & kpm & KQB  |  KQA & KPM & KQB  ; 
assign lqa = ~LQA; //complement 
assign lqm =  KQA & kpm & kqb  |  kqa & KPM & kqb  |  kqa & kpm & KQB  |  kqa & kpm & kqb  ; 
assign LQM = ~lqm;  //complement 
assign qta = ~QTA;  //complement 
assign tta = ~TTA;  //complement 
assign ttb = ~TTB;  //complement 
assign opb = ~OPB;  //complement 
assign oqa = ~OQA;  //complement 
assign oqb = ~OQB;  //complement 
assign ora = ~ORA;  //complement 
assign JPA =  HON & hpb & hpc  |  hon & HPB & hpc  |  hon & hpb & HPC  |  HON & HPB & HPC  ; 
assign jpa = ~JPA; //complement 
assign jpm =  HON & hpb & hpc  |  hon & HPB & hpc  |  hon & hpb & HPC  |  hon & hpb & hpc  ; 
assign JPM = ~jpm;  //complement 
assign kqa = ~KQA;  //complement 
assign KQM = ~kqm;  //complement 
assign oib = ~OIB;  //complement 
assign oja = ~OJA;  //complement 
assign okb = ~OKB;  //complement 
assign oma = ~OMA;  //complement 
assign kra = ~KRA;  //complement 
assign mrb = ~MRB;  //complement 
assign msa = ~MSA;  //complement 
assign LRA =  KQM & kra & krb  |  kqm & KRA & krb  |  kqm & kra & KRB  |  KQM & KRA & KRB  ; 
assign lra = ~LRA; //complement 
assign lrm =  KQM & kra & krb  |  kqm & KRA & krb  |  kqm & kra & KRB  |  kqm & kra & krb  ; 
assign LRM = ~lrm;  //complement 
assign ccu = ~CCU;  //complement 
assign orb = ~ORB;  //complement 
assign osa = ~OSA;  //complement 
assign JEA =  HDM & heb & hea  |  hdm & HEB & hea  |  hdm & heb & HEA  |  HDM & HEB & HEA  ; 
assign jea = ~JEA; //complement 
assign jem =  HDM & heb & hea  |  hdm & HEB & hea  |  hdm & heb & HEA  |  hdm & heb & hea  ; 
assign JEM = ~jem;  //complement 
assign ELL =  CDZ & DDL  ; 
assign ell = ~ELL;  //complement 
assign JCA =  HCA & hce & hbm  |  hca & HCE & hbm  |  hca & hce & HBM  |  HCA & HCE & HBM  ; 
assign jca = ~JCA; //complement 
assign jcm =  HCA & hce & hbm  |  hca & HCE & hbm  |  hca & hce & HBM  |  hca & hce & hbm  ; 
assign JCM = ~jcm;  //complement 
assign JDA =  HDA & hdd & hcm  |  hda & HDD & hcm  |  hda & hdd & HCM  |  HDA & HDD & HCM  ; 
assign jda = ~JDA; //complement 
assign jdm =  HDA & hdd & hcm  |  hda & HDD & hcm  |  hda & hdd & HCM  |  hda & hdd & hcm  ; 
assign JDM = ~jdm;  //complement 
assign kda = ~KDA;  //complement 
assign KDM = ~kdm;  //complement 
assign kaa = ~KAA;  //complement 
assign KAM = ~kam;  //complement 
assign kac = ~KAC;  //complement 
assign kca = ~KCA;  //complement 
assign KCM = ~kcm;  //complement 
assign kdc = ~KDC;  //complement 
assign kea = ~KEA;  //complement 
assign KEM = ~kem;  //complement 
assign kdb = ~KDB;  //complement 
assign oba = ~OBA;  //complement 
assign OBM = ~obm;  //complement 
assign maa = ~MAA;  //complement 
assign MAM = ~mam;  //complement 
assign LDA =  KCM & kdc & kdb  |  kcm & KDC & kdb  |  kcm & kdc & KDB  |  KCM & KDC & KDB  ; 
assign lda = ~LDA; //complement 
assign ldm =  KCM & kdc & kdb  |  kcm & KDC & kdb  |  kcm & kdc & KDB  |  kcm & kdc & kdb  ; 
assign LDM = ~ldm;  //complement 
assign NAA =  MAA & mac & mab  |  maa & MAC & mab  |  maa & mac & MAB  |  MAA & MAC & MAB  ; 
assign naa = ~NAA; //complement 
assign nam =  MAA & mac & mab  |  maa & MAC & mab  |  maa & mac & MAB  |  maa & mac & mab  ; 
assign NAM = ~nam;  //complement 
assign oaa = ~OAA;  //complement 
assign OAM = ~oam;  //complement 
assign NBA =  MAM & mba & mbb  |  mam & MBA & mbb  |  mam & mba & MBB  |  MAM & MBA & MBB  ; 
assign nba = ~NBA; //complement 
assign nbm =  MAM & mba & mbb  |  mam & MBA & mbb  |  mam & mba & MBB  |  mam & mba & mbb  ; 
assign NBM = ~nbm;  //complement 
assign JBB =  HAO & hbb & hbd  |  hao & HBB & hbd  |  hao & hbb & HBD  |  HAO & HBB & HBD  ; 
assign jbb = ~JBB; //complement 
assign jbn =  HAO & hbb & hbd  |  hao & HBB & hbd  |  hao & hbb & HBD  |  hao & hbb & hbd  ; 
assign JBN = ~jbn;  //complement 
assign LEA =  KDM & kea & keb  |  kdm & KEA & keb  |  kdm & kea & KEB  |  KDM & KEA & KEB  ; 
assign lea = ~LEA; //complement 
assign lem =  KDM & kea & keb  |  kdm & KEA & keb  |  kdm & kea & KEB  |  kdm & kea & keb  ; 
assign LEM = ~lem;  //complement 
assign JGB =  HFN & hge & hga  |  hfn & HGE & hga  |  hfn & hge & HGA  |  HFN & HGE & HGA  ; 
assign jgb = ~JGB; //complement 
assign jgn =  HFN & hge & hga  |  hfn & HGE & hga  |  hfn & hge & HGA  |  hfn & hge & hga  ; 
assign JGN = ~jgn;  //complement 
assign JCB =  HBN & hcc & hcb  |  hbn & HCC & hcb  |  hbn & hcc & HCB  |  HBN & HCC & HCB  ; 
assign jcb = ~JCB; //complement 
assign jcn =  HBN & hcc & hcb  |  hbn & HCC & hcb  |  hbn & hcc & HCB  |  hbn & hcc & hcb  ; 
assign JCN = ~jcn;  //complement 
assign mac = ~MAC;  //complement 
assign oca = ~OCA;  //complement 
assign OCM = ~ocm;  //complement 
assign JDC =  HCO & hdc & hcp  |  hco & HDC & hcp  |  hco & hdc & HCP  |  HCO & HDC & HCP  ; 
assign jdc = ~JDC; //complement 
assign jdo =  HCO & hdc & hcp  |  hco & HDC & hcp  |  hco & hdc & HCP  |  hco & hdc & hcp  ; 
assign JDO = ~jdo;  //complement 
assign kha = ~KHA;  //complement 
assign KHM = ~khm;  //complement 
assign meb = ~MEB;  //complement 
assign EPQ =  CDY & DDQ  ; 
assign epq = ~EPQ;  //complement 
assign EJP =  CDT & DDP  ; 
assign ejp = ~EJP;  //complement 
assign kcb = ~KCB;  //complement 
assign KCN = ~kcn;  //complement 
assign mda = ~MDA;  //complement 
assign MDM = ~mdm;  //complement 
assign mea = ~MEA;  //complement 
assign NEA =  MEB & mdm & mea  |  meb & MDM & mea  |  meb & mdm & MEA  |  MEB & MDM & MEA  ; 
assign nea = ~NEA; //complement 
assign nem =  MEB & mdm & mea  |  meb & MDM & mea  |  meb & mdm & MEA  |  meb & mdm & mea  ; 
assign NEM = ~nem;  //complement 
assign JMA =  HLM & hmc & hma  |  hlm & HMC & hma  |  hlm & hmc & HMA  |  HLM & HMC & HMA  ; 
assign jma = ~JMA; //complement 
assign jmm =  HLM & hmc & hma  |  hlm & HMC & hma  |  hlm & hmc & HMA  |  hlm & hmc & hma  ; 
assign JMM = ~jmm;  //complement 
assign kma = ~KMA;  //complement 
assign KMM = ~kmm;  //complement 
assign knb = ~KNB;  //complement 
assign LNA =  KMM & knb & kna  |  kmm & KNB & kna  |  kmm & knb & KNA  |  KMM & KNB & KNA  ; 
assign lna = ~LNA; //complement 
assign lnm =  KMM & knb & kna  |  kmm & KNB & kna  |  kmm & knb & KNA  |  kmm & knb & kna  ; 
assign LNM = ~lnm;  //complement 
assign JIA =  HIA & hhn & hib  |  hia & HHN & hib  |  hia & hhn & HIB  |  HIA & HHN & HIB  ; 
assign jia = ~JIA; //complement 
assign jim =  HIA & hhn & hib  |  hia & HHN & hib  |  hia & hhn & HIB  |  hia & hhn & hib  ; 
assign JIM = ~jim;  //complement 
assign LMA =  KMA & kmb & klm  |  kma & KMB & klm  |  kma & kmb & KLM  |  KMA & KMB & KLM  ; 
assign lma = ~LMA; //complement 
assign lmm =  KMA & kmb & klm  |  kma & KMB & klm  |  kma & kmb & KLM  |  kma & kmb & klm  ; 
assign LMM = ~lmm;  //complement 
assign JNA =  HNA & hmm & hnc  |  hna & HMM & hnc  |  hna & hmm & HNC  |  HNA & HMM & HNC  ; 
assign jna = ~JNA; //complement 
assign jnm =  HNA & hmm & hnc  |  hna & HMM & hnc  |  hna & hmm & HNC  |  hna & hmm & hnc  ; 
assign JNM = ~jnm;  //complement 
assign kja = ~KJA;  //complement 
assign KJM = ~kjm;  //complement 
assign kjc = ~KJC;  //complement 
assign LJA =  KJA & kjc & kim  |  kja & KJC & kim  |  kja & kjc & KIM  |  KJA & KJC & KIM  ; 
assign lja = ~LJA; //complement 
assign ljm =  KJA & kjc & kim  |  kja & KJC & kim  |  kja & kjc & KIM  |  kja & kjc & kim  ; 
assign LJM = ~ljm;  //complement 
assign kla = ~KLA;  //complement 
assign KLM = ~klm;  //complement 
assign kmb = ~KMB;  //complement 
assign kia = ~KIA;  //complement 
assign KIM = ~kim;  //complement 
assign kjb = ~KJB;  //complement 
assign mja = ~MJA;  //complement 
assign MJM = ~mjm;  //complement 
assign JLB =  HKO & hkn & hlc  |  hko & HKN & hlc  |  hko & hkn & HLC  |  HKO & HKN & HLC  ; 
assign jlb = ~JLB; //complement 
assign jln =  HKO & hkn & hlc  |  hko & HKN & hlc  |  hko & hkn & HLC  |  hko & hkn & hlc  ; 
assign JLN = ~jln;  //complement 
assign LOA =  KNM & kob & koa  |  knm & KOB & koa  |  knm & kob & KOA  |  KNM & KOB & KOA  ; 
assign loa = ~LOA; //complement 
assign lom =  KNM & kob & koa  |  knm & KOB & koa  |  knm & kob & KOA  |  knm & kob & koa  ; 
assign LOM = ~lom;  //complement 
assign JIB =  HID & hic & hho  |  hid & HIC & hho  |  hid & hic & HHO  |  HID & HIC & HHO  ; 
assign jib = ~JIB; //complement 
assign jin =  HID & hic & hho  |  hid & HIC & hho  |  hid & hic & HHO  |  hid & hic & hho  ; 
assign JIN = ~jin;  //complement 
assign JJB =  HJB & hio & hjd  |  hjb & HIO & hjd  |  hjb & hio & HJD  |  HJB & HIO & HJD  ; 
assign jjb = ~JJB; //complement 
assign jjn =  HJB & hio & hjd  |  hjb & HIO & hjd  |  hjb & hio & HJD  |  hjb & hio & hjd  ; 
assign JJN = ~jjn;  //complement 
assign JKA =  HJN & hkb & hkc  |  hjn & HKB & hkc  |  hjn & hkb & HKC  |  HJN & HKB & HKC  ; 
assign jka = ~JKA; //complement 
assign jkm =  HJN & hkb & hkc  |  hjn & HKB & hkc  |  hjn & hkb & HKC  |  hjn & hkb & hkc  ; 
assign JKM = ~jkm;  //complement 
assign kna = ~KNA;  //complement 
assign KNM = ~knm;  //complement 
assign kob = ~KOB;  //complement 
assign JHB =  HGN & hhc & hgo  |  hgn & HHC & hgo  |  hgn & hhc & HGO  |  HGN & HHC & HGO  ; 
assign jhb = ~JHB; //complement 
assign jhn =  HGN & hhc & hgo  |  hgn & HHC & hgo  |  hgn & hhc & HGO  |  hgn & hhc & hgo  ; 
assign JHN = ~jhn;  //complement 
assign kkb = ~KKB;  //complement 
assign kkc = ~KKC;  //complement 
assign JMB =  HMB & hlo & hln  |  hmb & HLO & hln  |  hmb & hlo & HLN  |  HMB & HLO & HLN  ; 
assign jmb = ~JMB; //complement 
assign jmn =  HMB & hlo & hln  |  hmb & HLO & hln  |  hmb & hlo & HLN  |  hmb & hlo & hln  ; 
assign JMN = ~jmn;  //complement 
assign oeb = ~OEB;  //complement 
assign ofa = ~OFA;  //complement 
assign mvb = ~MVB;  //complement 
assign mwa = ~MWA;  //complement 
assign mya = ~MYA;  //complement 
assign cay = ~CAY;  //complement 
assign cby = ~CBY;  //complement 
assign ccy = ~CCY;  //complement 
assign cdy = ~CDY;  //complement 
assign ovb = ~OVB;  //complement 
assign owa = ~OWA;  //complement 
assign oya = ~OYA;  //complement 
assign mma = ~MMA;  //complement 
assign mna = ~MNA;  //complement 
assign mnb = ~MNB;  //complement 
assign moa = ~MOA;  //complement 
assign kva = ~KVA;  //complement 
assign KVM = ~kvm;  //complement 
assign dbd = ~DBD;  //complement 
assign dcd = ~DCD;  //complement 
assign ddd = ~DDD;  //complement 
assign ona = ~ONA;  //complement 
assign onb = ~ONB;  //complement 
assign ooa = ~OOA;  //complement 
assign kta = ~KTA;  //complement 
assign KTM = ~ktm;  //complement 
assign kua = ~KUA;  //complement 
assign KUM = ~kum;  //complement 
assign kya = ~KYA;  //complement 
assign kza = ~KZA;  //complement 
assign kzb = ~KZB;  //complement 
assign daz = ~DAZ;  //complement 
assign dbz = ~DBZ;  //complement 
assign dcz = ~DCZ;  //complement 
assign mtb = ~MTB;  //complement 
assign mua = ~MUA;  //complement 
assign mub = ~MUB;  //complement 
assign mva = ~MVA;  //complement 
assign JUA =  HUB & huc & htm  |  hub & HUC & htm  |  hub & huc & HTM  |  HUB & HUC & HTM  ; 
assign jua = ~JUA; //complement 
assign jum =  HUB & huc & htm  |  hub & HUC & htm  |  hub & huc & HTM  |  hub & huc & htm  ; 
assign JUM = ~jum;  //complement 
assign otb = ~OTB;  //complement 
assign oua = ~OUA;  //complement 
assign oub = ~OUB;  //complement 
assign ova = ~OVA;  //complement 
assign ksa = ~KSA;  //complement 
assign KSM = ~ksm;  //complement 
assign mob = ~MOB;  //complement 
assign mpa = ~MPA;  //complement 
assign msb = ~MSB;  //complement 
assign mta = ~MTA;  //complement 
assign cak = ~CAK;  //complement 
assign cbk = ~CBK;  //complement 
assign cck = ~CCK;  //complement 
assign cdk = ~CDK;  //complement 
assign ojb = ~OJB;  //complement 
assign oka = ~OKA;  //complement 
assign JSA =  HRM & hrn & hsb  |  hrm & HRN & hsb  |  hrm & hrn & HSB  |  HRM & HRN & HSB  ; 
assign jsa = ~JSA; //complement 
assign jsm =  HRM & hrn & hsb  |  hrm & HRN & hsb  |  hrm & hrn & HSB  |  hrm & hrn & hsb  ; 
assign JSM = ~jsm;  //complement 
assign cao = ~CAO;  //complement 
assign cbo = ~CBO;  //complement 
assign cco = ~CCO;  //complement 
assign cdo = ~CDO;  //complement 
assign DHZ = ~dhz;  //complement 
assign trg = ~TRG;  //complement 
assign ota = ~OTA;  //complement 
assign omb = ~OMB;  //complement 
assign oob = ~OOB;  //complement 
assign opa = ~OPA;  //complement 
assign osb = ~OSB;  //complement 
assign ddz = ~DDZ;  //complement 
assign cam = ~CAM;  //complement 
assign cbm = ~CBM;  //complement 
assign ccm = ~CCM;  //complement 
assign cdm = ~CDM;  //complement 
assign mza = ~MZA;  //complement 
assign mzb = ~MZB;  //complement 
assign oza = ~OZA;  //complement 
assign ozb = ~OZB;  //complement 
assign JNB =  HNB & hmn & hnd  |  hnb & HMN & hnd  |  hnb & hmn & HND  |  HNB & HMN & HND  ; 
assign jnb = ~JNB; //complement 
assign jnn =  HNB & hmn & hnd  |  hnb & HMN & hnd  |  hnb & hmn & HND  |  hnb & hmn & hnd  ; 
assign JNN = ~jnn;  //complement 
assign can = ~CAN;  //complement 
assign cbn = ~CBN;  //complement 
assign ccn = ~CCN;  //complement 
assign cdn = ~CDN;  //complement 
assign DEZ = ~dez;  //complement 
assign DFZ = ~dfz;  //complement 
assign DGZ = ~dgz;  //complement 
assign hgc = ~HGC;  //complement 
assign HGO = ~hgo;  //complement 
assign GCA =  FCE & fbo & fcg  |  fce & FBO & fcg  |  fce & fbo & FCG  |  FCE & FBO & FCG  ; 
assign gca = ~GCA; //complement 
assign gcm =  FCE & fbo & fcg  |  fce & FBO & fcg  |  fce & fbo & FCG  |  fce & fbo & fcg  ; 
assign GCM = ~gcm;  //complement 
assign GDA =  FDG & fcs & fcq  |  fdg & FCS & fcq  |  fdg & fcs & FCQ  |  FDG & FCS & FCQ  ; 
assign gda = ~GDA; //complement 
assign gdm =  FDG & fcs & fcq  |  fdg & FCS & fcq  |  fdg & fcs & FCQ  |  fdg & fcs & fcq  ; 
assign GDM = ~gdm;  //complement 
assign GHA =  FHE & fgq & fgo  |  fhe & FGQ & fgo  |  fhe & fgq & FGO  |  FHE & FGQ & FGO  ; 
assign gha = ~GHA; //complement 
assign ghm =  FHE & fgq & fgo  |  fhe & FGQ & fgo  |  fhe & fgq & FGO  |  fhe & fgq & fgo  ; 
assign GHM = ~ghm;  //complement 
assign GBB =  FAM & fbe & fat  |  fam & FBE & fat  |  fam & fbe & FAT  |  FAM & FBE & FAT  ; 
assign gbb = ~GBB; //complement 
assign gbn =  FAM & fbe & fat  |  fam & FBE & fat  |  fam & fbe & FAT  |  fam & fbe & fat  ; 
assign GBN = ~gbn;  //complement 
assign hca = ~HCA;  //complement 
assign HCM = ~hcm;  //complement 
assign hce = ~HCE;  //complement 
assign hda = ~HDA;  //complement 
assign HDM = ~hdm;  //complement 
assign hdd = ~HDD;  //complement 
assign GGA =  FFO & fge & ffr  |  ffo & FGE & ffr  |  ffo & fge & FFR  |  FFO & FGE & FFR  ; 
assign gga = ~GGA; //complement 
assign ggm =  FFO & fge & ffr  |  ffo & FGE & ffr  |  ffo & fge & FFR  |  ffo & fge & ffr  ; 
assign GGM = ~ggm;  //complement 
assign hdc = ~HDC;  //complement 
assign HDO = ~hdo;  //complement 
assign heb = ~HEB;  //complement 
assign HEN = ~hen;  //complement 
assign hge = ~HGE;  //complement 
assign hhb = ~HHB;  //complement 
assign HHN = ~hhn;  //complement 
assign GBC =  FBG & faq & fba  |  fbg & FAQ & fba  |  fbg & faq & FBA  |  FBG & FAQ & FBA  ; 
assign gbc = ~GBC; //complement 
assign gbo =  FBG & faq & fba  |  fbg & FAQ & fba  |  fbg & faq & FBA  |  fbg & faq & fba  ; 
assign GBO = ~gbo;  //complement 
assign GDC =  FDE & fcm & fdd  |  fde & FCM & fdd  |  fde & fcm & FDD  |  FDE & FCM & FDD  ; 
assign gdc = ~GDC; //complement 
assign gdo =  FDE & fcm & fdd  |  fde & FCM & fdd  |  fde & fcm & FDD  |  fde & fcm & fdd  ; 
assign GDO = ~gdo;  //complement 
assign GEC =  FED & fdq & feg  |  fed & FDQ & feg  |  fed & fdq & FEG  |  FED & FDQ & FEG  ; 
assign gec = ~GEC; //complement 
assign geo =  FED & fdq & feg  |  fed & FDQ & feg  |  fed & fdq & FEG  |  fed & fdq & feg  ; 
assign GEO = ~geo;  //complement 
assign GHB =  FHC & fhh & fgm  |  fhc & FHH & fgm  |  fhc & fhh & FGM  |  FHC & FHH & FGM  ; 
assign ghb = ~GHB; //complement 
assign ghn =  FHC & fhh & fgm  |  fhc & FHH & fgm  |  fhc & fhh & FGM  |  fhc & fhh & fgm  ; 
assign GHN = ~ghn;  //complement 
assign GAB =  FAI & fae & faf  |  fai & FAE & faf  |  fai & fae & FAF  |  FAI & FAE & FAF  ; 
assign gab = ~GAB; //complement 
assign gan =  FAI & fae & faf  |  fai & FAE & faf  |  fai & fae & FAF  |  fai & fae & faf  ; 
assign GAN = ~gan;  //complement 
assign hbb = ~HBB;  //complement 
assign HBN = ~hbn;  //complement 
assign hbd = ~HBD;  //complement 
assign hfb = ~HFB;  //complement 
assign HFN = ~hfn;  //complement 
assign GFC =  FFG & fes & feq  |  ffg & FES & feq  |  ffg & fes & FEQ  |  FFG & FES & FEQ  ; 
assign gfc = ~GFC; //complement 
assign gfo =  FFG & fes & feq  |  ffg & FES & feq  |  ffg & fes & FEQ  |  ffg & fes & feq  ; 
assign GFO = ~gfo;  //complement 
assign GBD =  FAU & far & fbb  |  fau & FAR & fbb  |  fau & far & FBB  |  FAU & FAR & FBB  ; 
assign gbd = ~GBD; //complement 
assign gbp =  FAU & far & fbb  |  fau & FAR & fbb  |  fau & far & FBB  |  fau & far & fbb  ; 
assign GBP = ~gbp;  //complement 
assign hcc = ~HCC;  //complement 
assign HCO = ~hco;  //complement 
assign GED =  FEI & fee & fdr  |  fei & FEE & fdr  |  fei & fee & FDR  |  FEI & FEE & FDR  ; 
assign ged = ~GED; //complement 
assign gep =  FEI & fee & fdr  |  fei & FEE & fdr  |  fei & fee & FDR  |  fei & fee & fdr  ; 
assign GEP = ~gep;  //complement 
assign GHD =  FHD & fgn & fgs  |  fhd & FGN & fgs  |  fhd & fgn & FGS  |  FHD & FGN & FGS  ; 
assign ghd = ~GHD; //complement 
assign ghp =  FHD & fgn & fgs  |  fhd & FGN & fgs  |  fhd & fgn & FGS  |  fhd & fgn & fgs  ; 
assign GHP = ~ghp;  //complement 
assign hab = ~HAB;  //complement 
assign HAN = ~han;  //complement 
assign GDE =  FDH & fct & fdb  |  fdh & FCT & fdb  |  fdh & fct & FDB  |  FDH & FCT & FDB  ; 
assign gde = ~GDE; //complement 
assign gdq =  FDH & fct & fdb  |  fdh & FCT & fdb  |  fdh & fct & FDB  |  fdh & fct & fdb  ; 
assign GDQ = ~gdq;  //complement 
assign GCB =  FBS & fbq & fcc  |  fbs & FBQ & fcc  |  fbs & fbq & FCC  |  FBS & FBQ & FCC  ; 
assign gcb = ~GCB; //complement 
assign gcn =  FBS & fbq & fcc  |  fbs & FBQ & fcc  |  fbs & fbq & FCC  |  fbs & fbq & fcc  ; 
assign GCN = ~gcn;  //complement 
assign GBE =  FAS & fan & fbj  |  fas & FAN & fbj  |  fas & fan & FBJ  |  FAS & FAN & FBJ  ; 
assign gbe = ~GBE; //complement 
assign gbq =  FAS & fan & fbj  |  fas & FAN & fbj  |  fas & fan & FBJ  |  fas & fan & fbj  ; 
assign GBQ = ~gbq;  //complement 
assign GCE =  FBR & fcf & fbp  |  fbr & FCF & fbp  |  fbr & fcf & FBP  |  FBR & FCF & FBP  ; 
assign gce = ~GCE; //complement 
assign gcq =  FBR & fcf & fbp  |  fbr & FCF & fbp  |  fbr & fcf & FBP  |  fbr & fcf & fbp  ; 
assign GCQ = ~gcq;  //complement 
assign hcd = ~HCD;  //complement 
assign HCP = ~hcp;  //complement 
assign GFE =  FFE & fen & ffh  |  ffe & FEN & ffh  |  ffe & fen & FFH  |  FFE & FEN & FFH  ; 
assign gfe = ~GFE; //complement 
assign gfq =  FFE & fen & ffh  |  ffe & FEN & ffh  |  ffe & fen & FFH  |  ffe & fen & ffh  ; 
assign GFQ = ~gfq;  //complement 
assign GKA =  FJO & fkc & fkg  |  fjo & FKC & fkg  |  fjo & fkc & FKG  |  FJO & FKC & FKG  ; 
assign gka = ~GKA; //complement 
assign gkm =  FJO & fkc & fkg  |  fjo & FKC & fkg  |  fjo & fkc & FKG  |  fjo & fkc & fkg  ; 
assign GKM = ~gkm;  //complement 
assign hla = ~HLA;  //complement 
assign HLM = ~hlm;  //complement 
assign hmc = ~HMC;  //complement 
assign GTA =  FTB & fso & ftd  |  ftb & FSO & ftd  |  ftb & fso & FTD  |  FTB & FSO & FTD  ; 
assign gta = ~GTA; //complement 
assign gtm =  FTB & fso & ftd  |  ftb & FSO & ftd  |  ftb & fso & FTD  |  ftb & fso & ftd  ; 
assign GTM = ~gtm;  //complement 
assign GIA =  FIA & fhq & fie  |  fia & FHQ & fie  |  fia & fhq & FIE  |  FIA & FHQ & FIE  ; 
assign gia = ~GIA; //complement 
assign gim =  FIA & fhq & fie  |  fia & FHQ & fie  |  fia & fhq & FIE  |  fia & fhq & fie  ; 
assign GIM = ~gim;  //complement 
assign GLA =  FKO & flf & fld  |  fko & FLF & fld  |  fko & flf & FLD  |  FKO & FLF & FLD  ; 
assign gla = ~GLA; //complement 
assign glm =  FKO & flf & fld  |  fko & FLF & fld  |  fko & flf & FLD  |  fko & flf & fld  ; 
assign GLM = ~glm;  //complement 
assign GQA =  FQA & fpp & fqc  |  fqa & FPP & fqc  |  fqa & fpp & FQC  |  FQA & FPP & FQC  ; 
assign gqa = ~GQA; //complement 
assign gqm =  FQA & fpp & fqc  |  fqa & FPP & fqc  |  fqa & fpp & FQC  |  fqa & fpp & fqc  ; 
assign GQM = ~gqm;  //complement 
assign hia = ~HIA;  //complement 
assign HIM = ~him;  //complement 
assign GMA =  FLO & fma & fme  |  flo & FMA & fme  |  flo & fma & FME  |  FLO & FMA & FME  ; 
assign gma = ~GMA; //complement 
assign gmm =  FLO & fma & fme  |  flo & FMA & fme  |  flo & fma & FME  |  flo & fma & fme  ; 
assign GMM = ~gmm;  //complement 
assign hna = ~HNA;  //complement 
assign HNM = ~hnm;  //complement 
assign hqc = ~HQC;  //complement 
assign GIB =  FHO & fig & fif  |  fho & FIG & fif  |  fho & fig & FIF  |  FHO & FIG & FIF  ; 
assign gib = ~GIB; //complement 
assign gin =  FHO & fig & fif  |  fho & FIG & fif  |  fho & fig & FIF  |  fho & fig & fif  ; 
assign GIN = ~gin;  //complement 
assign hib = ~HIB;  //complement 
assign HIN = ~hin;  //complement 
assign hjc = ~HJC;  //complement 
assign hma = ~HMA;  //complement 
assign HMM = ~hmm;  //complement 
assign GNB =  FND & fne & fna  |  fnd & FNE & fna  |  fnd & fne & FNA  |  FND & FNE & FNA  ; 
assign gnb = ~GNB; //complement 
assign gnn =  FND & fne & fna  |  fnd & FNE & fna  |  fnd & fne & FNA  |  fnd & fne & fna  ; 
assign GNN = ~gnn;  //complement 
assign hic = ~HIC;  //complement 
assign HIO = ~hio;  //complement 
assign GLB =  FKQ & flc & flb  |  fkq & FLC & flb  |  fkq & flc & FLB  |  FKQ & FLC & FLB  ; 
assign glb = ~GLB; //complement 
assign gln =  FKQ & flc & flb  |  fkq & FLC & flb  |  fkq & flc & FLB  |  fkq & flc & flb  ; 
assign GLN = ~gln;  //complement 
assign hkb = ~HKB;  //complement 
assign HKN = ~hkn;  //complement 
assign hnc = ~HNC;  //complement 
assign GIC =  FHN & fhp & fid  |  fhn & FHP & fid  |  fhn & fhp & FID  |  FHN & FHP & FID  ; 
assign gic = ~GIC; //complement 
assign gio =  FHN & fhp & fid  |  fhn & FHP & fid  |  fhn & fhp & FID  |  fhn & fhp & fid  ; 
assign GIO = ~gio;  //complement 
assign GKC =  FKA & fjp & fjr  |  fka & FJP & fjr  |  fka & fjp & FJR  |  FKA & FJP & FJR  ; 
assign gkc = ~GKC; //complement 
assign gko =  FKA & fjp & fjr  |  fka & FJP & fjr  |  fka & fjp & FJR  |  fka & fjp & fjr  ; 
assign GKO = ~gko;  //complement 
assign GMB =  FLQ & fmd & fln  |  flq & FMD & fln  |  flq & fmd & FLN  |  FLQ & FMD & FLN  ; 
assign gmb = ~GMB; //complement 
assign gmn =  FLQ & fmd & fln  |  flq & FMD & fln  |  flq & fmd & FLN  |  flq & fmd & fln  ; 
assign GMN = ~gmn;  //complement 
assign hhc = ~HHC;  //complement 
assign HHO = ~hho;  //complement 
assign hjd = ~HJD;  //complement 
assign hjb = ~HJB;  //complement 
assign HJN = ~hjn;  //complement 
assign hlc = ~HLC;  //complement 
assign HLO = ~hlo;  //complement 
assign hpc = ~HPC;  //complement 
assign GGD =  FFQ & fgf & ffp  |  ffq & FGF & ffp  |  ffq & fgf & FFP  |  FFQ & FGF & FFP  ; 
assign ggd = ~GGD; //complement 
assign ggp =  FFQ & fgf & ffp  |  ffq & FGF & ffp  |  ffq & fgf & FFP  |  ffq & fgf & ffp  ; 
assign GGP = ~ggp;  //complement 
assign GJD =  FIO & fin & fje  |  fio & FIN & fje  |  fio & fin & FJE  |  FIO & FIN & FJE  ; 
assign gjd = ~GJD; //complement 
assign gjp =  FIO & fin & fje  |  fio & FIN & fje  |  fio & fin & FJE  |  fio & fin & fje  ; 
assign GJP = ~gjp;  //complement 
assign GLC =  FLE & fkp & fla  |  fle & FKP & fla  |  fle & fkp & FLA  |  FLE & FKP & FLA  ; 
assign glc = ~GLC; //complement 
assign glo =  FLE & fkp & fla  |  fle & FKP & fla  |  fle & fkp & FLA  |  fle & fkp & fla  ; 
assign GLO = ~glo;  //complement 
assign GXA =  FXA & fxb & fwm  |  fxa & FXB & fwm  |  fxa & fxb & FWM  |  FXA & FXB & FWM  ; 
assign gxa = ~GXA; //complement 
assign gxm =  FXA & fxb & fwm  |  fxa & FXB & fwm  |  fxa & fxb & FWM  |  fxa & fxb & fwm  ; 
assign GXM = ~gxm;  //complement 
assign hua = ~HUA;  //complement 
assign HUM = ~hum;  //complement 
assign htc = ~HTC;  //complement 
assign qax = ~QAX;  //complement 
assign caz = ~CAZ;  //complement 
assign cbz = ~CBZ;  //complement 
assign ccz = ~CCZ;  //complement 
assign cdz = ~CDZ;  //complement 
assign GUA =  FUB & fua & fuc  |  fub & FUA & fuc  |  fub & fua & FUC  |  FUB & FUA & FUC  ; 
assign gua = ~GUA; //complement 
assign gum =  FUB & fua & fuc  |  fub & FUA & fuc  |  fub & fua & FUC  |  fub & fua & fuc  ; 
assign GUM = ~gum;  //complement 
assign GZA =  FZA & fzb & fym  |  fza & FZB & fym  |  fza & fzb & FYM  |  FZA & FZB & FYM  ; 
assign gza = ~GZA; //complement 
assign gzm =  FZA & fzb & fym  |  fza & FZB & fym  |  fza & fzb & FYM  |  fza & fzb & fym  ; 
assign GZM = ~gzm;  //complement 
assign QAK = ~qak;  //complement 
assign QAL = ~qal;  //complement 
assign dae = ~DAE;  //complement 
assign dce = ~DCE;  //complement 
assign dde = ~DDE;  //complement 
assign hya = ~HYA;  //complement 
assign HYM = ~hym;  //complement 
assign hza = ~HZA;  //complement 
assign qao = ~QAO;  //complement 
assign qar = ~QAR;  //complement 
assign qau = ~QAU;  //complement 
assign qaz = ~QAZ;  //complement 
assign kzm = ~KZM;  //complement 
assign ozm = ~OZM;  //complement 
assign qia = ~QIA;  //complement 
assign GTB =  FSN & ftc & fta  |  fsn & FTC & fta  |  fsn & ftc & FTA  |  FSN & FTC & FTA  ; 
assign gtb = ~GTB; //complement 
assign gtn =  FSN & ftc & fta  |  fsn & FTC & fta  |  fsn & ftc & FTA  |  fsn & ftc & fta  ; 
assign GTN = ~gtn;  //complement 
assign hub = ~HUB;  //complement 
assign huc = ~HUC;  //complement 
assign hxb = ~HXB;  //complement 
assign QAH = ~qah;  //complement 
assign QAI = ~qai;  //complement 
assign caw = ~CAW;  //complement 
assign cbw = ~CBW;  //complement 
assign ccw = ~CCW;  //complement 
assign cdw = ~CDW;  //complement 
assign GRB =  FRC & frd & fqn  |  frc & FRD & fqn  |  frc & frd & FQN  |  FRC & FRD & FQN  ; 
assign grb = ~GRB; //complement 
assign grn =  FRC & frd & fqn  |  frc & FRD & fqn  |  frc & frd & FQN  |  frc & frd & fqn  ; 
assign GRN = ~grn;  //complement 
assign qib = ~QIB;  //complement 
assign qic = ~QIC;  //complement 
assign qid = ~QID;  //complement 
assign qie = ~QIE;  //complement 
assign car = ~CAR;  //complement 
assign cbr = ~CBR;  //complement 
assign ccr = ~CCR;  //complement 
assign cdr = ~CDR;  //complement 
assign hrb = ~HRB;  //complement 
assign HRN = ~hrn;  //complement 
assign hsb = ~HSB;  //complement 
assign QAE = ~qae;  //complement 
assign QAF = ~qaf;  //complement 
assign GOC =  FOD & foe & fno  |  fod & FOE & fno  |  fod & foe & FNO  |  FOD & FOE & FNO  ; 
assign goc = ~GOC; //complement 
assign goo =  FOD & foe & fno  |  fod & FOE & fno  |  fod & foe & FNO  |  fod & foe & fno  ; 
assign GOO = ~goo;  //complement 
assign hzm = ~HZM;  //complement 
assign mzm = ~MZM;  //complement 
assign hmb = ~HMB;  //complement 
assign HMN = ~hmn;  //complement 
assign hnd = ~HND;  //complement 
assign trh = ~TRH;  //complement 
assign QAA = ~qaa;  //complement 
assign QAB = ~qab;  //complement 
assign QAC = ~qac;  //complement 
assign cal = ~CAL;  //complement 
assign cbl = ~CBL;  //complement 
assign ccl = ~CCL;  //complement 
assign cdl = ~CDL;  //complement 
assign EBW =  CCE & DGW  ; 
assign ebw = ~EBW;  //complement 
assign EBX =  CCD & DGX  ; 
assign ebx = ~EBX;  //complement 
assign EBY =  CCC & DGY  ; 
assign eby = ~EBY;  //complement 
assign ECC =  CCZ & DCC  ; 
assign ecc = ~ECC;  //complement 
assign ECD =  CCY & DCD  ; 
assign ecd = ~ECD;  //complement 
assign ECE =  CCX & DCE  ; 
assign ece = ~ECE;  //complement 
assign EGG =  CCZ & DCG  ; 
assign egg = ~EGG;  //complement 
assign EGH =  CCY & DCH  ; 
assign egh = ~EGH;  //complement 
assign EGI =  CCX & DCI  ; 
assign egi = ~EGI;  //complement 
assign EKK =  CCZ & DCK  ; 
assign ekk = ~EKK;  //complement 
assign EKL =  CCY & DCL  ; 
assign ekl = ~EKL;  //complement 
assign EKM =  CCX & DCM  ; 
assign ekm = ~EKM;  //complement 
assign fbe = ~FBE;  //complement 
assign FBQ = ~fbq;  //complement 
assign fce = ~FCE;  //complement 
assign FCQ = ~fcq;  //complement 
assign fge = ~FGE;  //complement 
assign FGQ = ~fgq;  //complement 
assign fkc = ~FKC;  //complement 
assign FKO = ~fko;  //complement 
assign EAS =  CCH & DGS  ; 
assign eas = ~EAS;  //complement 
assign EAT =  CCG & DGT  ; 
assign eat = ~EAT;  //complement 
assign EAU =  CCF & DGU  ; 
assign eau = ~EAU;  //complement 
assign EDG =  CCW & DCG  ; 
assign edg = ~EDG;  //complement 
assign EDH =  CCV & DCH  ; 
assign edh = ~EDH;  //complement 
assign EDI =  CCU & DCI  ; 
assign edi = ~EDI;  //complement 
assign EEW =  CCH & DGW  ; 
assign eew = ~EEW;  //complement 
assign EEX =  CCG & DGX  ; 
assign eex = ~EEX;  //complement 
assign EEY =  CCF & DGY  ; 
assign eey = ~EEY;  //complement 
assign EHK =  CCW & DCK  ; 
assign ehk = ~EHK;  //complement 
assign EHL =  CCV & DCL  ; 
assign ehl = ~EHL;  //complement 
assign EHM =  CCU & DCM  ; 
assign ehm = ~EHM;  //complement 
assign fae = ~FAE;  //complement 
assign FAQ = ~faq;  //complement 
assign fei = ~FEI;  //complement 
assign fde = ~FDE;  //complement 
assign FDQ = ~fdq;  //complement 
assign fed = ~FED;  //complement 
assign FEP = ~fep;  //complement 
assign fhc = ~FHC;  //complement 
assign FHO = ~fho;  //complement 
assign fhh = ~FHH;  //complement 
assign EAG =  CCT & DCG  ; 
assign eag = ~EAG;  //complement 
assign EAH =  CCS & DCH  ; 
assign eah = ~EAH;  //complement 
assign EAI =  CCR & DCI  ; 
assign eai = ~EAI;  //complement 
assign EDS =  CCK & DGS  ; 
assign eds = ~EDS;  //complement 
assign EDT =  CCJ & DGT  ; 
assign edt = ~EDT;  //complement 
assign EDU =  CCI & DGU  ; 
assign edu = ~EDU;  //complement 
assign EEK =  CCT & DGK  ; 
assign eek = ~EEK;  //complement 
assign EEL =  CCS & DGL  ; 
assign eel = ~EEL;  //complement 
assign EEM =  CCR & DGM  ; 
assign eem = ~EEM;  //complement 
assign EHW =  CCK & DGW  ; 
assign ehw = ~EHW;  //complement 
assign EHX =  CCJ & DGX  ; 
assign ehx = ~EHX;  //complement 
assign EHY =  CCI & DGY  ; 
assign ehy = ~EHY;  //complement 
assign faf = ~FAF;  //complement 
assign FAR = ~far;  //complement 
assign fdf = ~FDF;  //complement 
assign FDR = ~fdr;  //complement 
assign fee = ~FEE;  //complement 
assign FEQ = ~feq;  //complement 
assign fhd = ~FHD;  //complement 
assign FHP = ~fhp;  //complement 
assign ffh = ~FFH;  //complement 
assign EAY =  CCB & DKY  ; 
assign eay = ~EAY;  //complement 
assign EAZ =  CCA & DGZ  ; 
assign eaz = ~EAZ;  //complement 
assign EBK =  CCQ & DGK  ; 
assign ebk = ~EBK;  //complement 
assign EBL =  CCP & DGL  ; 
assign ebl = ~EBL;  //complement 
assign EBM =  CCO & DGM  ; 
assign ebm = ~EBM;  //complement 
assign ECO =  CCN & DGO  ; 
assign eco = ~ECO;  //complement 
assign ECP =  CCM & DGP  ; 
assign ecp = ~ECP;  //complement 
assign ECQ =  CCL & DGQ  ; 
assign ecq = ~ECQ;  //complement 
assign EFO =  CCQ & DGO  ; 
assign efo = ~EFO;  //complement 
assign EFP =  CCP & DGP  ; 
assign efp = ~EFP;  //complement 
assign EFQ =  CCO & DGQ  ; 
assign efq = ~EFQ;  //complement 
assign fag = ~FAG;  //complement 
assign FAS = ~fas;  //complement 
assign fbj = ~FBJ;  //complement 
assign fbf = ~FBF;  //complement 
assign FBR = ~fbr;  //complement 
assign fci = ~FCI;  //complement 
assign fcf = ~FCF;  //complement 
assign FCR = ~fcr;  //complement 
assign ffe = ~FFE;  //complement 
assign FFQ = ~ffq;  //complement 
assign EOO =  CCZ & DCO  ; 
assign eoo = ~EOO;  //complement 
assign EOP =  CCY & DCP  ; 
assign eop = ~EOP;  //complement 
assign EOQ =  CCX & DCQ  ; 
assign eoq = ~EOQ;  //complement 
assign hxa = ~HXA;  //complement 
assign ESS =  CCZ & DCS  ; 
assign ess = ~ESS;  //complement 
assign EST =  CCY & DCT  ; 
assign est = ~EST;  //complement 
assign ESU =  CCX & DCU  ; 
assign esu = ~ESU;  //complement 
assign EWW =  CCZ & DCW  ; 
assign eww = ~EWW;  //complement 
assign EWX =  CCY & DCX  ; 
assign ewx = ~EWX;  //complement 
assign EWY =  CCX & DCY  ; 
assign ewy = ~EWY;  //complement 
assign foc = ~FOC;  //complement 
assign FOO = ~foo;  //complement 
assign fkg = ~FKG;  //complement 
assign fsc = ~FSC;  //complement 
assign FSO = ~fso;  //complement 
assign flf = ~FLF;  //complement 
assign fwa = ~FWA;  //complement 
assign FWM = ~fwm;  //complement 
assign fzb = ~FZB;  //complement 
assign ELO =  CCW & DCO  ; 
assign elo = ~ELO;  //complement 
assign ELP =  CCV & DCP  ; 
assign elp = ~ELP;  //complement 
assign ELQ =  CCU & DCQ  ; 
assign elq = ~ELQ;  //complement 
assign EJS =  CCQ & DCS  ; 
assign ejs = ~EJS;  //complement 
assign EJT =  CCP & DCT  ; 
assign ejt = ~EJT;  //complement 
assign EJU =  CCO & DCU  ; 
assign eju = ~EJU;  //complement 
assign EPS =  CCW & DCS  ; 
assign eps = ~EPS;  //complement 
assign EPT =  CCV & DCT  ; 
assign ept = ~EPT;  //complement 
assign EPU =  CCU & DCU  ; 
assign epu = ~EPU;  //complement 
assign ETW =  CCW & DCW  ; 
assign etw = ~ETW;  //complement 
assign ETX =  CCV & DCX  ; 
assign etx = ~ETX;  //complement 
assign ETY =  CCU & DCY  ; 
assign ety = ~ETY;  //complement 
assign flc = ~FLC;  //complement 
assign FLO = ~flo;  //complement 
assign fig = ~FIG;  //complement 
assign fpc = ~FPC;  //complement 
assign FPO = ~fpo;  //complement 
assign fta = ~FTA;  //complement 
assign FTM = ~ftm;  //complement 
assign fne = ~FNE;  //complement 
assign EIO =  CCT & DGO  ; 
assign eio = ~EIO;  //complement 
assign EIP =  CCS & DCP  ; 
assign eip = ~EIP;  //complement 
assign EIQ =  CCR & DCQ  ; 
assign eiq = ~EIQ;  //complement 
assign EMS =  CCT & DCS  ; 
assign ems = ~EMS;  //complement 
assign EMT =  CCS & DCT  ; 
assign emt = ~EMT;  //complement 
assign EMU =  CCR & DCU  ; 
assign emu = ~EMU;  //complement 
assign ENZ =  CCN & DCZ  ; 
assign enz = ~ENZ;  //complement 
assign fid = ~FID;  //complement 
assign FIP = ~fip;  //complement 
assign fmd = ~FMD;  //complement 
assign FMP = ~fmp;  //complement 
assign EGS =  CCN & DGS  ; 
assign egs = ~EGS;  //complement 
assign EGT =  CCM & DGT  ; 
assign egt = ~EGT;  //complement 
assign EGU =  CCL & DGU  ; 
assign egu = ~EGU;  //complement 
assign EKW =  CCN & DCW  ; 
assign ekw = ~EKW;  //complement 
assign EKX =  CCM & DCX  ; 
assign ekx = ~EKX;  //complement 
assign EKY =  CCL & DCY  ; 
assign eky = ~EKY;  //complement 
assign fgf = ~FGF;  //complement 
assign FGR = ~fgr;  //complement 
assign fje = ~FJE;  //complement 
assign FJQ = ~fjq;  //complement 
assign fkd = ~FKD;  //complement 
assign FKP = ~fkp;  //complement 
assign EZZ =  CCZ & DCZ  ; 
assign ezz = ~EZZ;  //complement 
assign cae = ~CAE;  //complement 
assign cbe = ~CBE;  //complement 
assign cce = ~CCE;  //complement 
assign cbc = ~CBC;  //complement 
assign ccc = ~CCC;  //complement 
assign cdc = ~CDC;  //complement 
assign dai = ~DAI;  //complement 
assign dci = ~DCI;  //complement 
assign ddi = ~DDI;  //complement 
assign CDE = ~cde;  //complement 
assign CDH = ~cdh;  //complement 
assign cat = ~CAT;  //complement 
assign dbh = ~DBH;  //complement 
assign dch = ~DCH;  //complement 
assign ddh = ~DDH;  //complement 
assign EQX =  CCS & DCX  ; 
assign eqx = ~EQX;  //complement 
assign DGU = ~dgu;  //complement 
assign DGX = ~dgx;  //complement 
assign DHU = ~dhu;  //complement 
assign DHX = ~dhx;  //complement 
assign DGL = ~dgl;  //complement 
assign DHL = ~dhl;  //complement 
assign DKY = ~dky;  //complement 
assign cah = ~CAH;  //complement 
assign cbh = ~CBH;  //complement 
assign cch = ~CCH;  //complement 
assign dam = ~DAM;  //complement 
assign dcm = ~DCM;  //complement 
assign ddm = ~DDM;  //complement 
assign dem = ~DEM;  //complement 
assign DGM = ~dgm;  //complement 
assign DGY = ~dgy;  //complement 
assign DHM = ~dhm;  //complement 
assign DHY = ~dhy;  //complement 
assign cas = ~CAS;  //complement 
assign cbs = ~CBS;  //complement 
assign ccs = ~CCS;  //complement 
assign cds = ~CDS;  //complement 
assign EQW =  CCT & DCW  ; 
assign eqw = ~EQW;  //complement 
assign EQY =  CCR & DCY  ; 
assign eqy = ~EQY;  //complement 
assign day = ~DAY;  //complement 
assign dcy = ~DCY;  //complement 
assign ddy = ~DDY;  //complement 
assign dey = ~DEY;  //complement 
assign caj = ~CAJ;  //complement 
assign cbj = ~CBJ;  //complement 
assign ccj = ~CCJ;  //complement 
assign cca = ~CCA;  //complement 
assign CDJ = ~cdj;  //complement 
assign fqb = ~FQB;  //complement 
assign FQN = ~fqn;  //complement 
assign dau = ~DAU;  //complement 
assign dcu = ~DCU;  //complement 
assign ddu = ~DDU;  //complement 
assign deu = ~DEU;  //complement 
assign cbt = ~CBT;  //complement 
assign cct = ~CCT;  //complement 
assign cdt = ~CDT;  //complement 
assign trc = ~TRC;  //complement 
assign ENW =  CCQ & DCW  ; 
assign enw = ~ENW;  //complement 
assign ENX =  CCP & DCX  ; 
assign enx = ~ENX;  //complement 
assign ENY =  CCO & DCY  ; 
assign eny = ~ENY;  //complement 
assign dbx = ~DBX;  //complement 
assign dcx = ~DCX;  //complement 
assign ddx = ~DDX;  //complement 
assign dfx = ~DFX;  //complement 
assign dbl = ~DBL;  //complement 
assign dcl = ~DCL;  //complement 
assign ddl = ~DDL;  //complement 
assign dfl = ~DFL;  //complement 
assign fnc = ~FNC;  //complement 
assign FNO = ~fno;  //complement 
assign dbt = ~DBT;  //complement 
assign dct = ~DCT;  //complement 
assign ddt = ~DDT;  //complement 
assign dft = ~DFT;  //complement 
assign DGT = ~dgt;  //complement 
assign DHT = ~dht;  //complement 
assign fcg = ~FCG;  //complement 
assign FCS = ~fcs;  //complement 
assign fbi = ~FBI;  //complement 
assign fdg = ~FDG;  //complement 
assign FDS = ~fds;  //complement 
assign fhe = ~FHE;  //complement 
assign FHQ = ~fhq;  //complement 
assign EBZ =  CDB & DHZ  ; 
assign ebz = ~EBZ;  //complement 
assign ECX =  CDE & DHX  ; 
assign ecx = ~ECX;  //complement 
assign ECY =  CDD & DHY  ; 
assign ecy = ~ECY;  //complement 
assign ECZ =  CDC & DHZ  ; 
assign ecz = ~ECZ;  //complement 
assign EDD =  CDZ & DDD  ; 
assign edd = ~EDD;  //complement 
assign EDE =  CDY & DDE  ; 
assign ede = ~EDE;  //complement 
assign EDF =  CDX & DDF  ; 
assign edf = ~EDF;  //complement 
assign EHH =  CDZ & DDH  ; 
assign ehh = ~EHH;  //complement 
assign EHI =  CDY & DDI  ; 
assign ehi = ~EHI;  //complement 
assign EHJ =  CDX & DDJ  ; 
assign ehj = ~EHJ;  //complement 
assign fah = ~FAH;  //complement 
assign FAT = ~fat;  //complement 
assign fbg = ~FBG;  //complement 
assign FBS = ~fbs;  //complement 
assign fef = ~FEF;  //complement 
assign FER = ~fer;  //complement 
assign fff = ~FFF;  //complement 
assign FFR = ~ffr;  //complement 
assign EAD =  CDW & DDD  ; 
assign ead = ~EAD;  //complement 
assign EAE =  CDV & DDE  ; 
assign eae = ~EAE;  //complement 
assign EAF =  CDU & DDF  ; 
assign eaf = ~EAF;  //complement 
assign EBT =  CDH & DHT  ; 
assign ebt = ~EBT;  //complement 
assign EBU =  CDG & DHU  ; 
assign ebu = ~EBU;  //complement 
assign EBV =  CDF & DHV  ; 
assign ebv = ~EBV;  //complement 
assign EEH =  CDW & DDH  ; 
assign eeh = ~EEH;  //complement 
assign EEI =  CDV & DDI  ; 
assign eei = ~EEI;  //complement 
assign EEJ =  CDU & DDJ  ; 
assign eej = ~EEJ;  //complement 
assign EFX =  CDH & DHX  ; 
assign efx = ~EFX;  //complement 
assign EFY =  CDG & DHY  ; 
assign efy = ~EFY;  //complement 
assign EFZ =  CDF & DHZ  ; 
assign efz = ~EFZ;  //complement 
assign fai = ~FAI;  //complement 
assign FAU = ~fau;  //complement 
assign fbh = ~FBH;  //complement 
assign FBT = ~fbt;  //complement 
assign feg = ~FEG;  //complement 
assign FES = ~fes;  //complement 
assign ffg = ~FFG;  //complement 
assign FFS = ~ffs;  //complement 
assign EAQ =  CDJ & DHQ  ; 
assign eaq = ~EAQ;  //complement 
assign EAR =  CDI & DHR  ; 
assign ear = ~EAR;  //complement 
assign EAP =  CDK & DHP  ; 
assign eap = ~EAP;  //complement 
assign EBH =  CDT & DDH  ; 
assign ebh = ~EBH;  //complement 
assign EBI =  CDS & DDI  ; 
assign ebi = ~EBI;  //complement 
assign EBJ =  CDR & DDJ  ; 
assign ebj = ~EBJ;  //complement 
assign EET =  CDK & DHT  ; 
assign eet = ~EET;  //complement 
assign EEU =  CDJ & DHU  ; 
assign eeu = ~EEU;  //complement 
assign EEV =  CDI & DHV  ; 
assign eev = ~EEV;  //complement 
assign EFL =  CDT & DHL  ; 
assign efl = ~EFL;  //complement 
assign EFM =  CDS & DHM  ; 
assign efm = ~EFM;  //complement 
assign EFN =  CDR & DHN  ; 
assign efn = ~EFN;  //complement 
assign fch = ~FCH;  //complement 
assign FCT = ~fct;  //complement 
assign fdh = ~FDH;  //complement 
assign FDT = ~fdt;  //complement 
assign fgg = ~FGG;  //complement 
assign FGS = ~fgs;  //complement 
assign fhf = ~FHF;  //complement 
assign FHR = ~fhr;  //complement 
assign ECL =  CDQ & DHL  ; 
assign ecl = ~ECL;  //complement 
assign ECM =  CDP & DHM  ; 
assign ecm = ~ECM;  //complement 
assign ECN =  CDO & DHN  ; 
assign ecn = ~ECN;  //complement 
assign EDP =  CDN & DHP  ; 
assign edp = ~EDP;  //complement 
assign EDQ =  CDM & DHQ  ; 
assign edq = ~EDQ;  //complement 
assign EDR =  CDL & DHR  ; 
assign edr = ~EDR;  //complement 
assign EGP =  CDQ & DHP  ; 
assign egp = ~EGP;  //complement 
assign EGQ =  CDP & DHQ  ; 
assign egq = ~EGQ;  //complement 
assign EGR =  CDO & DHR  ; 
assign egr = ~EGR;  //complement 
assign EHT =  CDN & DHT  ; 
assign eht = ~EHT;  //complement 
assign EHU =  CDM & DHU  ; 
assign ehu = ~EHU;  //complement 
assign EHV =  CDL & DHV  ; 
assign ehv = ~EHV;  //complement 
assign fld = ~FLD;  //complement 
assign FLP = ~flp;  //complement 
assign fpd = ~FPD;  //complement 
assign FPP = ~fpp;  //complement 
assign ftb = ~FTB;  //complement 
assign FTN = ~ftn;  //complement 
assign ELM =  CDY & DDM  ; 
assign elm = ~ELM;  //complement 
assign EPP =  CDZ & DDP  ; 
assign epp = ~EPP;  //complement 
assign EPR =  CDX & DDR  ; 
assign epr = ~EPR;  //complement 
assign ETT =  CDZ & DDT  ; 
assign ett = ~ETT;  //complement 
assign ETU =  CDY & DDU  ; 
assign etu = ~ETU;  //complement 
assign ETV =  CDX & DDV  ; 
assign etv = ~ETV;  //complement 
assign fie = ~FIE;  //complement 
assign FIQ = ~fiq;  //complement 
assign fme = ~FME;  //complement 
assign FMQ = ~fmq;  //complement 
assign fqc = ~FQC;  //complement 
assign FQO = ~fqo;  //complement 
assign EIL =  CDW & DDL  ; 
assign eil = ~EIL;  //complement 
assign EIM =  CDV & DDM  ; 
assign eim = ~EIM;  //complement 
assign EIN =  CDU & DDN  ; 
assign ein = ~EIN;  //complement 
assign EMP =  CDW & DDP  ; 
assign emp = ~EMP;  //complement 
assign EMQ =  CDV & DDQ  ; 
assign emq = ~EMQ;  //complement 
assign EMR =  CDU & DDR  ; 
assign emr = ~EMR;  //complement 
assign EQT =  CDW & DDT  ; 
assign eqt = ~EQT;  //complement 
assign EQU =  CDV & DDU  ; 
assign equ = ~EQU;  //complement 
assign EQV =  CDU & DDV  ; 
assign eqv = ~EQV;  //complement 
assign fif = ~FIF;  //complement 
assign FIR = ~fir;  //complement 
assign fjf = ~FJF;  //complement 
assign FJR = ~fjr;  //complement 
assign fnd = ~FND;  //complement 
assign FNP = ~fnp;  //complement 
assign frd = ~FRD;  //complement 
assign EIX =  CDK & DHX  ; 
assign eix = ~EIX;  //complement 
assign EIY =  CDJ & DHY  ; 
assign eiy = ~EIY;  //complement 
assign EIZ =  CDI & DHZ  ; 
assign eiz = ~EIZ;  //complement 
assign EJQ =  CDS & DDQ  ; 
assign ejq = ~EJQ;  //complement 
assign EJR =  CDR & DDR  ; 
assign ejr = ~EJR;  //complement 
assign ENT =  CDT & DDT  ; 
assign ent = ~ENT;  //complement 
assign ENU =  CDS & DDU  ; 
assign enu = ~ENU;  //complement 
assign ENV =  CDR & DDV  ; 
assign env = ~ENV;  //complement 
assign fke = ~FKE;  //complement 
assign FKQ = ~fkq;  //complement 
assign fle = ~FLE;  //complement 
assign FLQ = ~flq;  //complement 
assign fod = ~FOD;  //complement 
assign FOP = ~fop;  //complement 
assign foe = ~FOE;  //complement 
assign EKT =  CDQ & DHT  ; 
assign ekt = ~EKT;  //complement 
assign EKV =  CDO & DHV  ; 
assign ekv = ~EKV;  //complement 
assign EKU =  CDP & DHU  ; 
assign eku = ~EKU;  //complement 
assign ELX =  CDN & DDX  ; 
assign elx = ~ELX;  //complement 
assign ELY =  CDM & DDY  ; 
assign ely = ~ELY;  //complement 
assign ELZ =  CDL & DDZ  ; 
assign elz = ~ELZ;  //complement 
assign EOX =  CDQ & DDX  ; 
assign eox = ~EOX;  //complement 
assign EOY =  CDP & DDY  ; 
assign eoy = ~EOY;  //complement 
assign EOZ =  CDO & DDZ  ; 
assign eoz = ~EOZ;  //complement 
assign fxa = ~FXA;  //complement 
assign FXM = ~fxm;  //complement 
assign fza = ~FZA;  //complement 
assign EXX =  CDZ & DDX  ; 
assign exx = ~EXX;  //complement 
assign EXY =  CDY & DDY  ; 
assign exy = ~EXY;  //complement 
assign EXZ =  CDX & DDZ  ; 
assign exz = ~EXZ;  //complement 
assign fub = ~FUB;  //complement 
assign FUN = ~fun;  //complement 
assign LKA =  KKA & kkb & kkc  |  kka & KKB & kkc  |  kka & kkb & KKC  |  KKA & KKB & KKC  ; 
assign lka = ~LKA; //complement 
assign lkm =  KKA & kkb & kkc  |  kka & KKB & kkc  |  kka & kkb & KKC  |  kka & kkb & kkc  ; 
assign LKM = ~lkm;  //complement 
assign EUX =  CDW & DDX  ; 
assign eux = ~EUX;  //complement 
assign EUY =  CDV & DDY  ; 
assign euy = ~EUY;  //complement 
assign EUZ =  CDU & DDZ  ; 
assign euz = ~EUZ;  //complement 
assign ccb = ~CCB;  //complement 
assign cdb = ~CDB;  //complement 
assign frc = ~FRC;  //complement 
assign FRO = ~fro;  //complement 
assign ERX =  CDT & DDX  ; 
assign erx = ~ERX;  //complement 
assign ERY =  CDS & DDY  ; 
assign ery = ~ERY;  //complement 
assign ERZ =  CDR & DDZ  ; 
assign erz = ~ERZ;  //complement 
assign trd = ~TRD;  //complement 
assign dbp = ~DBP;  //complement 
assign dcp = ~DCP;  //complement 
assign ddp = ~DDP;  //complement 
assign dfp = ~DFP;  //complement 
assign DGP = ~dgp;  //complement 
assign DHP = ~dhp;  //complement 
assign daq = ~DAQ;  //complement 
assign dcq = ~DCQ;  //complement 
assign ddq = ~DDQ;  //complement 
assign deq = ~DEQ;  //complement 
assign DGQ = ~dgq;  //complement 
assign DHQ = ~dhq;  //complement 
assign iaa = ~IAA; //complement 
assign iab = ~IAB; //complement 
assign iac = ~IAC; //complement 
assign iad = ~IAD; //complement 
assign iae = ~IAE; //complement 
assign iaf = ~IAF; //complement 
assign iag = ~IAG; //complement 
assign iah = ~IAH; //complement 
assign iai = ~IAI; //complement 
assign iaj = ~IAJ; //complement 
assign iak = ~IAK; //complement 
assign ial = ~IAL; //complement 
assign iam = ~IAM; //complement 
assign ian = ~IAN; //complement 
assign iao = ~IAO; //complement 
assign iap = ~IAP; //complement 
assign iaq = ~IAQ; //complement 
assign iar = ~IAR; //complement 
assign ias = ~IAS; //complement 
assign iat = ~IAT; //complement 
assign iau = ~IAU; //complement 
assign iav = ~IAV; //complement 
assign iaw = ~IAW; //complement 
assign iax = ~IAX; //complement 
assign iay = ~IAY; //complement 
assign iaz = ~IAZ; //complement 
assign iba = ~IBA; //complement 
assign ibb = ~IBB; //complement 
assign ibc = ~IBC; //complement 
assign ibd = ~IBD; //complement 
assign ibe = ~IBE; //complement 
assign ibf = ~IBF; //complement 
assign ibg = ~IBG; //complement 
assign ibh = ~IBH; //complement 
assign ibi = ~IBI; //complement 
assign ibj = ~IBJ; //complement 
assign ibk = ~IBK; //complement 
assign ibl = ~IBL; //complement 
assign ibm = ~IBM; //complement 
assign ibn = ~IBN; //complement 
assign ibo = ~IBO; //complement 
assign ibp = ~IBP; //complement 
assign ibq = ~IBQ; //complement 
assign ibr = ~IBR; //complement 
assign ibs = ~IBS; //complement 
assign ibt = ~IBT; //complement 
assign ibu = ~IBU; //complement 
assign ibv = ~IBV; //complement 
assign ibw = ~IBW; //complement 
assign ibx = ~IBX; //complement 
assign iby = ~IBY; //complement 
assign ibz = ~IBZ; //complement 
assign ica = ~ICA; //complement 
assign icb = ~ICB; //complement 
assign icc = ~ICC; //complement 
assign icd = ~ICD; //complement 
assign ice = ~ICE; //complement 
assign icf = ~ICF; //complement 
assign icg = ~ICG; //complement 
assign ich = ~ICH; //complement 
assign ici = ~ICI; //complement 
assign icj = ~ICJ; //complement 
assign iia = ~IIA; //complement 
assign ika = ~IKA; //complement 
assign ikb = ~IKB; //complement 
assign ikc = ~IKC; //complement 
assign ikd = ~IKD; //complement 
assign ike = ~IKE; //complement 
assign ikf = ~IKF; //complement 
assign ikg = ~IKG; //complement 
assign ikh = ~IKH; //complement 
assign iki = ~IKI; //complement 
assign ikj = ~IKJ; //complement 
assign ikk = ~IKK; //complement 
assign ikl = ~IKL; //complement 
assign ikm = ~IKM; //complement 
assign ila = ~ILA; //complement 
assign ilb = ~ILB; //complement 
assign ilc = ~ILC; //complement 
assign ild = ~ILD; //complement 
assign ile = ~ILE; //complement 
assign ilf = ~ILF; //complement 
assign ilg = ~ILG; //complement 
assign ilh = ~ILH; //complement 
assign ili = ~ILI; //complement 
assign ima = ~IMA; //complement 
assign imb = ~IMB; //complement 
assign imc = ~IMC; //complement 
assign imd = ~IMD; //complement 
assign ime = ~IME; //complement 
assign imf = ~IMF; //complement 
assign img = ~IMG; //complement 
assign imh = ~IMH; //complement 
assign ina = ~INA; //complement 
assign inb = ~INB; //complement 
assign inc = ~INC; //complement 
assign ind = ~IND; //complement 
assign ioa = ~IOA; //complement 
assign iob = ~IOB; //complement 
assign ira = ~IRA; //complement 
assign isa = ~ISA; //complement 
assign isb = ~ISB; //complement 
assign isc = ~ISC; //complement 
assign ita = ~ITA; //complement 
always@(posedge IZZ )
   begin 
 FAA <=  EAA & eab & eac  |  eaa & EAB & eac  |  eaa & eab & EAC  |  EAA & EAB & EAC  ;
 fam <=  EAA & eab & eac  |  eaa & EAB & eac  |  eaa & eab & EAC  |  eaa & eab & eac  ;
 FDA <=  EDY & edz & qad  |  edy & EDZ & qad  |  edy & edz & QAD  |  EDY & EDZ & QAD  ;
 fdm <=  EDY & edz & qad  |  edy & EDZ & qad  |  edy & edz & QAD  |  edy & edz & qad  ;
 FEA <=  EEE & eef & eeg  |  eee & EEF & eeg  |  eee & eef & EEG  |  EEE & EEF & EEG  ;
 fem <=  EEE & eef & eeg  |  eee & EEF & eeg  |  eee & eef & EEG  |  eee & eef & eeg  ;
 FIA <=  EII & eij & eik  |  eii & EIJ & eik  |  eii & eij & EIK  |  EII & EIJ & EIK  ;
 fim <=  EII & eij & eik  |  eii & EIJ & eik  |  eii & eij & EIK  |  eii & eij & eik  ;
 FBA <=  EBE & ebf & ebg  |  ebe & EBF & ebg  |  ebe & ebf & EBG  |  EBE & EBF & EBG  ;
 fbm <=  EBE & ebf & ebg  |  ebe & EBF & ebg  |  ebe & ebf & EBG  |  ebe & ebf & ebg  ;
 FCA <=  ECU & ecv & ecw  |  ecu & ECV & ecw  |  ecu & ecv & ECW  |  ECU & ECV & ECW  ;
 fcm <=  ECU & ecv & ecw  |  ecu & ECV & ecw  |  ecu & ecv & ECW  |  ecu & ecv & ecw  ;
 FFA <=  EFI & efj & efk  |  efi & EFJ & efk  |  efi & efj & EFK  |  EFI & EFJ & EFK  ;
 ffm <=  EFI & efj & efk  |  efi & EFJ & efk  |  efi & efj & EFK  |  efi & efj & efk  ;
 FGA <=  EGY & egz & qag  |  egy & EGZ & qag  |  egy & egz & QAG  |  EGY & EGZ & QAG  ;
 fgm <=  EGY & egz & qag  |  egy & EGZ & qag  |  egy & egz & QAG  |  egy & egz & qag  ;
 FBB <=  EBQ & ebr & ebs  |  ebq & EBR & ebs  |  ebq & ebr & EBS  |  EBQ & EBR & EBS  ;
 fbn <=  EBQ & ebr & ebs  |  ebq & EBR & ebs  |  ebq & ebr & EBS  |  ebq & ebr & ebs  ;
 FCB <=  ECI & ecj & eck  |  eci & ECJ & eck  |  eci & ecj & ECK  |  ECI & ECJ & ECK  ;
 fcn <=  ECI & ecj & eck  |  eci & ECJ & eck  |  eci & ecj & ECK  |  eci & ecj & eck  ;
 FFB <=  EFU & efv & efw  |  efu & EFV & efw  |  efu & efv & EFW  |  EFU & EFV & EFW  ;
 ffn <=  EFU & efv & efw  |  efu & EFV & efw  |  efu & efv & EFW  |  efu & efv & efw  ;
 FGB <=  EGM & egn & ego  |  egm & EGN & ego  |  egm & egn & EGO  |  EGM & EGN & EGO  ;
 fgn <=  EGM & egn & ego  |  egm & EGN & ego  |  egm & egn & EGO  |  egm & egn & ego  ;
 FAB <=  EAM & ean & eao  |  eam & EAN & eao  |  eam & ean & EAO  |  EAM & EAN & EAO  ;
 fan <=  EAM & ean & eao  |  eam & EAN & eao  |  eam & ean & EAO  |  eam & ean & eao  ;
 FDB <=  EDM & edn & edo  |  edm & EDN & edo  |  edm & edn & EDO  |  EDM & EDN & EDO  ;
 fdn <=  EDM & edn & edo  |  edm & EDN & edo  |  edm & edn & EDO  |  edm & edn & edo  ;
 FEB <=  EEQ & eer & ees  |  eeq & EER & ees  |  eeq & eer & EES  |  EEQ & EER & EES  ;
 fen <=  EEQ & eer & ees  |  eeq & EER & ees  |  eeq & eer & EES  |  eeq & eer & ees  ;
 FHA <=  EHQ & ehr & ehs  |  ehq & EHR & ehs  |  ehq & ehr & EHS  |  EHQ & EHR & EHS  ;
 fhm <=  EHQ & ehr & ehs  |  ehq & EHR & ehs  |  ehq & ehr & EHS  |  ehq & ehr & ehs  ;
 FMA <=  EMM & emn & emo  |  emm & EMN & emo  |  emm & emn & EMO  |  EMM & EMN & EMO  ;
 fmm <=  EMM & emn & emo  |  emm & EMN & emo  |  emm & emn & EMO  |  emm & emn & emo  ;
 FQA <=  EQQ & eqr & eqs  |  eqq & EQR & eqs  |  eqq & eqr & EQS  |  EQQ & EQR & EQS  ;
 fqm <=  EQQ & eqr & eqs  |  eqq & EQR & eqs  |  eqq & eqr & EQS  |  eqq & eqr & eqs  ;
 FUA <=  EUU & euv & euw  |  euu & EUV & euw  |  euu & euv & EUW  |  EUU & EUV & EUW  ;
 fum <=  EUU & euv & euw  |  euu & EUV & euw  |  euu & euv & EUW  |  euu & euv & euw  ;
 FJA <=  EJM & ejn & ejo  |  ejm & EJN & ejo  |  ejm & ejn & EJO  |  EJM & EJN & EJO  ;
 fjm <=  EJM & ejn & ejo  |  ejm & EJN & ejo  |  ejm & ejn & EJO  |  ejm & ejn & ejo  ;
 FNA <=  ENQ & enr & ens  |  enq & ENR & ens  |  enq & enr & ENS  |  ENQ & ENR & ENS  ;
 fnm <=  ENQ & enr & ens  |  enq & ENR & ens  |  enq & enr & ENS  |  enq & enr & ens  ;
 FRA <=  ERU & erv & erw  |  eru & ERV & erw  |  eru & erv & ERW  |  ERU & ERV & ERW  ;
 frm <=  ERU & erv & erw  |  eru & ERV & erw  |  eru & erv & ERW  |  eru & erv & erw  ;
 FJB <=  EJY & ejz & qaj  |  ejy & EJZ & qaj  |  ejy & ejz & QAJ  |  EJY & EJZ & QAJ  ;
 fjn <=  EJY & ejz & qaj  |  ejy & EJZ & qaj  |  ejy & ejz & QAJ  |  ejy & ejz & qaj  ;
 FKA <=  EKQ & ekr & eks  |  ekq & EKR & eks  |  ekq & ekr & EKS  |  EKQ & EKR & EKS  ;
 fkm <=  EKQ & ekr & eks  |  ekq & EKR & eks  |  ekq & ekr & EKS  |  ekq & ekr & eks  ;
 FOA <=  EOU & eov & eow  |  eou & EOV & eow  |  eou & eov & EOW  |  EOU & EOV & EOW  ;
 fom <=  EOU & eov & eow  |  eou & EOV & eow  |  eou & eov & EOW  |  eou & eov & eow  ;
 FIB <=  EIU & eiv & eiw  |  eiu & EIV & eiw  |  eiu & eiv & EIW  |  EIU & EIV & EIW  ;
 fin <=  EIU & eiv & eiw  |  eiu & EIV & eiw  |  eiu & eiv & EIW  |  eiu & eiv & eiw  ;
 FLA <=  ELU & elv & elw  |  elu & ELV & elw  |  elu & elv & ELW  |  ELU & ELV & ELW  ;
 flm <=  ELU & elv & elw  |  elu & ELV & elw  |  elu & elv & ELW  |  elu & elv & elw  ;
 FMB <=  EMY & emz & qam  |  emy & EMZ & qam  |  emy & emz & QAM  |  EMY & EMZ & QAM  ;
 fmn <=  EMY & emz & qam  |  emy & EMZ & qam  |  emy & emz & QAM  |  emy & emz & qam  ;
 DAA <= IBA ; 
 DAB <= IBB ; 
 DBB <= IBB ; 
 FYA <=  EYY & eyz & qay  |  eyy & EYZ & qay  |  eyy & eyz & QAY  |  EYY & EYZ & QAY  ;
 fym <=  EYY & eyz & qay  |  eyy & EYZ & qay  |  eyy & eyz & QAY  |  eyy & eyz & qay  ;
 FVA <=  EVY & evz & qav  |  evy & EVZ & qav  |  evy & evz & QAV  |  EVY & EVZ & QAV  ;
 fvm <=  EVY & evz & qav  |  evy & EVZ & qav  |  evy & evz & QAV  |  evy & evz & qav  ;
 QRA <= IRA ; 
 FSA <=  ESY & esz & qas  |  esy & ESZ & qas  |  esy & esz & QAS  |  ESY & ESZ & QAS  ;
 fsm <=  ESY & esz & qas  |  esy & ESZ & qas  |  esy & esz & QAS  |  esy & esz & qas  ;
 TRA <= QRA ; 
 FPA <=  EPY & epz & qap  |  epy & EPZ & qap  |  epy & epz & QAP  |  EPY & EPZ & QAP  ;
 fpm <=  EPY & epz & qap  |  epy & EPZ & qap  |  epy & epz & QAP  |  epy & epz & qap  ;
 FAC <=  EAV & eaw & eax  |  eav & EAW & eax  |  eav & eaw & EAX  |  EAV & EAW & EAX  ;
 fao <=  EAV & eaw & eax  |  eav & EAW & eax  |  eav & eaw & EAX  |  eav & eaw & eax  ;
 FBC <=  EBB & ebc & ebd  |  ebb & EBC & ebd  |  ebb & ebc & EBD  |  EBB & EBC & EBD  ;
 fbo <=  EBB & ebc & ebd  |  ebb & EBC & ebd  |  ebb & ebc & EBD  |  ebb & ebc & ebd  ;
 FFC <=  EFF & efg & efh  |  eff & EFG & efh  |  eff & efg & EFH  |  EFF & EFG & EFH  ;
 ffo <=  EFF & efg & efh  |  eff & EFG & efh  |  eff & efg & EFH  |  eff & efg & efh  ;
 FCC <=  ECF & ecg & ech  |  ecf & ECG & ech  |  ecf & ecg & ECH  |  ECF & ECG & ECH  ;
 fco <=  ECF & ecg & ech  |  ecf & ECG & ech  |  ecf & ecg & ECH  |  ecf & ecg & ech  ;
 FDC <=  EDV & edw & edx  |  edv & EDW & edx  |  edv & edw & EDX  |  EDV & EDW & EDX  ;
 fdo <=  EDV & edw & edx  |  edv & EDW & edx  |  edv & edw & EDX  |  edv & edw & edx  ;
 FGC <=  EGJ & egk & egl  |  egj & EGK & egl  |  egj & egk & EGL  |  EGJ & EGK & EGL  ;
 fgo <=  EGJ & egk & egl  |  egj & EGK & egl  |  egj & egk & EGL  |  egj & egk & egl  ;
 FEH <= EEZ ; 
 FEC <=  EEN & eeo & eep  |  een & EEO & eep  |  een & eeo & EEP  |  EEN & EEO & EEP  ;
 feo <=  EEN & eeo & eep  |  een & EEO & eep  |  een & eeo & EEP  |  een & eeo & eep  ;
 FCD <=  ECR & ecs & ect  |  ecr & ECS & ect  |  ecr & ecs & ECT  |  ECR & ECS & ECT  ;
 fcp <=  ECR & ecs & ect  |  ecr & ECS & ect  |  ecr & ecs & ECT  |  ecr & ecs & ect  ;
 FDD <=  EDJ & edk & edl  |  edj & EDK & edl  |  edj & edk & EDL  |  EDJ & EDK & EDL  ;
 fdp <=  EDJ & edk & edl  |  edj & EDK & edl  |  edj & edk & EDL  |  edj & edk & edl  ;
 FGD <=  EGV & egw & egx  |  egv & EGW & egx  |  egv & egw & EGX  |  EGV & EGW & EGX  ;
 fgp <=  EGV & egw & egx  |  egv & EGW & egx  |  egv & egw & EGX  |  egv & egw & egx  ;
 FHB <=  EHN & eho & ehp  |  ehn & EHO & ehp  |  ehn & eho & EHP  |  EHN & EHO & EHP  ;
 fhn <=  EHN & eho & ehp  |  ehn & EHO & ehp  |  ehn & eho & EHP  |  ehn & eho & ehp  ;
 FHG <= EHZ ; 
 FAD <=  EAJ & eak & eal  |  eaj & EAK & eal  |  eaj & eak & EAL  |  EAJ & EAK & EAL  ;
 fap <=  EAJ & eak & eal  |  eaj & EAK & eal  |  eaj & eak & EAL  |  eaj & eak & eal  ;
 FBD <=  EBN & ebo & ebp  |  ebn & EBO & ebp  |  ebn & ebo & EBP  |  EBN & EBO & EBP  ;
 fbp <=  EBN & ebo & ebp  |  ebn & EBO & ebp  |  ebn & ebo & EBP  |  ebn & ebo & ebp  ;
 FFD <=  EFR & efs & eft  |  efr & EFS & eft  |  efr & efs & EFT  |  EFR & EFS & EFT  ;
 ffp <=  EFR & efs & eft  |  efr & EFS & eft  |  efr & efs & EFT  |  efr & efs & eft  ;
 FJC <=  EJJ & ejk & ejl  |  ejj & EJK & ejl  |  ejj & ejk & EJL  |  EJJ & EJK & EJL  ;
 fjo <=  EJJ & ejk & ejl  |  ejj & EJK & ejl  |  ejj & ejk & EJL  |  ejj & ejk & ejl  ;
 FNB <=  ENN & eno & enp  |  enn & ENO & enp  |  enn & eno & ENP  |  ENN & ENO & ENP  ;
 fnn <=  ENN & eno & enp  |  enn & ENO & enp  |  enn & eno & ENP  |  enn & eno & enp  ;
 FRB <=  ERR & ers & ert  |  err & ERS & ert  |  err & ers & ERT  |  ERR & ERS & ERT  ;
 frn <=  ERR & ers & ert  |  err & ERS & ert  |  err & ers & ERT  |  err & ers & ert  ;
 FWC <= QAW ; 
 FKB <=  EKN & eko & ekp  |  ekn & EKO & ekp  |  ekn & eko & EKP  |  EKN & EKO & EKP  ;
 fkn <=  EKN & eko & ekp  |  ekn & EKO & ekp  |  ekn & eko & EKP  |  ekn & eko & ekp  ;
 FKF <= EKZ ; 
 FJD <=  EJV & ejw & ejx  |  ejv & EJW & ejx  |  ejv & ejw & EJX  |  EJV & EJW & EJX  ;
 fjp <=  EJV & ejw & ejx  |  ejv & EJW & ejx  |  ejv & ejw & EJX  |  ejv & ejw & ejx  ;
 FOB <=  EOR & eos & eot  |  eor & EOS & eot  |  eor & eos & EOT  |  EOR & EOS & EOT  ;
 fon <=  EOR & eos & eot  |  eor & EOS & eot  |  eor & eos & EOT  |  eor & eos & eot  ;
 FSB <=  ESV & esw & esx  |  esv & ESW & esx  |  esv & esw & ESX  |  ESV & ESW & ESX  ;
 fsn <=  ESV & esw & esx  |  esv & ESW & esx  |  esv & esw & ESX  |  esv & esw & esx  ;
 FTD <= QAT ; 
 FLB <=  ELR & els & elt  |  elr & ELS & elt  |  elr & els & ELT  |  ELR & ELS & ELT  ;
 fln <=  ELR & els & elt  |  elr & ELS & elt  |  elr & els & ELT  |  elr & els & elt  ;
 FPB <=  EPV & epw & epx  |  epv & EPW & epx  |  epv & epw & EPX  |  EPV & EPW & EPX  ;
 fpn <=  EPV & epw & epx  |  epv & EPW & epx  |  epv & epw & EPX  |  epv & epw & epx  ;
 FQE <= QAQ ; 
 FIC <=  EIR & eis & eit  |  eir & EIS & eit  |  eir & eis & EIT  |  EIR & EIS & EIT  ;
 fio <=  EIR & eis & eit  |  eir & EIS & eit  |  eir & eis & EIT  |  eir & eis & eit  ;
 FMC <=  EMV & emw & emx  |  emv & EMW & emx  |  emv & emw & EMX  |  EMV & EMW & EMX  ;
 fmo <=  EMV & emw & emx  |  emv & EMW & emx  |  emv & emw & EMX  |  emv & emw & emx  ;
 FNF <= QAN ; 
 FVB <=  EVV & evw & evx  |  evv & EVW & evx  |  evv & evw & EVX  |  EVV & EVW & EVX  ;
 fvn <=  EVV & evw & evx  |  evv & EVW & evx  |  evv & evw & EVX  |  evv & evw & evx  ;
 DAF <= IBF ; 
 DBF <= IBF ; 
 DDF <= IBF ; 
 DAJ <= IBJ ; 
 DBJ <= IBJ ; 
 DDJ <= IBJ ; 
 DFJ <= IBJ ; 
 DAG <= IBG ; 
 DBG <= IBG ; 
 DCG <= IBG ; 
 DDR <= IBR ; 
 DDV <= IBV ; 
 dgk <= ibk ; 
 DAK <= IBK ; 
 DBK <= IBK ; 
 DCK <= IBK ; 
 DFK <= IBK ; 
 cdf <= iaf & TRB |  icf & trb ; 
 cdg <= iag & TRB |  icg & trb ; 
 DAO <= IBO ; 
 DBO <= IBO ; 
 DCO <= IBO ; 
 DEO <= IBO ; 
 CAG <=  IAG & TRB  |  ICG & trb  ; 
 CBG <=  IAG & TRB  |  ICG & trb  ; 
 CCG <=  IAG & TRB  |  ICG & trb  ; 
 CAF <=  IAF & TRB  |  ICF & trb  ; 
 CBF <=  IAF & TRB  |  ICF & trb  ; 
 CCF <=  IAF & TRB  |  ICF & trb  ; 
 FTC <= ETZ ; 
 FUC <= QAU ; 
 FWB <= EWZ ; 
 dfn <= ibn ; 
 dfo <= ibo ; 
 dgo <= ibo ; 
 dhn <= ibn ; 
 cdi <= iai & TRB |  ici & trb ; 
 CAI <=  IAI & TRB  |  ICI & trb  ; 
 CBI <=  IAI & TRB  |  ICI & trb  ; 
 CCI <=  IAI & TRB  |  ICI & trb  ; 
 dfv <= ibv ; 
 dfw <= ibw ; 
 dgw <= ibw ; 
 dhv <= ibv ; 
 DAN <= IBN ; 
 DBN <= IBN ; 
 DDN <= IBN ; 
 DEN <= IBN ; 
 TRB <= QRA ; 
 FQD <= EQZ ; 
 DAW <= IBW ; 
 DBW <= IBW ; 
 DCW <= IBW ; 
 DEW <= IBW ; 
 DAV <= IBV ; 
 DBV <= IBV ; 
 DEV <= IBV ; 
 dfr <= ibr ; 
 dfs <= ibs ; 
 dgs <= ibs ; 
 dhr <= ibr ; 
 DAR <= IBR ; 
 DBR <= IBR ; 
 DER <= IBR ; 
 DAS <= IBS ; 
 DBS <= IBS ; 
 DCS <= IBS ; 
 DES <= IBS ; 
 HAA <=  GAA & ilf & ila  |  gaa & ILF & ila  |  gaa & ilf & ILA  |  GAA & ILF & ILA  ;
 ham <=  GAA & ilf & ila  |  gaa & ILF & ila  |  gaa & ilf & ILA  |  gaa & ilf & ila  ;
 HEA <=  GEA & gdn & gdm  |  gea & GDN & gdm  |  gea & gdn & GDM  |  GEA & GDN & GDM  ;
 hem <=  GEA & gdn & gdm  |  gea & GDN & gdm  |  gea & gdn & GDM  |  gea & gdn & gdm  ;
 HGD <= GFM ; 
 HBA <=  GBA & gam & gbb  |  gba & GAM & gbb  |  gba & gam & GBB  |  GBA & GAM & GBB  ;
 hbm <=  GBA & gam & gbb  |  gba & GAM & gbb  |  gba & gam & GBB  |  gba & gam & gbb  ;
 HHA <=  GGM & gha & ggn  |  ggm & GHA & ggn  |  ggm & gha & GGN  |  GGM & GHA & GGN  ;
 hhm <=  GGM & gha & ggn  |  ggm & GHA & ggn  |  ggm & gha & GGN  |  ggm & gha & ggn  ;
 HAD <=  GAC & ili & ile  |  gac & ILI & ile  |  gac & ili & ILE  |  GAC & ILI & ILE  ;
 hap <=  GAC & ili & ile  |  gac & ILI & ile  |  gac & ili & ILE  |  gac & ili & ile  ;
 HED <=  GEE & gdq & fdt  |  gee & GDQ & fdt  |  gee & gdq & FDT  |  GEE & GDQ & FDT  ;
 hep <=  GEE & gdq & fdt  |  gee & GDQ & fdt  |  gee & gdq & FDT  |  gee & gdq & fdt  ;
 HFA <=  GEM & gen & gfb  |  gem & GEN & gfb  |  gem & gen & GFB  |  GEM & GEN & GFB  ;
 hfm <=  GEM & gen & gfb  |  gem & GEN & gfb  |  gem & gen & GFB  |  gem & gen & gfb  ;
 HFD <= GFA ; 
 HAC <=  GAB & ild & ilh  |  gab & ILD & ilh  |  gab & ild & ILH  |  GAB & ILD & ILH  ;
 hao <=  GAB & ild & ilh  |  gab & ILD & ilh  |  gab & ild & ILH  |  gab & ild & ilh  ;
 HCB <=  GCC & fcd & gcb  |  gcc & FCD & gcb  |  gcc & fcd & GCB  |  GCC & FCD & GCB  ;
 hcn <=  GCC & fcd & gcb  |  gcc & FCD & gcb  |  gcc & fcd & GCB  |  gcc & fcd & gcb  ;
 HDE <= GDB ; 
 HEC <=  GED & fdp & gdp  |  ged & FDP & gdp  |  ged & fdp & GDP  |  GED & FDP & GDP  ;
 heo <=  GED & fdp & gdp  |  ged & FDP & gdp  |  ged & fdp & GDP  |  ged & fdp & gdp  ;
 HGA <=  GFN & ggb & fgd  |  gfn & GGB & fgd  |  gfn & ggb & FGD  |  GFN & GGB & FGD  ;
 hgm <=  GFN & ggb & fgd  |  gfn & GGB & fgd  |  gfn & ggb & FGD  |  gfn & ggb & fgd  ;
 HDB <=  GCO & gdd & gcp  |  gco & GDD & gcp  |  gco & gdd & GCP  |  GCO & GDD & GCP  ;
 hdn <=  GCO & gdd & gcp  |  gco & GDD & gcp  |  gco & gdd & GCP  |  gco & gdd & gcp  ;
 HBC <=  GBF & gao & gbe  |  gbf & GAO & gbe  |  gbf & gao & GBE  |  GBF & GAO & GBE  ;
 hbo <=  GBF & gao & gbe  |  gbf & GAO & gbe  |  gbf & gao & GBE  |  gbf & gao & gbe  ;
 HFC <=  GFE & geq & gfd  |  gfe & GEQ & gfd  |  gfe & geq & GFD  |  GFE & GEQ & GFD  ;
 hfo <=  GFE & geq & gfd  |  gfe & GEQ & gfd  |  gfe & geq & GFD  |  gfe & geq & gfd  ;
 HKA <=  GKA & gjm & gjn  |  gka & GJM & gjn  |  gka & gjm & GJN  |  GKA & GJM & GJN  ;
 hkm <=  GKA & gjm & gjn  |  gka & GJM & gjn  |  gka & gjm & GJN  |  gka & gjm & gjn  ;
 FXB <= QAX ; 
 HJA <=  GJA & gjb & gim  |  gja & GJB & gim  |  gja & gjb & GIM  |  GJA & GJB & GIM  ;
 hjm <=  GJA & gjb & gim  |  gja & GJB & gim  |  gja & gjb & GIM  |  gja & gjb & gim  ;
 HOA <=  GOA & gnm & gnn  |  goa & GNM & gnn  |  goa & gnm & GNN  |  GOA & GNM & GNN  ;
 hom <=  GOA & gnm & gnn  |  goa & GNM & gnn  |  goa & gnm & GNN  |  goa & gnm & gnn  ;
 HQB <= GPM ; 
 HPA <=  FPD & gom & foo  |  fpd & GOM & foo  |  fpd & gom & FOO  |  FPD & GOM & FOO  ;
 hpm <=  FPD & gom & foo  |  fpd & GOM & foo  |  fpd & gom & FOO  |  fpd & gom & foo  ;
 HRA <=  GRA & gqm & fra  |  gra & GQM & fra  |  gra & gqm & FRA  |  GRA & GQM & FRA  ;
 hrm <=  GRA & gqm & fra  |  gra & GQM & fra  |  gra & gqm & FRA  |  gra & gqm & fra  ;
 HLB <=  GKN & glb & fkm  |  gkn & GLB & fkm  |  gkn & glb & FKM  |  GKN & GLB & FKM  ;
 hln <=  GKN & glb & fkm  |  gkn & GLB & fkm  |  gkn & glb & FKM  |  gkn & glb & fkm  ;
 HGB <=  GGC & gfp & gfo  |  ggc & GFP & gfo  |  ggc & gfp & GFO  |  GGC & GFP & GFO  ;
 hgn <=  GGC & gfp & gfo  |  ggc & GFP & gfo  |  ggc & gfp & GFO  |  ggc & gfp & gfo  ;
 HID <= GHQ ; 
 HKC <=  GJO & gkd & gjp  |  gjo & GKD & gjp  |  gjo & gkd & GJP  |  GJO & GKD & GJP  ;
 hko <=  GJO & gkd & gjp  |  gjo & GKD & gjp  |  gjo & gkd & GJP  |  gjo & gkd & gjp  ;
 HNB <=  GMN & gnc & gmo  |  gmn & GNC & gmo  |  gmn & gnc & GMO  |  GMN & GNC & GMO  ;
 hnn <=  GMN & gnc & gmo  |  gmn & GNC & gmo  |  gmn & gnc & GMO  |  gmn & gnc & gmo  ;
 HWA <=  GWA & gvm & fvm  |  gwa & GVM & fvm  |  gwa & gvm & FVM  |  GWA & GVM & FVM  ;
 hwm <=  GWA & gvm & fvm  |  gwa & GVM & fvm  |  gwa & gvm & FVM  |  gwa & gvm & fvm  ;
 QAW <=  IKI & TTB  |  IKJ & ttb  |  QIB  ; 
 DAC <= IBC ; 
 DBC <= IBC ; 
 DCC <= IBC ; 
 HVA <=  GVA & gum & fva  |  gva & GUM & fva  |  gva & gum & FVA  |  GVA & GUM & FVA  ;
 hvm <=  GVA & gum & fva  |  gva & GUM & fva  |  gva & gum & FVA  |  gva & gum & fva  ;
 QAY <=  IKK & TTB  |  IKL & ttb  |  QIB  ; 
 CAD <=  IAD & TRE  |  ICD & tre  ; 
 CBD <=  IAD & TRE  |  ICD & tre  ; 
 CCD <=  IAD & TRE  |  ICD & tre  ; 
 HSA <=  GSA & grm & gsb  |  gsa & GRM & gsb  |  gsa & grm & GSB  |  GSA & GRM & GSB  ;
 hsm <=  GSA & grm & gsb  |  gsa & GRM & gsb  |  gsa & grm & GSB  |  gsa & grm & gsb  ;
 HTB <= GSM ; 
 qaj <= qie ; 
 qam <= qie ; 
 QBC <= QBB ; 
 QBE <= QBD ; 
 qad <= qic ; 
 qag <= qic ; 
 OZN <= QBE ; 
 QBB <= QBA ; 
 QBD <= QBC ; 
 HTA <=  FSM & gtb & gsn  |  fsm & GTB & gsn  |  fsm & gtb & GSN  |  FSM & GTB & GSN  ;
 htm <=  FSM & gtb & gsn  |  fsm & GTB & gsn  |  fsm & gtb & GSN  |  fsm & gtb & gsn  ;
 QAT <=  IKF & TTB  |  IKG & ttb  |  QIC  ; 
 QAV <=  IKH & TTB  |  IKI & ttb  |  QIC  ; 
 cdd <= iad & TRE |  icd & tre ; 
 HPB <=  GON & gpb & goo  |  gon & GPB & goo  |  gon & gpb & GOO  |  GON & GPB & GOO  ;
 hpn <=  GON & gpb & goo  |  gon & GPB & goo  |  gon & gpb & GOO  |  gon & gpb & goo  ;
 HWB <= FWB ; 
 QBA <=  IKM & TTB  |  QIB  ; 
 HOB <=  GOB & gno & goc  |  gob & GNO & goc  |  gob & gno & GOC  |  GOB & GNO & GOC  ;
 hon <=  GOB & gno & goc  |  gob & GNO & goc  |  gob & gno & GOC  |  gob & gno & goc  ;
 TRF <= QRA ; 
 QAQ <=  IKC & TTA  |  IKD & tta  |  QID  ; 
 QAS <=  IKE & TTA  |  IKF & tta  |  QID  ; 
 TRE <= QRA ; 
 HQA <=  GQB & gpn & gqc  |  gqb & GPN & gqc  |  gqb & gpn & GQC  |  GQB & GPN & GQC  ;
 hqm <=  GQB & gpn & gqc  |  gqb & GPN & gqc  |  gqb & gpn & GQC  |  gqb & gpn & gqc  ;
 CAQ <= IAQ ; 
 CBQ <= IAQ ; 
 CCQ <= IAQ ; 
 CDQ <= IAQ ; 
 QAN <=  ZZI & TTA  |  IKA & tta  |  QIE  ; 
 QAP <=  IKB & TTA  |  IKC & tta  |  QIE  ; 
 CAP <= IAP ; 
 CBP <= IAP ; 
 CCP <= IAP ; 
 CDP <= IAP ; 
 KFA <=  JFA & jem & hem  |  jfa & JEM & hem  |  jfa & jem & HEM  |  JFA & JEM & HEM  ;
 kfm <=  JFA & jem & hem  |  jfa & JEM & hem  |  jfa & jem & HEM  |  jfa & jem & hem  ;
 MAB <= INA ; 
 MGA <=  LGA & lfm & kfn  |  lga & LFM & kfn  |  lga & lfm & KFN  |  LGA & LFM & KFN  ;
 mgm <=  LGA & lfm & kfn  |  lga & LFM & kfn  |  lga & lfm & KFN  |  lga & lfm & kfn  ;
 KGA <=  JFM & hfm & hgd  |  jfm & HFM & hgd  |  jfm & hfm & HGD  |  JFM & HFM & HGD  ;
 kgm <=  JFM & hfm & hgd  |  jfm & HFM & hgd  |  jfm & hfm & HGD  |  jfm & hfm & hgd  ;
 KIB <= HHM ; 
 KEB <=  JDO & jeb & hdo  |  jdo & JEB & hdo  |  jdo & jeb & HDO  |  JDO & JEB & HDO  ;
 ken <=  JDO & jeb & hdo  |  jdo & JEB & hdo  |  jdo & jeb & HDO  |  jdo & jeb & hdo  ;
 MBC <= IND ; 
 MBA <=  KBA & kam & lam  |  kba & KAM & lam  |  kba & kam & LAM  |  KBA & KAM & LAM  ;
 mbm <=  KBA & kam & lam  |  kba & KAM & lam  |  kba & kam & LAM  |  kba & kam & lam  ;
 MBB <= LBA ; 
 MFA <=  LFA & kfb & lem  |  lfa & KFB & lem  |  lfa & kfb & LEM  |  LFA & KFB & LEM  ;
 mfm <=  LFA & kfb & lem  |  lfa & KFB & lem  |  lfa & kfb & LEM  |  lfa & kfb & lem  ;
 KGB <=  JFN & jga & jgb  |  jfn & JGA & jgb  |  jfn & jga & JGB  |  JFN & JGA & JGB  ;
 kgn <=  JFN & jga & jgb  |  jfn & JGA & jgb  |  jfn & jga & JGB  |  jfn & jga & jgb  ;
 KHB <= JHA ; 
 KAB <=  HAD & imf & imc  |  had & IMF & imc  |  had & imf & IMC  |  HAD & IMF & IMC  ;
 kan <=  HAD & imf & imc  |  had & IMF & imc  |  had & imf & IMC  |  had & imf & imc  ;
 KAD <= IMD ; 
 KBB <=  HAP & hbc & jbb  |  hap & HBC & jbb  |  hap & hbc & JBB  |  HAP & HBC & JBB  ;
 kbn <=  HAP & hbc & jbb  |  hap & HBC & jbb  |  hap & hbc & JBB  |  hap & hbc & jbb  ;
 KBC <= IMH ; 
 KBA <=  IMG & jba & jam  |  img & JBA & jam  |  img & jba & JAM  |  IMG & JBA & JAM  ;
 kbm <=  IMG & jba & jam  |  img & JBA & jam  |  img & jba & JAM  |  img & jba & jam  ;
 MCA <=  LCA & lbm & kcb  |  lca & LBM & kcb  |  lca & lbm & KCB  |  LCA & LBM & KCB  ;
 mcm <=  LCA & lbm & kcb  |  lca & LBM & kcb  |  lca & lbm & KCB  |  lca & lbm & kcb  ;
 MDB <= LCM ; 
 KFB <=  HFC & jfb & jen  |  hfc & JFB & jen  |  hfc & jfb & JEN  |  HFC & JFB & JEN  ;
 kfn <=  HFC & jfb & jen  |  hfc & JFB & jen  |  hfc & jfb & JEN  |  hfc & jfb & jen  ;
 MHA <=  LGM & kgm & lha  |  lgm & KGM & lha  |  lgm & kgm & LHA  |  LGM & KGM & LHA  ;
 mhm <=  LGM & kgm & lha  |  lgm & KGM & lha  |  lgm & kgm & LHA  |  lgm & kgm & lha  ;
 KIC <= JHM ; 
 KKA <=  JJM & hjm & hka  |  jjm & HJM & hka  |  jjm & hjm & HKA  |  JJM & HJM & HKA  ;
 kkm <=  JJM & hjm & hka  |  jjm & HJM & hka  |  jjm & hjm & HKA  |  jjm & hjm & hka  ;
 MKA <=  LKA & ljm & kjm  |  lka & LJM & kjm  |  lka & ljm & KJM  |  LKA & LJM & KJM  ;
 mkm <=  LKA & ljm & kjm  |  lka & LJM & kjm  |  lka & ljm & KJM  |  lka & ljm & kjm  ;
 MLA <=  KKM & lkm & kla  |  kkm & LKM & kla  |  kkm & lkm & KLA  |  KKM & LKM & KLA  ;
 mlm <=  KKM & lkm & kla  |  kkm & LKM & kla  |  kkm & lkm & KLA  |  kkm & lkm & kla  ;
 KOA <=  JOA & jnm & hoa  |  joa & JNM & hoa  |  joa & jnm & HOA  |  JOA & JNM & HOA  ;
 kom <=  JOA & jnm & hoa  |  joa & JNM & hoa  |  joa & jnm & HOA  |  joa & jnm & hoa  ;
 KPB <= HOM ; 
 KPA <=  JOM & jpa & hpa  |  jom & JPA & hpa  |  jom & jpa & HPA  |  JOM & JPA & HPA  ;
 kpm <=  JOM & jpa & hpa  |  jom & JPA & hpa  |  jom & jpa & HPA  |  jom & jpa & hpa  ;
 KQB <= JQA ; 
 MIA <=  LIA & lhm & khm  |  lia & LHM & khm  |  lia & lhm & KHM  |  LIA & LHM & KHM  ;
 mim <=  LIA & lhm & khm  |  lia & LHM & khm  |  lia & lhm & KHM  |  lia & lhm & khm  ;
 ODA <= NDA ; 
 OEA <= NDM ; 
 CAX <= IAX ; 
 CBX <= IAX ; 
 CCX <= IAX ; 
 CDX <= IAX ; 
 MWB <= KWA ; 
 MXA <= KXA ; 
 MXB <= KXB ; 
 MYB <= KYB ; 
 OWB <= MWB ; 
 OXA <= MXA ; 
 OXB <= MXB ; 
 OYB <= MYB ; 
 KWA <= JWA ; 
 KXA <= JWM ; 
 KXB <= JXA ; 
 KYB <= JXM ; 
 OGB <= MGA ; 
 OHA <= MGM ; 
 OHB <= MHA ; 
 OIA <= MHM ; 
 CAU <= IAU ; 
 CBU <= IAU ; 
 CDU <= IAU ; 
 CAV <= IAV ; 
 CBV <= IAV ; 
 CCV <= IAV ; 
 CDV <= IAV ; 
 KRB <= JRA ; 
 MPB <= LPA ; 
 MQA <= LPM ; 
 MQB <= LQA ; 
 MRA <= LQM ; 
 OFB <= MFA ; 
 OGA <= MFM ; 
 OLA <= MKM ; 
 OLB <= MLA ; 
 QTA <= ITA ; 
 TTA <= QTA ; 
 TTB <= QTA ; 
 OPB <= MPB ; 
 OQA <= MQA ; 
 OQB <= MQB ; 
 ORA <= MRA ; 
 KQA <=  JPM & hpn & hqa  |  jpm & HPN & hqa  |  jpm & hpn & HQA  |  JPM & HPN & HQA  ;
 kqm <=  JPM & hpn & hqa  |  jpm & HPN & hqa  |  jpm & hpn & HQA  |  jpm & hpn & hqa  ;
 OIB <= MIA ; 
 OJA <= MIM ; 
 OKB <= MKA ; 
 OMA <= MLM ; 
 KRA <= JQM ; 
 MRB <= LRA ; 
 MSA <= LRM ; 
 CCU <= IAU ; 
 ORB <= MRB ; 
 OSA <= MSA ; 
 KDA <=  JCN & jdc & jdb  |  jcn & JDC & jdb  |  jcn & jdc & JDB  |  JCN & JDC & JDB  ;
 kdm <=  JCN & jdc & jdb  |  jcn & JDC & jdb  |  jcn & jdc & JDB  |  jcn & jdc & jdb  ;
 KAA <=  IME & ima & jaa  |  ime & IMA & jaa  |  ime & ima & JAA  |  IME & IMA & JAA  ;
 kam <=  IME & ima & jaa  |  ime & IMA & jaa  |  ime & ima & JAA  |  ime & ima & jaa  ;
 KAC <= IMB ; 
 KCA <=  JCA & jbn & jbm  |  jca & JBN & jbm  |  jca & jbn & JBM  |  JCA & JBN & JBM  ;
 kcm <=  JCA & jbn & jbm  |  jca & JBN & jbm  |  jca & jbn & JBM  |  jca & jbn & jbm  ;
 KDC <= JCM ; 
 KEA <=  JEA & jdm & jdn  |  jea & JDM & jdn  |  jea & jdm & JDN  |  JEA & JDM & JDN  ;
 kem <=  JEA & jdm & jdn  |  jea & JDM & jdn  |  jea & jdm & JDN  |  jea & jdm & jdn  ;
 KDB <= JDA ; 
 OBA <=  NAM & nba & mbc  |  nam & NBA & mbc  |  nam & nba & MBC  |  NAM & NBA & MBC  ;
 obm <=  NAM & nba & mbc  |  nam & NBA & mbc  |  nam & nba & MBC  |  nam & nba & mbc  ;
 MAA <=  LAA & kaa & inc  |  laa & KAA & inc  |  laa & kaa & INC  |  LAA & KAA & INC  ;
 mam <=  LAA & kaa & inc  |  laa & KAA & inc  |  laa & kaa & INC  |  laa & kaa & inc  ;
 OAA <=  NAA & ioa & iob  |  naa & IOA & iob  |  naa & ioa & IOB  |  NAA & IOA & IOB  ;
 oam <=  NAA & ioa & iob  |  naa & IOA & iob  |  naa & ioa & IOB  |  naa & ioa & iob  ;
 MAC <= INB ; 
 OCA <=  NBM & mbm & mca  |  nbm & MBM & mca  |  nbm & mbm & MCA  |  NBM & MBM & MCA  ;
 ocm <=  NBM & mbm & mca  |  nbm & MBM & mca  |  nbm & mbm & MCA  |  nbm & mbm & mca  ;
 KHA <=  JGN & jhb & jgm  |  jgn & JHB & jgm  |  jgn & jhb & JGM  |  JGN & JHB & JGM  ;
 khm <=  JGN & jhb & jgm  |  jgn & JHB & jgm  |  jgn & jhb & JGM  |  jgn & jhb & jgm  ;
 MEB <= LDM ; 
 KCB <=  JCB & hcd & hbo  |  jcb & HCD & hbo  |  jcb & hcd & HBO  |  JCB & HCD & HBO  ;
 kcn <=  JCB & hcd & hbo  |  jcb & HCD & hbo  |  jcb & hcd & HBO  |  jcb & hcd & hbo  ;
 MDA <=  KCN & kda & lda  |  kcn & KDA & lda  |  kcn & kda & LDA  |  KCN & KDA & LDA  ;
 mdm <=  KCN & kda & lda  |  kcn & KDA & lda  |  kcn & kda & LDA  |  kcn & kda & lda  ;
 MEA <= LEA ; 
 KMA <=  JMA & jlm & jln  |  jma & JLM & jln  |  jma & jlm & JLN  |  JMA & JLM & JLN  ;
 kmm <=  JMA & jlm & jln  |  jma & JLM & jln  |  jma & jlm & JLN  |  jma & jlm & jln  ;
 KNB <= JMM ; 
 KJA <=  JIM & jja & hjc  |  jim & JJA & hjc  |  jim & jja & HJC  |  JIM & JJA & HJC  ;
 kjm <=  JIM & jja & hjc  |  jim & JJA & hjc  |  jim & jja & HJC  |  jim & jja & hjc  ;
 KJC <= JJB ; 
 KLA <=  JKM & jlb & jla  |  jkm & JLB & jla  |  jkm & jlb & JLA  |  JKM & JLB & JLA  ;
 klm <=  JKM & jlb & jla  |  jkm & JLB & jla  |  jkm & jlb & JLA  |  jkm & jlb & jla  ;
 KMB <= JMB ; 
 KIA <=  JIA & jib & jhn  |  jia & JIB & jhn  |  jia & jib & JHN  |  JIA & JIB & JHN  ;
 kim <=  JIA & jib & jhn  |  jia & JIB & jhn  |  jia & jib & JHN  |  jia & jib & jhn  ;
 KJB <= JIN ; 
 MJA <=  LJA & kjb & lim  |  lja & KJB & lim  |  lja & kjb & LIM  |  LJA & KJB & LIM  ;
 mjm <=  LJA & kjb & lim  |  lja & KJB & lim  |  lja & kjb & LIM  |  lja & kjb & lim  ;
 KNA <=  JNA & jmn & jnb  |  jna & JMN & jnb  |  jna & jmn & JNB  |  JNA & JMN & JNB  ;
 knm <=  JNA & jmn & jnb  |  jna & JMN & jnb  |  jna & jmn & JNB  |  jna & jmn & jnb  ;
 KOB <= JNN ; 
 KKB <= JKA ; 
 KKC <= JJN ; 
 OEB <= NEA ; 
 OFA <= NEM ; 
 MVB <= KVA ; 
 MWA <= KVM ; 
 MYA <= KYA ; 
 CAY <= IAY ; 
 CBY <= IAY ; 
 CCY <= IAY ; 
 CDY <= IAY ; 
 OVB <= MVB ; 
 OWA <= MWA ; 
 OYA <= MYA ; 
 MMA <= LMA ; 
 MNA <= LMM ; 
 MNB <= LNA ; 
 MOA <= LNM ; 
 KVA <=  JUM & hum & hva  |  jum & HUM & hva  |  jum & hum & HVA  |  JUM & HUM & HVA  ;
 kvm <=  JUM & hum & hva  |  jum & HUM & hva  |  jum & hum & HVA  |  jum & hum & hva  ;
 DBD <= IBD ; 
 DCD <= IBD ; 
 DDD <= IBD ; 
 ONA <= MNA ; 
 ONB <= MNB ; 
 OOA <= MOA ; 
 KTA <=  JTA & htc & jsm  |  jta & HTC & jsm  |  jta & htc & JSM  |  JTA & HTC & JSM  ;
 ktm <=  JTA & htc & jsm  |  jta & HTC & jsm  |  jta & htc & JSM  |  jta & htc & jsm  ;
 KUA <=  JUA & jtm & hua  |  jua & JTM & hua  |  jua & jtm & HUA  |  JUA & JTM & HUA  ;
 kum <=  JUA & jtm & hua  |  jua & JTM & hua  |  jua & jtm & HUA  |  jua & jtm & hua  ;
 KYA <= HYA ; 
 KZA <= HYM ; 
 KZB <= HZA ; 
 DAZ <= IBZ ; 
 DBZ <= IBZ ; 
 DCZ <= IBZ ; 
 MTB <= KTA ; 
 MUA <= KTM ; 
 MUB <= KUA ; 
 MVA <= KUM ; 
 OTB <= MTB ; 
 OUA <= MUA ; 
 OUB <= MUB ; 
 OVA <= MVA ; 
 KSA <=  JSA & hsa & jrm  |  jsa & HSA & jrm  |  jsa & hsa & JRM  |  JSA & HSA & JRM  ;
 ksm <=  JSA & hsa & jrm  |  jsa & HSA & jrm  |  jsa & hsa & JRM  |  jsa & hsa & jrm  ;
 MOB <= LOA ; 
 MPA <= LOM ; 
 MSB <= KSA ; 
 MTA <= KSM ; 
 CAK <= IAK ; 
 CBK <= IAK ; 
 CCK <= IAK ; 
 CDK <= IAK ; 
 OJB <= MJA ; 
 OKA <= MJM ; 
 CAO <= IAO ; 
 CBO <= IAO ; 
 CCO <= IAO ; 
 CDO <= IAO ; 
 dhz <= ibz ; 
 TRG <= QRA ; 
 OTA <= MTA ; 
 OMB <= MMA ; 
 OOB <= MOB ; 
 OPA <= MPA ; 
 OSB <= MSB ; 
 DDZ <= IBZ ; 
 CAM <= IAM ; 
 CBM <= IAM ; 
 CCM <= IAM ; 
 CDM <= IAM ; 
 MZA <= KZA ; 
 MZB <= KZB ; 
 OZA <= MZA ; 
 OZB <= MZB ; 
 CAN <= IAN ; 
 CBN <= IAN ; 
 CCN <= IAN ; 
 CDN <= IAN ; 
 dez <= ibz ; 
 dfz <= ibz ; 
 dgz <= ibz ; 
 HGC <=  GFQ & ggd & fgg  |  gfq & GGD & fgg  |  gfq & ggd & FGG  |  GFQ & GGD & FGG  ;
 hgo <=  GFQ & ggd & fgg  |  gfq & GGD & fgg  |  gfq & ggd & FGG  |  gfq & ggd & fgg  ;
 HCA <=  GCA & gbn & gbm  |  gca & GBN & gbm  |  gca & gbn & GBM  |  GCA & GBN & GBM  ;
 hcm <=  GCA & gbn & gbm  |  gca & GBN & gbm  |  gca & gbn & GBM  |  gca & gbn & gbm  ;
 HCE <= GBO ; 
 HDA <=  GDA & gcm & gcn  |  gda & GCM & gcn  |  gda & gcm & GCN  |  GDA & GCM & GCN  ;
 hdm <=  GDA & gcm & gcn  |  gda & GCM & gcn  |  gda & gcm & GCN  |  gda & gcm & gcn  ;
 HDD <= GDC ; 
 HDC <=  GDE & gcq & fcr  |  gde & GCQ & fcr  |  gde & gcq & FCR  |  GDE & GCQ & FCR  ;
 hdo <=  GDE & gcq & fcr  |  gde & GCQ & fcr  |  gde & gcq & FCR  |  gde & gcq & fcr  ;
 HEB <=  GEB & gec & gdo  |  geb & GEC & gdo  |  geb & gec & GDO  |  GEB & GEC & GDO  ;
 hen <=  GEB & gec & gdo  |  geb & GEC & gdo  |  geb & gec & GDO  |  geb & gec & gdo  ;
 HGE <= GGA ; 
 HHB <=  GHC & ghb & ghd  |  ghc & GHB & ghd  |  ghc & ghb & GHD  |  GHC & GHB & GHD  ;
 hhn <=  GHC & ghb & ghd  |  ghc & GHB & ghd  |  ghc & ghb & GHD  |  ghc & ghb & ghd  ;
 HBB <=  GAN & gbd & fbh  |  gan & GBD & fbh  |  gan & gbd & FBH  |  GAN & GBD & FBH  ;
 hbn <=  GAN & gbd & fbh  |  gan & GBD & fbh  |  gan & gbd & FBH  |  gan & gbd & fbh  ;
 HBD <= GBC ; 
 HFB <=  GEO & gfc & gep  |  geo & GFC & gep  |  geo & gfc & GEP  |  GEO & GFC & GEP  ;
 hfn <=  GEO & gfc & gep  |  geo & GFC & gep  |  geo & gfc & GEP  |  geo & gfc & gep  ;
 HCC <=  GBP & gbr & gcd  |  gbp & GBR & gcd  |  gbp & gbr & GCD  |  GBP & GBR & GCD  ;
 hco <=  GBP & gbr & gcd  |  gbp & GBR & gcd  |  gbp & gbr & GCD  |  gbp & gbr & gcd  ;
 HAB <=  ILC & ilg & ilb  |  ilc & ILG & ilb  |  ilc & ilg & ILB  |  ILC & ILG & ILB  ;
 han <=  ILC & ilg & ilb  |  ilc & ILG & ilb  |  ilc & ilg & ILB  |  ilc & ilg & ilb  ;
 HCD <=  GCE & gbq & fci  |  gce & GBQ & fci  |  gce & gbq & FCI  |  GCE & GBQ & FCI  ;
 hcp <=  GCE & gbq & fci  |  gce & GBQ & fci  |  gce & gbq & FCI  |  gce & gbq & fci  ;
 HLA <=  GKM & gla & fkn  |  gkm & GLA & fkn  |  gkm & gla & FKN  |  GKM & GLA & FKN  ;
 hlm <=  GKM & gla & fkn  |  gkm & GLA & fkn  |  gkm & gla & FKN  |  gkm & gla & fkn  ;
 HMC <= FLP ; 
 HIA <=  GHM & gia & gho  |  ghm & GIA & gho  |  ghm & gia & GHO  |  GHM & GIA & GHO  ;
 him <=  GHM & gia & gho  |  ghm & GIA & gho  |  ghm & gia & GHO  |  ghm & gia & gho  ;
 HNA <=  GMM & gnb & gna  |  gmm & GNB & gna  |  gmm & gnb & GNA  |  GMM & GNB & GNA  ;
 hnm <=  GMM & gnb & gna  |  gmm & GNB & gna  |  gmm & gnb & GNA  |  gmm & gnb & gna  ;
 HQC <= GQA ; 
 HIB <=  GHN & gib & fhr  |  ghn & GIB & fhr  |  ghn & gib & FHR  |  GHN & GIB & FHR  ;
 hin <=  GHN & gib & fhr  |  ghn & GIB & fhr  |  ghn & gib & FHR  |  ghn & gib & fhr  ;
 HJC <= GIN ; 
 HMA <=  GLM & gma & gln  |  glm & GMA & gln  |  glm & gma & GLN  |  GLM & GMA & GLN  ;
 hmm <=  GLM & gma & gln  |  glm & GMA & gln  |  glm & gma & GLN  |  glm & gma & gln  ;
 HIC <=  GHP & gic & gid  |  ghp & GIC & gid  |  ghp & gic & GID  |  GHP & GIC & GID  ;
 hio <=  GHP & gic & gid  |  ghp & GIC & gid  |  ghp & gic & GID  |  ghp & gic & gid  ;
 HKB <=  GKB & fke & gkc  |  gkb & FKE & gkc  |  gkb & fke & GKC  |  GKB & FKE & GKC  ;
 hkn <=  GKB & fke & gkc  |  gkb & FKE & gkc  |  gkb & fke & GKC  |  gkb & fke & gkc  ;
 HNC <= FMP ; 
 HHC <=  GGP & ghe & ggo  |  ggp & GHE & ggo  |  ggp & ghe & GGO  |  GGP & GHE & GGO  ;
 hho <=  GGP & ghe & ggo  |  ggp & GHE & ggo  |  ggp & ghe & GGO  |  ggp & ghe & ggo  ;
 HJD <= GIP ; 
 HJB <=  GJD & gio & gjc  |  gjd & GIO & gjc  |  gjd & gio & GJC  |  GJD & GIO & GJC  ;
 hjn <=  GJD & gio & gjc  |  gjd & GIO & gjc  |  gjd & gio & GJC  |  gjd & gio & gjc  ;
 HLC <=  GLC & gko & gkp  |  glc & GKO & gkp  |  glc & gko & GKP  |  GLC & GKO & GKP  ;
 hlo <=  GLC & gko & gkp  |  glc & GKO & gkp  |  glc & gko & GKP  |  glc & gko & gkp  ;
 HPC <= GPA ; 
 HUA <=  GTM & gua & ftn  |  gtm & GUA & ftn  |  gtm & gua & FTN  |  GTM & GUA & FTN  ;
 hum <=  GTM & gua & ftn  |  gtm & GUA & ftn  |  gtm & gua & FTN  |  gtm & gua & ftn  ;
 HTC <= GTA ; 
 QAX <=  IKJ & TTB  |  IKK & ttb  |  QIB  ; 
 CAZ <= IAZ ; 
 CBZ <= IAZ ; 
 CCZ <= IAZ ; 
 CDZ <= IAZ ; 
 qak <= qib ; 
 qal <= qib ; 
 DAE <= IBE ; 
 DCE <= IBE ; 
 DDE <= IBE ; 
 HYA <=  GXM & fxm & fya  |  gxm & FXM & fya  |  gxm & fxm & FYA  |  GXM & FXM & FYA  ;
 hym <=  GXM & fxm & fya  |  gxm & FXM & fya  |  gxm & fxm & FYA  |  gxm & fxm & fya  ;
 HZA <= GZA ; 
 QAO <=  IKA & TTA  |  IKB & tta  |  QIE  ; 
 QAR <=  IKD & TTA  |  IKE & tta  |  QIE  ; 
 QAU <=  IKG & TTB  |  IKH & ttb  |  QIC  ; 
 QAZ <=  IKL & TTB  |  IKM & ttb  |  QIC  ; 
 KZM <= HZM ; 
 OZM <= MZM ; 
 QIA <= IIA ; 
 HUB <= GTN ; 
 HUC <= FTM ; 
 HXB <= GXA ; 
 qah <= qic ; 
 qai <= qic ; 
 CAW <= IAW ; 
 CBW <= IAW ; 
 CCW <= IAW ; 
 CDW <= IAW ; 
 QIB <= QIA ; 
 QIC <= QIA ; 
 QID <= QIA ; 
 QIE <= QIA ; 
 CAR <= IAR ; 
 CBR <= IAR ; 
 CCR <= IAR ; 
 CDR <= IAR ; 
 HRB <=  GRB & gqn & gqo  |  grb & GQN & gqo  |  grb & gqn & GQO  |  GRB & GQN & GQO  ;
 hrn <=  GRB & gqn & gqo  |  grb & GQN & gqo  |  grb & gqn & GQO  |  grb & gqn & gqo  ;
 HSB <= GRN ; 
 qae <= qid ; 
 qaf <= qid ; 
 HZM <= GZM ; 
 MZM <= KZM ; 
 HMB <=  GLO & gmb & gmc  |  glo & GMB & gmc  |  glo & gmb & GMC  |  GLO & GMB & GMC  ;
 hmn <=  GLO & gmb & gmc  |  glo & GMB & gmc  |  glo & gmb & GMC  |  glo & gmb & gmc  ;
 HND <= FNC ; 
 TRH <= QRA ; 
 qaa <= qie & isa ; 
 qab <= qie & isb ; 
 qac <= qie & isc ; 
 CAL <= IAL ; 
 CBL <= IAL ; 
 CCL <= IAL ; 
 CDL <= IAL ; 
 FBE <=  EBW & ebx & eby  |  ebw & EBX & eby  |  ebw & ebx & EBY  |  EBW & EBX & EBY  ;
 fbq <=  EBW & ebx & eby  |  ebw & EBX & eby  |  ebw & ebx & EBY  |  ebw & ebx & eby  ;
 FCE <=  ECC & ecd & ece  |  ecc & ECD & ece  |  ecc & ecd & ECE  |  ECC & ECD & ECE  ;
 fcq <=  ECC & ecd & ece  |  ecc & ECD & ece  |  ecc & ecd & ECE  |  ecc & ecd & ece  ;
 FGE <=  EGG & egh & egi  |  egg & EGH & egi  |  egg & egh & EGI  |  EGG & EGH & EGI  ;
 fgq <=  EGG & egh & egi  |  egg & EGH & egi  |  egg & egh & EGI  |  egg & egh & egi  ;
 FKC <=  EKK & ekl & ekm  |  ekk & EKL & ekm  |  ekk & ekl & EKM  |  EKK & EKL & EKM  ;
 fko <=  EKK & ekl & ekm  |  ekk & EKL & ekm  |  ekk & ekl & EKM  |  ekk & ekl & ekm  ;
 FAE <=  EAS & eat & eau  |  eas & EAT & eau  |  eas & eat & EAU  |  EAS & EAT & EAU  ;
 faq <=  EAS & eat & eau  |  eas & EAT & eau  |  eas & eat & EAU  |  eas & eat & eau  ;
 FEI <= QAE ; 
 FDE <=  EDG & edh & edi  |  edg & EDH & edi  |  edg & edh & EDI  |  EDG & EDH & EDI  ;
 fdq <=  EDG & edh & edi  |  edg & EDH & edi  |  edg & edh & EDI  |  edg & edh & edi  ;
 FED <=  EEW & eex & eey  |  eew & EEX & eey  |  eew & eex & EEY  |  EEW & EEX & EEY  ;
 fep <=  EEW & eex & eey  |  eew & EEX & eey  |  eew & eex & EEY  |  eew & eex & eey  ;
 FHC <=  EHK & ehl & ehm  |  ehk & EHL & ehm  |  ehk & ehl & EHM  |  EHK & EHL & EHM  ;
 fho <=  EHK & ehl & ehm  |  ehk & EHL & ehm  |  ehk & ehl & EHM  |  ehk & ehl & ehm  ;
 FHH <= QAH ; 
 FAF <=  EAG & eah & eai  |  eag & EAH & eai  |  eag & eah & EAI  |  EAG & EAH & EAI  ;
 far <=  EAG & eah & eai  |  eag & EAH & eai  |  eag & eah & EAI  |  eag & eah & eai  ;
 FDF <=  EDS & edt & edu  |  eds & EDT & edu  |  eds & edt & EDU  |  EDS & EDT & EDU  ;
 fdr <=  EDS & edt & edu  |  eds & EDT & edu  |  eds & edt & EDU  |  eds & edt & edu  ;
 FEE <=  EEK & eel & eem  |  eek & EEL & eem  |  eek & eel & EEM  |  EEK & EEL & EEM  ;
 feq <=  EEK & eel & eem  |  eek & EEL & eem  |  eek & eel & EEM  |  eek & eel & eem  ;
 FHD <=  EHW & ehx & ehy  |  ehw & EHX & ehy  |  ehw & ehx & EHY  |  EHW & EHX & EHY  ;
 fhp <=  EHW & ehx & ehy  |  ehw & EHX & ehy  |  ehw & ehx & EHY  |  ehw & ehx & ehy  ;
 FFH <= QAF ; 
 FAG <=  EAY & eaz & qaa  |  eay & EAZ & qaa  |  eay & eaz & QAA  |  EAY & EAZ & QAA  ;
 fas <=  EAY & eaz & qaa  |  eay & EAZ & qaa  |  eay & eaz & QAA  |  eay & eaz & qaa  ;
 FBJ <= QAB ; 
 FBF <=  EBK & ebl & ebm  |  ebk & EBL & ebm  |  ebk & ebl & EBM  |  EBK & EBL & EBM  ;
 fbr <=  EBK & ebl & ebm  |  ebk & EBL & ebm  |  ebk & ebl & EBM  |  ebk & ebl & ebm  ;
 FCI <= QAC ; 
 FCF <=  ECO & ecp & ecq  |  eco & ECP & ecq  |  eco & ecp & ECQ  |  ECO & ECP & ECQ  ;
 fcr <=  ECO & ecp & ecq  |  eco & ECP & ecq  |  eco & ecp & ECQ  |  eco & ecp & ecq  ;
 FFE <=  EFO & efp & efq  |  efo & EFP & efq  |  efo & efp & EFQ  |  EFO & EFP & EFQ  ;
 ffq <=  EFO & efp & efq  |  efo & EFP & efq  |  efo & efp & EFQ  |  efo & efp & efq  ;
 HXA <= GWM ; 
 FOC <=  EOO & eop & eoq  |  eoo & EOP & eoq  |  eoo & eop & EOQ  |  EOO & EOP & EOQ  ;
 foo <=  EOO & eop & eoq  |  eoo & EOP & eoq  |  eoo & eop & EOQ  |  eoo & eop & eoq  ;
 FKG <= QAK ; 
 FSC <=  ESS & est & esu  |  ess & EST & esu  |  ess & est & ESU  |  ESS & EST & ESU  ;
 fso <=  ESS & est & esu  |  ess & EST & esu  |  ess & est & ESU  |  ess & est & esu  ;
 FLF <= QAL ; 
 FWA <=  EWW & ewx & ewy  |  eww & EWX & ewy  |  eww & ewx & EWY  |  EWW & EWX & EWY  ;
 fwm <=  EWW & ewx & ewy  |  eww & EWX & ewy  |  eww & ewx & EWY  |  eww & ewx & ewy  ;
 FZB <= QAZ ; 
 FLC <=  ELO & elp & elq  |  elo & ELP & elq  |  elo & elp & ELQ  |  ELO & ELP & ELQ  ;
 flo <=  ELO & elp & elq  |  elo & ELP & elq  |  elo & elp & ELQ  |  elo & elp & elq  ;
 FIG <= QAI ; 
 FPC <=  EPS & ept & epu  |  eps & EPT & epu  |  eps & ept & EPU  |  EPS & EPT & EPU  ;
 fpo <=  EPS & ept & epu  |  eps & EPT & epu  |  eps & ept & EPU  |  eps & ept & epu  ;
 FTA <=  ETW & etx & ety  |  etw & ETX & ety  |  etw & etx & ETY  |  ETW & ETX & ETY  ;
 ftm <=  ETW & etx & ety  |  etw & ETX & ety  |  etw & etx & ETY  |  etw & etx & ety  ;
 FNE <= ENZ ; 
 FID <=  EIO & eip & eiq  |  eio & EIP & eiq  |  eio & eip & EIQ  |  EIO & EIP & EIQ  ;
 fip <=  EIO & eip & eiq  |  eio & EIP & eiq  |  eio & eip & EIQ  |  eio & eip & eiq  ;
 FMD <=  EMS & emt & emu  |  ems & EMT & emu  |  ems & emt & EMU  |  EMS & EMT & EMU  ;
 fmp <=  EMS & emt & emu  |  ems & EMT & emu  |  ems & emt & EMU  |  ems & emt & emu  ;
 FGF <=  EGS & egt & egu  |  egs & EGT & egu  |  egs & egt & EGU  |  EGS & EGT & EGU  ;
 fgr <=  EGS & egt & egu  |  egs & EGT & egu  |  egs & egt & EGU  |  egs & egt & egu  ;
 FJE <=  EJS & ejt & eju  |  ejs & EJT & eju  |  ejs & ejt & EJU  |  EJS & EJT & EJU  ;
 fjq <=  EJS & ejt & eju  |  ejs & EJT & eju  |  ejs & ejt & EJU  |  ejs & ejt & eju  ;
 FKD <=  EKW & ekx & eky  |  ekw & EKX & eky  |  ekw & ekx & EKY  |  EKW & EKX & EKY  ;
 fkp <=  EKW & ekx & eky  |  ekw & EKX & eky  |  ekw & ekx & EKY  |  ekw & ekx & eky  ;
 CAE <=  IAE & TRC  |  ICE & trc  ; 
 CBE <=  IAE & TRC  |  ICE & trc  ; 
 CCE <=  IAE & TRC  |  ICE & trc  ; 
 CBC <=  IAC & TRC  |  ICC & trc  ; 
 CCC <=  IAC & TRC  |  ICC & trc  ; 
 CDC <=  IAC & TRC  |  ICC & trc  ; 
 DAI <= IBI ; 
 DCI <= IBI ; 
 DDI <= IBI ; 
 cde <= iae & TRC |  ice & trc ; 
 cdh <= iah & TRC |  ich & trc ; 
 CAT <= IAT ; 
 DBH <= IBH ; 
 DCH <= IBH ; 
 DDH <= IBH ; 
 dgu <= ibu ; 
 dgx <= ibx ; 
 dhu <= ibu ; 
 dhx <= ibx ; 
 dgl <= ibl ; 
 dhl <= ibl ; 
 dky <= iby ; 
 CAH <=  IAH & TRC  |  ICH & trc  ; 
 CBH <=  IAH & TRC  |  ICH & trc  ; 
 CCH <=  IAH & TRC  |  ICH & trc  ; 
 DAM <= IBM ; 
 DCM <= IBM ; 
 DDM <= IBM ; 
 DEM <= IBM ; 
 dgm <= ibm ; 
 dgy <= iby ; 
 dhm <= ibm ; 
 dhy <= iby ; 
 CAS <= IAS ; 
 CBS <= IAS ; 
 CCS <= IAS ; 
 CDS <= IAS ; 
 DAY <= IBY ; 
 DCY <= IBY ; 
 DDY <= IBY ; 
 DEY <= IBY ; 
 CAJ <=  IAJ & TRC  |  ICJ & trc  ; 
 CBJ <=  IAJ & TRC  |  ICJ & trc  ; 
 CCJ <=  IAJ & TRC  |  ICJ & trc  ; 
 CCA <= IAA & TRC |  ICA & trc ; 
 cdj <= iaj & TRC |  icj & trc ; 
 FQB <=  EQW & eqx & eqy  |  eqw & EQX & eqy  |  eqw & eqx & EQY  |  EQW & EQX & EQY  ;
 fqn <=  EQW & eqx & eqy  |  eqw & EQX & eqy  |  eqw & eqx & EQY  |  eqw & eqx & eqy  ;
 DAU <= IBU ; 
 DCU <= IBU ; 
 DDU <= IBU ; 
 DEU <= IBU ; 
 CBT <= IAT ; 
 CCT <= IAT ; 
 CDT <= IAT ; 
 TRC <= QRA ; 
 DBX <= IBX ; 
 DCX <= IBX ; 
 DDX <= IBX ; 
 DFX <= IBX ; 
 DBL <= IBL ; 
 DCL <= IBL ; 
 DDL <= IBL ; 
 DFL <= IBL ; 
 FNC <=  ENW & enx & eny  |  enw & ENX & eny  |  enw & enx & ENY  |  ENW & ENX & ENY  ;
 fno <=  ENW & enx & eny  |  enw & ENX & eny  |  enw & enx & ENY  |  enw & enx & eny  ;
 DBT <= IBT ; 
 DCT <= IBT ; 
 DDT <= IBT ; 
 DFT <= IBT ; 
 dgt <= ibt ; 
 dht <= ibt ; 
 FCG <=  ECX & ecy & ecz  |  ecx & ECY & ecz  |  ecx & ecy & ECZ  |  ECX & ECY & ECZ  ;
 fcs <=  ECX & ecy & ecz  |  ecx & ECY & ecz  |  ecx & ecy & ECZ  |  ecx & ecy & ecz  ;
 FBI <= EBZ ; 
 FDG <=  EDD & ede & edf  |  edd & EDE & edf  |  edd & ede & EDF  |  EDD & EDE & EDF  ;
 fds <=  EDD & ede & edf  |  edd & EDE & edf  |  edd & ede & EDF  |  edd & ede & edf  ;
 FHE <=  EHH & ehi & ehj  |  ehh & EHI & ehj  |  ehh & ehi & EHJ  |  EHH & EHI & EHJ  ;
 fhq <=  EHH & ehi & ehj  |  ehh & EHI & ehj  |  ehh & ehi & EHJ  |  ehh & ehi & ehj  ;
 FAH <=  EAD & eae & eaf  |  ead & EAE & eaf  |  ead & eae & EAF  |  EAD & EAE & EAF  ;
 fat <=  EAD & eae & eaf  |  ead & EAE & eaf  |  ead & eae & EAF  |  ead & eae & eaf  ;
 FBG <=  EBT & ebu & ebv  |  ebt & EBU & ebv  |  ebt & ebu & EBV  |  EBT & EBU & EBV  ;
 fbs <=  EBT & ebu & ebv  |  ebt & EBU & ebv  |  ebt & ebu & EBV  |  ebt & ebu & ebv  ;
 FEF <=  EEH & eei & eej  |  eeh & EEI & eej  |  eeh & eei & EEJ  |  EEH & EEI & EEJ  ;
 fer <=  EEH & eei & eej  |  eeh & EEI & eej  |  eeh & eei & EEJ  |  eeh & eei & eej  ;
 FFF <=  EFX & efy & efz  |  efx & EFY & efz  |  efx & efy & EFZ  |  EFX & EFY & EFZ  ;
 ffr <=  EFX & efy & efz  |  efx & EFY & efz  |  efx & efy & EFZ  |  efx & efy & efz  ;
 FAI <=  EAP & eaq & ear  |  eap & EAQ & ear  |  eap & eaq & EAR  |  EAP & EAQ & EAR  ;
 fau <=  EAP & eaq & ear  |  eap & EAQ & ear  |  eap & eaq & EAR  |  eap & eaq & ear  ;
 FBH <=  EBH & ebi & ebj  |  ebh & EBI & ebj  |  ebh & ebi & EBJ  |  EBH & EBI & EBJ  ;
 fbt <=  EBH & ebi & ebj  |  ebh & EBI & ebj  |  ebh & ebi & EBJ  |  ebh & ebi & ebj  ;
 FEG <=  EET & eeu & eev  |  eet & EEU & eev  |  eet & eeu & EEV  |  EET & EEU & EEV  ;
 fes <=  EET & eeu & eev  |  eet & EEU & eev  |  eet & eeu & EEV  |  eet & eeu & eev  ;
 FFG <=  EFL & efm & efn  |  efl & EFM & efn  |  efl & efm & EFN  |  EFL & EFM & EFN  ;
 ffs <=  EFL & efm & efn  |  efl & EFM & efn  |  efl & efm & EFN  |  efl & efm & efn  ;
 FCH <=  ECL & ecm & ecn  |  ecl & ECM & ecn  |  ecl & ecm & ECN  |  ECL & ECM & ECN  ;
 fct <=  ECL & ecm & ecn  |  ecl & ECM & ecn  |  ecl & ecm & ECN  |  ecl & ecm & ecn  ;
 FDH <=  EDP & edq & edr  |  edp & EDQ & edr  |  edp & edq & EDR  |  EDP & EDQ & EDR  ;
 fdt <=  EDP & edq & edr  |  edp & EDQ & edr  |  edp & edq & EDR  |  edp & edq & edr  ;
 FGG <=  EGP & egq & egr  |  egp & EGQ & egr  |  egp & egq & EGR  |  EGP & EGQ & EGR  ;
 fgs <=  EGP & egq & egr  |  egp & EGQ & egr  |  egp & egq & EGR  |  egp & egq & egr  ;
 FHF <=  EHT & ehu & ehv  |  eht & EHU & ehv  |  eht & ehu & EHV  |  EHT & EHU & EHV  ;
 fhr <=  EHT & ehu & ehv  |  eht & EHU & ehv  |  eht & ehu & EHV  |  eht & ehu & ehv  ;
 FLD <=  ELL & elm & eln  |  ell & ELM & eln  |  ell & elm & ELN  |  ELL & ELM & ELN  ;
 flp <=  ELL & elm & eln  |  ell & ELM & eln  |  ell & elm & ELN  |  ell & elm & eln  ;
 FPD <=  EPP & epq & epr  |  epp & EPQ & epr  |  epp & epq & EPR  |  EPP & EPQ & EPR  ;
 fpp <=  EPP & epq & epr  |  epp & EPQ & epr  |  epp & epq & EPR  |  epp & epq & epr  ;
 FTB <=  ETT & etu & etv  |  ett & ETU & etv  |  ett & etu & ETV  |  ETT & ETU & ETV  ;
 ftn <=  ETT & etu & etv  |  ett & ETU & etv  |  ett & etu & ETV  |  ett & etu & etv  ;
 FIE <=  EIL & eim & ein  |  eil & EIM & ein  |  eil & eim & EIN  |  EIL & EIM & EIN  ;
 fiq <=  EIL & eim & ein  |  eil & EIM & ein  |  eil & eim & EIN  |  eil & eim & ein  ;
 FME <=  EMP & emq & emr  |  emp & EMQ & emr  |  emp & emq & EMR  |  EMP & EMQ & EMR  ;
 fmq <=  EMP & emq & emr  |  emp & EMQ & emr  |  emp & emq & EMR  |  emp & emq & emr  ;
 FQC <=  EQT & equ & eqv  |  eqt & EQU & eqv  |  eqt & equ & EQV  |  EQT & EQU & EQV  ;
 fqo <=  EQT & equ & eqv  |  eqt & EQU & eqv  |  eqt & equ & EQV  |  eqt & equ & eqv  ;
 FIF <=  EIX & eiy & eiz  |  eix & EIY & eiz  |  eix & eiy & EIZ  |  EIX & EIY & EIZ  ;
 fir <=  EIX & eiy & eiz  |  eix & EIY & eiz  |  eix & eiy & EIZ  |  eix & eiy & eiz  ;
 FJF <=  EJP & ejq & ejr  |  ejp & EJQ & ejr  |  ejp & ejq & EJR  |  EJP & EJQ & EJR  ;
 fjr <=  EJP & ejq & ejr  |  ejp & EJQ & ejr  |  ejp & ejq & EJR  |  ejp & ejq & ejr  ;
 FND <=  ENT & enu & env  |  ent & ENU & env  |  ent & enu & ENV  |  ENT & ENU & ENV  ;
 fnp <=  ENT & enu & env  |  ent & ENU & env  |  ent & enu & ENV  |  ent & enu & env  ;
 FRD <= QAR ; 
 FKE <=  EKT & eku & ekv  |  ekt & EKU & ekv  |  ekt & eku & EKV  |  EKT & EKU & EKV  ;
 fkq <=  EKT & eku & ekv  |  ekt & EKU & ekv  |  ekt & eku & EKV  |  ekt & eku & ekv  ;
 FLE <=  ELX & ely & elz  |  elx & ELY & elz  |  elx & ely & ELZ  |  ELX & ELY & ELZ  ;
 flq <=  ELX & ely & elz  |  elx & ELY & elz  |  elx & ely & ELZ  |  elx & ely & elz  ;
 FOD <=  EOX & eoy & eoz  |  eox & EOY & eoz  |  eox & eoy & EOZ  |  EOX & EOY & EOZ  ;
 fop <=  EOX & eoy & eoz  |  eox & EOY & eoz  |  eox & eoy & EOZ  |  eox & eoy & eoz  ;
 FOE <= QAO ; 
 FXA <=  EXX & exy & exz  |  exx & EXY & exz  |  exx & exy & EXZ  |  EXX & EXY & EXZ  ;
 fxm <=  EXX & exy & exz  |  exx & EXY & exz  |  exx & exy & EXZ  |  exx & exy & exz  ;
 FZA <= EZZ ; 
 FUB <=  EUX & euy & euz  |  eux & EUY & euz  |  eux & euy & EUZ  |  EUX & EUY & EUZ  ;
 fun <=  EUX & euy & euz  |  eux & EUY & euz  |  eux & euy & EUZ  |  eux & euy & euz  ;
 CCB <= IAB & TRD |  ICB & trd ; 
 CDB <= IAB & TRD |  ICB & trd ; 
 FRC <=  ERX & ery & erz  |  erx & ERY & erz  |  erx & ery & ERZ  |  ERX & ERY & ERZ  ;
 fro <=  ERX & ery & erz  |  erx & ERY & erz  |  erx & ery & ERZ  |  erx & ery & erz  ;
 TRD <= QRA ; 
 DBP <= IBP ; 
 DCP <= IBP ; 
 DDP <= IBP ; 
 DFP <= IBP ; 
 dgp <= ibp ; 
 dhp <= ibp ; 
 DAQ <= IBQ ; 
 DCQ <= IBQ ; 
 DDQ <= IBQ ; 
 DEQ <= IBQ ; 
 dgq <= ibq ; 
 dhq <= ibq ; 
end 
endmodule;
