module td( IZZ,
 IAA, 
 IAB, 
 IAC, 
 IAD, 
 IAE, 
 IAF, 
 IAG, 
 IAH, 
 IAI, 
 IAJ, 
 IAK, 
 IAL, 
 IAM, 
 IAN, 
 IAO, 
 IAP, 
 IAQ, 
 IAR, 
 IAS, 
 IAT, 
 IAU, 
 IAV, 
 IAW, 
 IAX, 
 IBA, 
 IBB, 
 IBC, 
 IBD, 
 IBE, 
 IBF, 
 IBG, 
 IBH, 
 IBI, 
 IBJ, 
 IBK, 
 IBL, 
 IBM, 
 IBN, 
 IBO, 
 IBP, 
 IBQ, 
 IBR, 
 IBS, 
 IBT, 
 IBU, 
 IBV, 
 IBW, 
 IBX, 
 ICA, 
 ICB, 
 ICC, 
 ICD, 
 ICE, 
 ICF, 
 ICG, 
 ICH, 
 ICI, 
 ICJ, 
 ICK, 
 ICL, 
 ICM, 
 ICN, 
 ICO, 
 ICP, 
 ICQ, 
 ICR, 
 ICS, 
 ICT, 
 ICU, 
 ICV, 
 ICW, 
 ICX, 
 IDA, 
 IDB, 
 IDC, 
 IDD, 
 IDE, 
 IDF, 
 IDG, 
 IDH, 
 IDI, 
 IDJ, 
 IDK, 
 IDL, 
 IDM, 
 IDN, 
 IDO, 
 IDP, 
 IDQ, 
 IDR, 
 IDS, 
 IDT, 
 IDU, 
 IDV, 
 IDW, 
 IDX, 
 IEA, 
 IEB, 
 IEC, 
 IED, 
 IEE, 
 IEF, 
 IFA, 
 IFB, 
 IFC, 
 IFD, 
 IFE, 
 IFFF , 
 IGA, 
 IGB, 
 IGC, 
 IGD, 
 IGE, 
 IGF, 
 IHA, 
 IHB, 
 IHC, 
 IHD, 
 IHE, 
 IHF, 
 IIA, 
 IJA, 
 OAA, 
 OAB, 
 OAC, 
 OAD, 
 OAE, 
 OAF, 
 OAG, 
 OAH, 
 OAI, 
 OAJ, 
 OAK, 
 OAL, 
 OAM, 
 OAN, 
 OAO, 
 OAP, 
 OBA, 
 OBB, 
 OBC, 
 OBD, 
 OBE, 
 OBF, 
 OBG, 
 OBH, 
 OBI, 
 OBJ, 
 OBK, 
 OBL, 
 OBM, 
 OBN, 
 OBO, 
 OBP, 
 OCA, 
 OCB, 
 OCC, 
 OCD, 
 OCE, 
 OCF, 
 OCG, 
 OCH, 
 OCI, 
 OCJ, 
 OCK, 
 OCL, 
 OCM, 
 OCN, 
 OCO, 
 OCP, 
 ODA, 
 ODB, 
 ODC, 
 ODD, 
 ODE, 
 ODF, 
 ODG, 
 ODH, 
 ODI, 
 ODJ, 
 ODK, 
 ODL, 
 ODM, 
 ODN, 
 ODO, 
 ODP, 
 OEA, 
 OEB, 
 OEC, 
 OED, 
 OEE, 
 OEF, 
 OEG, 
 OEH, 
 OEI, 
 OEJ, 
 OEK, 
 OEL, 
 OEM, 
 OEN, 
 OEO, 
 OEP, 
 OFA, 
 OFB, 
 OFC, 
 OFD, 
 OFE, 
 OFF, 
 OFG, 
 OFH, 
 OFI, 
 OFJ, 
 OFK, 
 OFL, 
 OFM, 
 OFN, 
 OFO, 
 OFP, 
 OGA, 
 OGB, 
 OGC, 
 OGD, 
 OGE, 
 OGF, 
 OGG, 
 OGH, 
 OGI, 
 OGJ, 
 OGK, 
 OGL, 
 OGM, 
 OGN, 
 OGO, 
 OGP, 
 OHA, 
 OHB, 
 OHC, 
 OHD, 
 OHE, 
 OHF, 
 OHG, 
 OHH, 
 OHI, 
 OHJ, 
 OHK, 
 OHL, 
 OHM, 
 OHN, 
 OHO, 
 OHP, 
 OIA, 
 OIB, 
 OIC, 
 OID, 
 OIE, 
 OIF, 
 OIG, 
 OIH, 
 OJA, 
 OKA, 
 OKB, 
 OKC, 
 OKD, 
 OKE, 
 OLA, 
 OLB, 
 OLC, 
 OLD, 
 OLE, 
 OMA, 
 OMB, 
 OMC, 
 OMD, 
 ONA, 
 ONB, 
 ONC, 
 OOA, 
 OOB, 
 OOC, 
OPA ); 
    
 input IZZ; 
 input IAA; 
 input IAB; 
 input IAC; 
 input IAD; 
 input IAE; 
 input IAF; 
 input IAG; 
 input IAH; 
 input IAI; 
 input IAJ; 
 input IAK; 
 input IAL; 
 input IAM; 
 input IAN; 
 input IAO; 
 input IAP; 
 input IAQ; 
 input IAR; 
 input IAS; 
 input IAT; 
 input IAU; 
 input IAV; 
 input IAW; 
 input IAX; 
 input IBA; 
 input IBB; 
 input IBC; 
 input IBD; 
 input IBE; 
 input IBF; 
 input IBG; 
 input IBH; 
 input IBI; 
 input IBJ; 
 input IBK; 
 input IBL; 
 input IBM; 
 input IBN; 
 input IBO; 
 input IBP; 
 input IBQ; 
 input IBR; 
 input IBS; 
 input IBT; 
 input IBU; 
 input IBV; 
 input IBW; 
 input IBX; 
 input ICA; 
 input ICB; 
 input ICC; 
 input ICD; 
 input ICE; 
 input ICF; 
 input ICG; 
 input ICH; 
 input ICI; 
 input ICJ; 
 input ICK; 
 input ICL; 
 input ICM; 
 input ICN; 
 input ICO; 
 input ICP; 
 input ICQ; 
 input ICR; 
 input ICS; 
 input ICT; 
 input ICU; 
 input ICV; 
 input ICW; 
 input ICX; 
 input IDA; 
 input IDB; 
 input IDC; 
 input IDD; 
 input IDE; 
 input IDF; 
 input IDG; 
 input IDH; 
 input IDI; 
 input IDJ; 
 input IDK; 
 input IDL; 
 input IDM; 
 input IDN; 
 input IDO; 
 input IDP; 
 input IDQ; 
 input IDR; 
 input IDS; 
 input IDT; 
 input IDU; 
 input IDV; 
 input IDW; 
 input IDX; 
 input IEA; 
 input IEB; 
 input IEC; 
 input IED; 
 input IEE; 
 input IEF; 
 input IFA; 
 input IFB; 
 input IFC; 
 input IFD; 
 input IFE; 
 input IFFF ; 
 input IGA; 
 input IGB; 
 input IGC; 
 input IGD; 
 input IGE; 
 input IGF; 
 input IHA; 
 input IHB; 
 input IHC; 
 input IHD; 
 input IHE; 
 input IHF; 
 input IIA; 
 input IJA; 
 output OAA; 
 output OAB; 
 output OAC; 
 output OAD; 
 output OAE; 
 output OAF; 
 output OAG; 
 output OAH; 
 output OAI; 
 output OAJ; 
 output OAK; 
 output OAL; 
 output OAM; 
 output OAN; 
 output OAO; 
 output OAP; 
 output OBA; 
 output OBB; 
 output OBC; 
 output OBD; 
 output OBE; 
 output OBF; 
 output OBG; 
 output OBH; 
 output OBI; 
 output OBJ; 
 output OBK; 
 output OBL; 
 output OBM; 
 output OBN; 
 output OBO; 
 output OBP; 
 output OCA; 
 output OCB; 
 output OCC; 
 output OCD; 
 output OCE; 
 output OCF; 
 output OCG; 
 output OCH; 
 output OCI; 
 output OCJ; 
 output OCK; 
 output OCL; 
 output OCM; 
 output OCN; 
 output OCO; 
 output OCP; 
 output ODA; 
 output ODB; 
 output ODC; 
 output ODD; 
 output ODE; 
 output ODF; 
 output ODG; 
 output ODH; 
 output ODI; 
 output ODJ; 
 output ODK; 
 output ODL; 
 output ODM; 
 output ODN; 
 output ODO; 
 output ODP; 
 output OEA; 
 output OEB; 
 output OEC; 
 output OED; 
 output OEE; 
 output OEF; 
 output OEG; 
 output OEH; 
 output OEI; 
 output OEJ; 
 output OEK; 
 output OEL; 
 output OEM; 
 output OEN; 
 output OEO; 
 output OEP; 
 output OFA; 
 output OFB; 
 output OFC; 
 output OFD; 
 output OFE; 
 output OFF; 
 output OFG; 
 output OFH; 
 output OFI; 
 output OFJ; 
 output OFK; 
 output OFL; 
 output OFM; 
 output OFN; 
 output OFO; 
 output OFP; 
 output OGA; 
 output OGB; 
 output OGC; 
 output OGD; 
 output OGE; 
 output OGF; 
 output OGG; 
 output OGH; 
 output OGI; 
 output OGJ; 
 output OGK; 
 output OGL; 
 output OGM; 
 output OGN; 
 output OGO; 
 output OGP; 
 output OHA; 
 output OHB; 
 output OHC; 
 output OHD; 
 output OHE; 
 output OHF; 
 output OHG; 
 output OHH; 
 output OHI; 
 output OHJ; 
 output OHK; 
 output OHL; 
 output OHM; 
 output OHN; 
 output OHO; 
 output OHP; 
 output OIA; 
 output OIB; 
 output OIC; 
 output OID; 
 output OIE; 
 output OIF; 
 output OIG; 
 output OIH; 
 output OJA; 
 output OKA; 
 output OKB; 
 output OKC; 
 output OKD; 
 output OKE; 
 output OLA; 
 output OLB; 
 output OLC; 
 output OLD; 
 output OLE; 
 output OMA; 
 output OMB; 
 output OMC; 
 output OMD; 
 output ONA; 
 output ONB; 
 output ONC; 
 output OOA; 
 output OOB; 
 output OOC; 
 output OPA; 
  
  
reg  aaa ;
reg  aab ;
reg  aac ;
reg  aad ;
reg  aae ;
reg  aaf ;
reg  aag ;
reg  aah ;
reg  aai ;
reg  aaj ;
reg  aak ;
reg  aal ;
reg  aam ;
reg  aan ;
reg  aao ;
reg  aap ;
reg  aaq ;
reg  aar ;
reg  aas ;
reg  aat ;
reg  aau ;
reg  aav ;
reg  aaw ;
reg  aax ;
reg  aba ;
reg  abb ;
reg  abc ;
reg  abd ;
reg  abe ;
reg  abf ;
reg  abg ;
reg  abh ;
reg  abi ;
reg  abj ;
reg  abk ;
reg  abl ;
reg  abm ;
reg  abn ;
reg  abo ;
reg  abp ;
reg  abq ;
reg  abr ;
reg  abs ;
reg  abt ;
reg  abu ;
reg  abv ;
reg  abw ;
reg  abx ;
reg  aca ;
reg  acb ;
reg  acc ;
reg  acd ;
reg  ace ;
reg  acf ;
reg  acg ;
reg  ach ;
reg  aci ;
reg  acj ;
reg  ack ;
reg  acl ;
reg  acm ;
reg  acn ;
reg  aco ;
reg  acp ;
reg  acq ;
reg  acr ;
reg  acs ;
reg  act ;
reg  acu ;
reg  acv ;
reg  acw ;
reg  acx ;
reg  ada ;
reg  adb ;
reg  adc ;
reg  add ;
reg  ade ;
reg  adf ;
reg  adg ;
reg  adh ;
reg  adi ;
reg  adj ;
reg  adk ;
reg  adl ;
reg  adm ;
reg  adn ;
reg  ado ;
reg  adp ;
reg  adq ;
reg  adr ;
reg  ads ;
reg  adt ;
reg  adu ;
reg  adv ;
reg  adw ;
reg  adx ;
reg  BAA ;
reg  BAB ;
reg  BAC ;
reg  BAD ;
reg  BAE ;
reg  BAF ;
reg  BAG ;
reg  BAH ;
reg  BAI ;
reg  BAJ ;
reg  BAK ;
reg  BAL ;
reg  BAM ;
reg  BAN ;
reg  BAO ;
reg  BAP ;
reg  BAQ ;
reg  BAR ;
reg  BAS ;
reg  BAT ;
reg  BAU ;
reg  BAV ;
reg  BAW ;
reg  BAX ;
reg  BBA ;
reg  BBB ;
reg  BBC ;
reg  BBD ;
reg  BBE ;
reg  BBF ;
reg  BBG ;
reg  BBH ;
reg  BBI ;
reg  BBJ ;
reg  BBK ;
reg  BBL ;
reg  BBM ;
reg  BBN ;
reg  BBO ;
reg  BBP ;
reg  BBQ ;
reg  BBR ;
reg  BBS ;
reg  BBT ;
reg  BBU ;
reg  BBV ;
reg  BBW ;
reg  BBX ;
reg  BCA ;
reg  BCB ;
reg  BCC ;
reg  BCD ;
reg  BCE ;
reg  BCF ;
reg  BCG ;
reg  BCH ;
reg  BCI ;
reg  BCJ ;
reg  BCK ;
reg  BCL ;
reg  BCM ;
reg  BCN ;
reg  BCO ;
reg  BCP ;
reg  BCQ ;
reg  BCR ;
reg  BCS ;
reg  BCT ;
reg  BCU ;
reg  BCV ;
reg  BCW ;
reg  BCX ;
reg  BDA ;
reg  BDB ;
reg  BDC ;
reg  BDD ;
reg  BDE ;
reg  BDF ;
reg  BDG ;
reg  BDH ;
reg  BDI ;
reg  BDJ ;
reg  BDK ;
reg  BDL ;
reg  BDM ;
reg  BDN ;
reg  BDO ;
reg  BDP ;
reg  BDQ ;
reg  BDR ;
reg  BDS ;
reg  BDT ;
reg  BDU ;
reg  BDV ;
reg  BDW ;
reg  BDX ;
reg  CAA ;
reg  CAB ;
reg  CAC ;
reg  CAD ;
reg  CAE ;
reg  CAF ;
reg  CAG ;
reg  CAH ;
reg  CAI ;
reg  CAJ ;
reg  CAK ;
reg  CAL ;
reg  CAM ;
reg  CAN ;
reg  CAO ;
reg  CAP ;
reg  CBA ;
reg  CBB ;
reg  CBC ;
reg  CBD ;
reg  CBE ;
reg  CBF ;
reg  CBG ;
reg  CBH ;
reg  CBI ;
reg  CBJ ;
reg  CBK ;
reg  CBL ;
reg  CBM ;
reg  CBN ;
reg  CBO ;
reg  CBP ;
reg  CCA ;
reg  CCB ;
reg  CCC ;
reg  CCD ;
reg  CCE ;
reg  CCF ;
reg  CCG ;
reg  CCH ;
reg  CCI ;
reg  CCJ ;
reg  CCK ;
reg  CCL ;
reg  CCM ;
reg  CCN ;
reg  CCO ;
reg  CCP ;
reg  CDA ;
reg  CDB ;
reg  CDC ;
reg  CDD ;
reg  CDE ;
reg  CDF ;
reg  CDG ;
reg  CDH ;
reg  CDI ;
reg  CDJ ;
reg  CDK ;
reg  CDL ;
reg  CDM ;
reg  CDN ;
reg  CDO ;
reg  CDP ;
reg  CEA ;
reg  CEB ;
reg  CEC ;
reg  CED ;
reg  CEE ;
reg  CEF ;
reg  CEG ;
reg  CEH ;
reg  CEI ;
reg  CEJ ;
reg  CEK ;
reg  CEL ;
reg  CEM ;
reg  CEN ;
reg  CEO ;
reg  CEP ;
reg  CFA ;
reg  CFB ;
reg  CFC ;
reg  CFD ;
reg  CFE ;
reg  CFF ;
reg  CFG ;
reg  CFH ;
reg  CFI ;
reg  CFJ ;
reg  CFK ;
reg  CFL ;
reg  CFM ;
reg  CFN ;
reg  CFO ;
reg  CFP ;
reg  CGA ;
reg  CGB ;
reg  CGC ;
reg  CGD ;
reg  CGE ;
reg  CGF ;
reg  CGG ;
reg  CGH ;
reg  CGI ;
reg  CGJ ;
reg  CGK ;
reg  CGL ;
reg  CGM ;
reg  CGN ;
reg  CGO ;
reg  CGP ;
reg  CHA ;
reg  CHB ;
reg  CHC ;
reg  CHD ;
reg  CHE ;
reg  CHF ;
reg  CHG ;
reg  CHH ;
reg  CHI ;
reg  CHJ ;
reg  CHK ;
reg  CHL ;
reg  CHM ;
reg  CHN ;
reg  CHO ;
reg  CHP ;
reg  CIA ;
reg  CIB ;
reg  CIC ;
reg  CID ;
reg  CIE ;
reg  CIF ;
reg  CIG ;
reg  CIH ;
reg  DAA ;
reg  DAB ;
reg  DAC ;
reg  DAD ;
reg  DAE ;
reg  DAF ;
reg  DAG ;
reg  DAH ;
reg  DBA ;
reg  DBB ;
reg  DBC ;
reg  DBD ;
reg  DBE ;
reg  DBF ;
reg  DBG ;
reg  DBH ;
reg  DCA ;
reg  DCB ;
reg  DCC ;
reg  DCD ;
reg  DCE ;
reg  DCF ;
reg  DCG ;
reg  DCH ;
reg  DDA ;
reg  DDB ;
reg  DDC ;
reg  DDD ;
reg  DDE ;
reg  DDF ;
reg  DDG ;
reg  DDH ;
reg  DEA ;
reg  DEB ;
reg  DEC ;
reg  DED ;
reg  DEE ;
reg  DEF ;
reg  DEG ;
reg  DEH ;
reg  DFA ;
reg  DFB ;
reg  DFC ;
reg  DFD ;
reg  DFE ;
reg  DFF ;
reg  DFG ;
reg  DFH ;
reg  DGA ;
reg  DGB ;
reg  DGC ;
reg  DGD ;
reg  DGE ;
reg  DGF ;
reg  DGG ;
reg  DGH ;
reg  DHA ;
reg  DHB ;
reg  DHC ;
reg  DHD ;
reg  DHE ;
reg  DHF ;
reg  DHG ;
reg  DHH ;
reg  DIA ;
reg  DIB ;
reg  DIC ;
reg  DID ;
reg  DIE ;
reg  DIF ;
reg  DIG ;
reg  DIH ;
reg  DJA ;
reg  DJB ;
reg  DJC ;
reg  DJD ;
reg  DJE ;
reg  DKA ;
reg  DKB ;
reg  DKC ;
reg  DKD ;
reg  DKE ;
reg  DLA ;
reg  DLB ;
reg  DLC ;
reg  DLD ;
reg  DLE ;
reg  DMA ;
reg  DMB ;
reg  DMC ;
reg  DMD ;
reg  DME ;
reg  DNA ;
reg  DNB ;
reg  DNC ;
reg  DND ;
reg  DNE ;
reg  DOA ;
reg  DOB ;
reg  DOC ;
reg  DOD ;
reg  DOE ;
reg  DPA ;
reg  DPB ;
reg  DPC ;
reg  DPD ;
reg  DPE ;
reg  DQA ;
reg  DQB ;
reg  DQC ;
reg  DQD ;
reg  DQE ;
reg  EAA ;
reg  EAB ;
reg  EAC ;
reg  EAD ;
reg  EAE ;
reg  EAF ;
reg  EAG ;
reg  EAH ;
reg  EBA ;
reg  EBB ;
reg  EBC ;
reg  EBD ;
reg  EBE ;
reg  EBF ;
reg  EBG ;
reg  EBH ;
reg  ECA ;
reg  ECB ;
reg  ECC ;
reg  ECD ;
reg  ECE ;
reg  ECF ;
reg  ECG ;
reg  ECH ;
reg  EDA ;
reg  EDB ;
reg  EDC ;
reg  EDD ;
reg  EDE ;
reg  EDF ;
reg  EDG ;
reg  EDH ;
reg  EEA ;
reg  EEB ;
reg  EEC ;
reg  EED ;
reg  EEE ;
reg  EEF ;
reg  EEG ;
reg  EEH ;
reg  EFA ;
reg  EFB ;
reg  EFC ;
reg  EFD ;
reg  EFE ;
reg  EFF ;
reg  EFG ;
reg  EFH ;
reg  EGA ;
reg  EGB ;
reg  EGC ;
reg  EGD ;
reg  EGE ;
reg  EGF ;
reg  EGG ;
reg  EGH ;
reg  EHA ;
reg  EHB ;
reg  EHC ;
reg  EHD ;
reg  EHE ;
reg  EHF ;
reg  EHG ;
reg  EHH ;
reg  EIA ;
reg  EIB ;
reg  EIC ;
reg  EID ;
reg  EIE ;
reg  EIF ;
reg  EIG ;
reg  EIH ;
reg  EJA ;
reg  EJB ;
reg  EJC ;
reg  EJD ;
reg  EJE ;
reg  EJF ;
reg  EJG ;
reg  EJH ;
reg  EKA ;
reg  EKB ;
reg  EKC ;
reg  EKD ;
reg  EKE ;
reg  EKF ;
reg  EKG ;
reg  EKH ;
reg  HAA ;
reg  HAB ;
reg  HAC ;
reg  HAD ;
reg  HAE ;
reg  HAF ;
reg  HAG ;
reg  HAH ;
reg  HBA ;
reg  HBB ;
reg  HBC ;
reg  HBD ;
reg  HBE ;
reg  HBF ;
reg  HBG ;
reg  HBH ;
reg  jja ;
reg  jjb ;
reg  LAA ;
reg  LAB ;
reg  LAC ;
reg  lba ;
reg  lbb ;
reg  lbc ;
reg  NAA ;
reg  NAB ;
reg  NAC ;
reg  NAD ;
reg  NAE ;
reg  NAF ;
reg  NBA ;
reg  NBB ;
reg  NBC ;
reg  NBD ;
reg  NBE ;
reg  NBF ;
reg  NCA ;
reg  NCB ;
reg  NCC ;
reg  NCD ;
reg  NCE ;
reg  NCF ;
reg  NDA ;
reg  NDB ;
reg  NDC ;
reg  NDD ;
reg  NDE ;
reg  NDF ;
reg  NEA ;
reg  NEB ;
reg  NEC ;
reg  NED ;
reg  NEE ;
reg  NEF ;
reg  NFA ;
reg  NFB ;
reg  NFC ;
reg  NFD ;
reg  NFE ;
reg  NFF ;
reg  NGA ;
reg  NGB ;
reg  NGC ;
reg  NGD ;
reg  NGE ;
reg  NGF ;
reg  NHA ;
reg  NHB ;
reg  NHC ;
reg  NHD ;
reg  NHE ;
reg  NHF ;
reg  NIA ;
reg  NIB ;
reg  NIC ;
reg  NID ;
reg  NIE ;
reg  NIF ;
reg  NJA ;
reg  NJB ;
reg  NJC ;
reg  NJD ;
reg  NJE ;
reg  NJF ;
reg  NKA ;
reg  NKB ;
reg  NKC ;
reg  NKD ;
reg  NKE ;
reg  NKF ;
reg  NLA ;
reg  NLB ;
reg  NLC ;
reg  NLD ;
reg  NLE ;
reg  NLF ;
reg  NMA ;
reg  NMB ;
reg  NMC ;
reg  NMD ;
reg  NME ;
reg  NMF ;
reg  NNA ;
reg  NNB ;
reg  NNC ;
reg  NND ;
reg  NNE ;
reg  NNF ;
reg  NOA ;
reg  NOB ;
reg  NOC ;
reg  NOD ;
reg  NOE ;
reg  NOF ;
reg  NPA ;
reg  NPB ;
reg  NPC ;
reg  NPD ;
reg  NPE ;
reg  NPF ;
reg  NQA ;
reg  NQB ;
reg  NQC ;
reg  NQD ;
reg  NQE ;
reg  NQF ;
reg  NRA ;
reg  NRB ;
reg  NRC ;
reg  NRD ;
reg  NRE ;
reg  NRF ;
reg  NSA ;
reg  NSB ;
reg  NSC ;
reg  NSD ;
reg  NSE ;
reg  NSF ;
reg  OAA ;
reg  OAB ;
reg  OAC ;
reg  OAD ;
reg  OAE ;
reg  OAF ;
reg  OAG ;
reg  OAH ;
reg  OAI ;
reg  OAJ ;
reg  OAK ;
reg  OAL ;
reg  OAM ;
reg  OAN ;
reg  OAO ;
reg  OAP ;
reg  OBA ;
reg  OBB ;
reg  OBC ;
reg  OBD ;
reg  OBE ;
reg  OBF ;
reg  OBG ;
reg  OBH ;
reg  OBI ;
reg  OBJ ;
reg  OBK ;
reg  OBL ;
reg  OBM ;
reg  OBN ;
reg  OBO ;
reg  OBP ;
reg  OCA ;
reg  OCB ;
reg  OCC ;
reg  OCD ;
reg  OCE ;
reg  OCF ;
reg  OCG ;
reg  OCH ;
reg  OCI ;
reg  OCJ ;
reg  OCK ;
reg  OCL ;
reg  OCM ;
reg  OCN ;
reg  OCO ;
reg  OCP ;
reg  ODA ;
reg  ODB ;
reg  ODC ;
reg  ODD ;
reg  ODE ;
reg  ODF ;
reg  ODG ;
reg  ODH ;
reg  ODI ;
reg  ODJ ;
reg  ODK ;
reg  ODL ;
reg  ODM ;
reg  ODN ;
reg  ODO ;
reg  ODP ;
reg  OEA ;
reg  OEB ;
reg  OEC ;
reg  OED ;
reg  OEE ;
reg  OEF ;
reg  OEG ;
reg  OEH ;
reg  OEI ;
reg  OEJ ;
reg  OEK ;
reg  OEL ;
reg  OEM ;
reg  OEN ;
reg  OEO ;
reg  OEP ;
reg  OFA ;
reg  OFB ;
reg  OFC ;
reg  OFD ;
reg  OFE ;
reg  OFF ;
reg  OFG ;
reg  OFH ;
reg  OFI ;
reg  OFJ ;
reg  OFK ;
reg  OFL ;
reg  OFM ;
reg  OFN ;
reg  OFO ;
reg  OFP ;
reg  OGA ;
reg  OGB ;
reg  OGC ;
reg  OGD ;
reg  OGE ;
reg  OGF ;
reg  OGG ;
reg  OGH ;
reg  OGI ;
reg  OGJ ;
reg  OGK ;
reg  OGL ;
reg  OGM ;
reg  OGN ;
reg  OGO ;
reg  OGP ;
reg  OHA ;
reg  OHB ;
reg  OHC ;
reg  OHD ;
reg  OHE ;
reg  OHF ;
reg  OHG ;
reg  OHH ;
reg  OHI ;
reg  OHJ ;
reg  OHK ;
reg  OHL ;
reg  OHM ;
reg  OHN ;
reg  OHO ;
reg  OHP ;
reg  OIA ;
reg  OIB ;
reg  OIC ;
reg  OID ;
reg  OIE ;
reg  OIF ;
reg  OIG ;
reg  OIH ;
reg  OJA ;
reg  ojb ;
reg  OKA ;
reg  OKB ;
reg  OKC ;
reg  OKD ;
reg  OKE ;
reg  OLA ;
reg  OLB ;
reg  OLC ;
reg  OLD ;
reg  OLE ;
reg  OMA ;
reg  OMB ;
reg  OMC ;
reg  OMD ;
reg  ONA ;
reg  ONB ;
reg  ONC ;
reg  OOA ;
reg  OOB ;
reg  OOC ;
reg  OPA ;
reg  PAD ;
reg  PAE ;
reg  PAF ;
reg  PCA ;
reg  PCB ;
reg  PCC ;
reg  PSD ;
reg  PSE ;
reg  PSF ;
reg  QAA ;
reg  QAB ;
reg  QAC ;
reg  QAD ;
reg  TAA ;
reg  TAB ;
reg  TAC ;
reg  TAD ;
reg  TAE ;
reg  TAF ;
reg  TAG ;
reg  TAH ;
reg  TAI ;
reg  TBA ;
reg  TBB ;
reg  TBC ;
reg  TBD ;
reg  TBE ;
reg  TBF ;
reg  TBG ;
reg  TBH ;
reg  TBI ;
reg  TCA ;
reg  TCB ;
reg  TCC ;
reg  TCD ;
reg  TCE ;
reg  TCF ;
reg  TCG ;
reg  TCH ;
reg  TCI ;
reg  TDA ;
reg  TDB ;
reg  TDC ;
reg  TDD ;
reg  TDE ;
reg  TDF ;
reg  TDG ;
reg  TDH ;
reg  TDI ;
wire  AAA ;
wire  AAB ;
wire  AAC ;
wire  AAD ;
wire  AAE ;
wire  AAF ;
wire  AAG ;
wire  AAH ;
wire  AAI ;
wire  AAJ ;
wire  AAK ;
wire  AAL ;
wire  AAM ;
wire  AAN ;
wire  AAO ;
wire  AAP ;
wire  AAQ ;
wire  AAR ;
wire  AAS ;
wire  AAT ;
wire  AAU ;
wire  AAV ;
wire  AAW ;
wire  AAX ;
wire  ABA ;
wire  ABB ;
wire  ABC ;
wire  ABD ;
wire  ABE ;
wire  ABF ;
wire  ABG ;
wire  ABH ;
wire  ABI ;
wire  ABJ ;
wire  ABK ;
wire  ABL ;
wire  ABM ;
wire  ABN ;
wire  ABO ;
wire  ABP ;
wire  ABQ ;
wire  ABR ;
wire  ABS ;
wire  ABT ;
wire  ABU ;
wire  ABV ;
wire  ABW ;
wire  ABX ;
wire  ACA ;
wire  ACB ;
wire  ACC ;
wire  ACD ;
wire  ACE ;
wire  ACF ;
wire  ACG ;
wire  ACH ;
wire  ACI ;
wire  ACJ ;
wire  ACK ;
wire  ACL ;
wire  ACM ;
wire  ACN ;
wire  ACO ;
wire  ACP ;
wire  ACQ ;
wire  ACR ;
wire  ACS ;
wire  ACT ;
wire  ACU ;
wire  ACV ;
wire  ACW ;
wire  ACX ;
wire  ADA ;
wire  ADB ;
wire  ADC ;
wire  ADD ;
wire  ADE ;
wire  ADF ;
wire  ADG ;
wire  ADH ;
wire  ADI ;
wire  ADJ ;
wire  ADK ;
wire  ADL ;
wire  ADM ;
wire  ADN ;
wire  ADO ;
wire  ADP ;
wire  ADQ ;
wire  ADR ;
wire  ADS ;
wire  ADT ;
wire  ADU ;
wire  ADV ;
wire  ADW ;
wire  ADX ;
wire  baa ;
wire  bab ;
wire  bac ;
wire  bad ;
wire  bae ;
wire  baf ;
wire  bag ;
wire  bah ;
wire  bai ;
wire  baj ;
wire  bak ;
wire  bal ;
wire  bam ;
wire  ban ;
wire  bao ;
wire  bap ;
wire  baq ;
wire  bar ;
wire  bas ;
wire  bat ;
wire  bau ;
wire  bav ;
wire  baw ;
wire  bax ;
wire  bba ;
wire  bbb ;
wire  bbc ;
wire  bbd ;
wire  bbe ;
wire  bbf ;
wire  bbg ;
wire  bbh ;
wire  bbi ;
wire  bbj ;
wire  bbk ;
wire  bbl ;
wire  bbm ;
wire  bbn ;
wire  bbo ;
wire  bbp ;
wire  bbq ;
wire  bbr ;
wire  bbs ;
wire  bbt ;
wire  bbu ;
wire  bbv ;
wire  bbw ;
wire  bbx ;
wire  bca ;
wire  bcb ;
wire  bcc ;
wire  bcd ;
wire  bce ;
wire  bcf ;
wire  bcg ;
wire  bch ;
wire  bci ;
wire  bcj ;
wire  bck ;
wire  bcl ;
wire  bcm ;
wire  bcn ;
wire  bco ;
wire  bcp ;
wire  bcq ;
wire  bcr ;
wire  bcs ;
wire  bct ;
wire  bcu ;
wire  bcv ;
wire  bcw ;
wire  bcx ;
wire  bda ;
wire  bdb ;
wire  bdc ;
wire  bdd ;
wire  bde ;
wire  bdf ;
wire  bdg ;
wire  bdh ;
wire  bdi ;
wire  bdj ;
wire  bdk ;
wire  bdl ;
wire  bdm ;
wire  bdn ;
wire  bdo ;
wire  bdp ;
wire  bdq ;
wire  bdr ;
wire  bds ;
wire  bdt ;
wire  bdu ;
wire  bdv ;
wire  bdw ;
wire  bdx ;
wire  caa ;
wire  cab ;
wire  cac ;
wire  cad ;
wire  cae ;
wire  caf ;
wire  cag ;
wire  cah ;
wire  cai ;
wire  caj ;
wire  cak ;
wire  cal ;
wire  cam ;
wire  can ;
wire  cao ;
wire  cap ;
wire  cba ;
wire  cbb ;
wire  cbc ;
wire  cbd ;
wire  cbe ;
wire  cbf ;
wire  cbg ;
wire  cbh ;
wire  cbi ;
wire  cbj ;
wire  cbk ;
wire  cbl ;
wire  cbm ;
wire  cbn ;
wire  cbo ;
wire  cbp ;
wire  cca ;
wire  ccb ;
wire  ccc ;
wire  ccd ;
wire  cce ;
wire  ccf ;
wire  ccg ;
wire  cch ;
wire  cci ;
wire  ccj ;
wire  cck ;
wire  ccl ;
wire  ccm ;
wire  ccn ;
wire  cco ;
wire  ccp ;
wire  cda ;
wire  cdb ;
wire  cdc ;
wire  cdd ;
wire  cde ;
wire  cdf ;
wire  cdg ;
wire  cdh ;
wire  cdi ;
wire  cdj ;
wire  cdk ;
wire  cdl ;
wire  cdm ;
wire  cdn ;
wire  cdo ;
wire  cdp ;
wire  cea ;
wire  ceb ;
wire  cec ;
wire  ced ;
wire  cee ;
wire  cef ;
wire  ceg ;
wire  ceh ;
wire  cei ;
wire  cej ;
wire  cek ;
wire  cel ;
wire  cem ;
wire  cen ;
wire  ceo ;
wire  cep ;
wire  cfa ;
wire  cfb ;
wire  cfc ;
wire  cfd ;
wire  cfe ;
wire  cff ;
wire  cfg ;
wire  cfh ;
wire  cfi ;
wire  cfj ;
wire  cfk ;
wire  cfl ;
wire  cfm ;
wire  cfn ;
wire  cfo ;
wire  cfp ;
wire  cga ;
wire  cgb ;
wire  cgc ;
wire  cgd ;
wire  cge ;
wire  cgf ;
wire  cgg ;
wire  cgh ;
wire  cgi ;
wire  cgj ;
wire  cgk ;
wire  cgl ;
wire  cgm ;
wire  cgn ;
wire  cgo ;
wire  cgp ;
wire  cha ;
wire  chb ;
wire  chc ;
wire  chd ;
wire  che ;
wire  chf ;
wire  chg ;
wire  chh ;
wire  chi ;
wire  chj ;
wire  chk ;
wire  chl ;
wire  chm ;
wire  chn ;
wire  cho ;
wire  chp ;
wire  cia ;
wire  cib ;
wire  cic ;
wire  cid ;
wire  cie ;
wire  cif ;
wire  cig ;
wire  cih ;
wire  daa ;
wire  dab ;
wire  dac ;
wire  dad ;
wire  dae ;
wire  daf ;
wire  dag ;
wire  dah ;
wire  dba ;
wire  dbb ;
wire  dbc ;
wire  dbd ;
wire  dbe ;
wire  dbf ;
wire  dbg ;
wire  dbh ;
wire  dca ;
wire  dcb ;
wire  dcc ;
wire  dcd ;
wire  dce ;
wire  dcf ;
wire  dcg ;
wire  dch ;
wire  dda ;
wire  ddb ;
wire  ddc ;
wire  ddd ;
wire  dde ;
wire  ddf ;
wire  ddg ;
wire  ddh ;
wire  dea ;
wire  deb ;
wire  dec ;
wire  ded ;
wire  dee ;
wire  def ;
wire  deg ;
wire  deh ;
wire  dfa ;
wire  dfb ;
wire  dfc ;
wire  dfd ;
wire  dfe ;
wire  dff ;
wire  dfg ;
wire  dfh ;
wire  dga ;
wire  dgb ;
wire  dgc ;
wire  dgd ;
wire  dge ;
wire  dgf ;
wire  dgg ;
wire  dgh ;
wire  dha ;
wire  dhb ;
wire  dhc ;
wire  dhd ;
wire  dhe ;
wire  dhf ;
wire  dhg ;
wire  dhh ;
wire  dia ;
wire  dib ;
wire  dic ;
wire  did ;
wire  die ;
wire  dif ;
wire  dig ;
wire  dih ;
wire  dja ;
wire  djb ;
wire  djc ;
wire  djd ;
wire  dje ;
wire  dka ;
wire  dkb ;
wire  dkc ;
wire  dkd ;
wire  dke ;
wire  dla ;
wire  dlb ;
wire  dlc ;
wire  dld ;
wire  dle ;
wire  dma ;
wire  dmb ;
wire  dmc ;
wire  dmd ;
wire  dme ;
wire  dna ;
wire  dnb ;
wire  dnc ;
wire  dnd ;
wire  dne ;
wire  doa ;
wire  dob ;
wire  doc ;
wire  dod ;
wire  doe ;
wire  dpa ;
wire  dpb ;
wire  dpc ;
wire  dpd ;
wire  dpe ;
wire  dqa ;
wire  dqb ;
wire  dqc ;
wire  dqd ;
wire  dqe ;
wire  eaa ;
wire  eab ;
wire  eac ;
wire  ead ;
wire  eae ;
wire  eaf ;
wire  eag ;
wire  eah ;
wire  eba ;
wire  ebb ;
wire  ebc ;
wire  ebd ;
wire  ebe ;
wire  ebf ;
wire  ebg ;
wire  ebh ;
wire  eca ;
wire  ecb ;
wire  ecc ;
wire  ecd ;
wire  ece ;
wire  ecf ;
wire  ecg ;
wire  ech ;
wire  eda ;
wire  edb ;
wire  edc ;
wire  edd ;
wire  ede ;
wire  edf ;
wire  edg ;
wire  edh ;
wire  eea ;
wire  eeb ;
wire  eec ;
wire  eed ;
wire  eee ;
wire  eef ;
wire  eeg ;
wire  eeh ;
wire  efa ;
wire  efb ;
wire  efc ;
wire  efd ;
wire  efe ;
wire  eff ;
wire  efg ;
wire  efh ;
wire  ega ;
wire  egb ;
wire  egc ;
wire  egd ;
wire  ege ;
wire  egf ;
wire  egg ;
wire  egh ;
wire  eha ;
wire  ehb ;
wire  ehc ;
wire  ehd ;
wire  ehe ;
wire  ehf ;
wire  ehg ;
wire  ehh ;
wire  eia ;
wire  eib ;
wire  eic ;
wire  eid ;
wire  eie ;
wire  eif ;
wire  eig ;
wire  eih ;
wire  eja ;
wire  ejb ;
wire  ejc ;
wire  ejd ;
wire  eje ;
wire  ejf ;
wire  ejg ;
wire  ejh ;
wire  eka ;
wire  ekb ;
wire  ekc ;
wire  ekd ;
wire  eke ;
wire  ekf ;
wire  ekg ;
wire  ekh ;
wire  faa ;
wire  FAA ;
wire  fab ;
wire  FAB ;
wire  fac ;
wire  FAC ;
wire  fad ;
wire  FAD ;
wire  fae ;
wire  FAE ;
wire  faf ;
wire  FAF ;
wire  fag ;
wire  FAG ;
wire  fah ;
wire  FAH ;
wire  fba ;
wire  FBA ;
wire  fbb ;
wire  FBB ;
wire  fbc ;
wire  FBC ;
wire  fbd ;
wire  FBD ;
wire  fbe ;
wire  FBE ;
wire  fbf ;
wire  FBF ;
wire  fbg ;
wire  FBG ;
wire  fbh ;
wire  FBH ;
wire  fca ;
wire  FCA ;
wire  fcb ;
wire  FCB ;
wire  fcc ;
wire  FCC ;
wire  fcd ;
wire  FCD ;
wire  fce ;
wire  FCE ;
wire  fcf ;
wire  FCF ;
wire  fcg ;
wire  FCG ;
wire  fch ;
wire  FCH ;
wire  gaa ;
wire  GAA ;
wire  gab ;
wire  GAB ;
wire  gac ;
wire  GAC ;
wire  gad ;
wire  GAD ;
wire  gae ;
wire  GAE ;
wire  gaf ;
wire  GAF ;
wire  gag ;
wire  GAG ;
wire  gah ;
wire  GAH ;
wire  gba ;
wire  GBA ;
wire  gbb ;
wire  GBB ;
wire  gbc ;
wire  GBC ;
wire  gbd ;
wire  GBD ;
wire  gbe ;
wire  GBE ;
wire  gbf ;
wire  GBF ;
wire  gbg ;
wire  GBG ;
wire  gbh ;
wire  GBH ;
wire  haa ;
wire  hab ;
wire  hac ;
wire  had ;
wire  hae ;
wire  haf ;
wire  hag ;
wire  hah ;
wire  hba ;
wire  hbb ;
wire  hbc ;
wire  hbd ;
wire  hbe ;
wire  hbf ;
wire  hbg ;
wire  hbh ;
wire  iaa ;
wire  iab ;
wire  iac ;
wire  iad ;
wire  iae ;
wire  iaf ;
wire  iag ;
wire  iah ;
wire  iai ;
wire  iaj ;
wire  iak ;
wire  ial ;
wire  iam ;
wire  ian ;
wire  iao ;
wire  iap ;
wire  iaq ;
wire  iar ;
wire  ias ;
wire  iat ;
wire  iau ;
wire  iav ;
wire  iaw ;
wire  iax ;
wire  iba ;
wire  ibb ;
wire  ibc ;
wire  ibd ;
wire  ibe ;
wire  ibf ;
wire  ibg ;
wire  ibh ;
wire  ibi ;
wire  ibj ;
wire  ibk ;
wire  ibl ;
wire  ibm ;
wire  ibn ;
wire  ibo ;
wire  ibp ;
wire  ibq ;
wire  ibr ;
wire  ibs ;
wire  ibt ;
wire  ibu ;
wire  ibv ;
wire  ibw ;
wire  ibx ;
wire  ica ;
wire  icb ;
wire  icc ;
wire  icd ;
wire  ice ;
wire  icf ;
wire  icg ;
wire  ich ;
wire  ici ;
wire  icj ;
wire  ick ;
wire  icl ;
wire  icm ;
wire  icn ;
wire  ico ;
wire  icp ;
wire  icq ;
wire  icr ;
wire  ics ;
wire  ict ;
wire  icu ;
wire  icv ;
wire  icw ;
wire  icx ;
wire  ida ;
wire  idb ;
wire  idc ;
wire  idd ;
wire  ide ;
wire  idf ;
wire  idg ;
wire  idh ;
wire  idi ;
wire  idj ;
wire  idk ;
wire  idl ;
wire  idm ;
wire  idn ;
wire  ido ;
wire  idp ;
wire  idq ;
wire  idr ;
wire  ids ;
wire  idt ;
wire  idu ;
wire  idv ;
wire  idw ;
wire  idx ;
wire  iea ;
wire  ieb ;
wire  iec ;
wire  ied ;
wire  iee ;
wire  ief ;
wire  ifa ;
wire  ifb ;
wire  ifc ;
wire  ifd ;
wire  ife ;
wire  ifff  ;
wire  iga ;
wire  igb ;
wire  igc ;
wire  igd ;
wire  ige ;
wire  igf ;
wire  iha ;
wire  ihb ;
wire  ihc ;
wire  ihd ;
wire  ihe ;
wire  ihf ;
wire  iia ;
wire  ija ;
wire  jaa ;
wire  JAA ;
wire  jab ;
wire  JAB ;
wire  jac ;
wire  JAC ;
wire  jad ;
wire  JAD ;
wire  jae ;
wire  JAE ;
wire  jaf ;
wire  JAF ;
wire  jag ;
wire  JAG ;
wire  jba ;
wire  JBA ;
wire  jbb ;
wire  JBB ;
wire  jbc ;
wire  JBC ;
wire  jbd ;
wire  JBD ;
wire  jbe ;
wire  JBE ;
wire  jbf ;
wire  JBF ;
wire  jbg ;
wire  JBG ;
wire  jca ;
wire  JCA ;
wire  jcb ;
wire  JCB ;
wire  jcc ;
wire  JCC ;
wire  jcd ;
wire  JCD ;
wire  jce ;
wire  JCE ;
wire  jcf ;
wire  JCF ;
wire  jcg ;
wire  JCG ;
wire  jda ;
wire  JDA ;
wire  jdb ;
wire  JDB ;
wire  jdc ;
wire  JDC ;
wire  jdd ;
wire  JDD ;
wire  jde ;
wire  JDE ;
wire  jdf ;
wire  JDF ;
wire  jdg ;
wire  JDG ;
wire  jea ;
wire  JEA ;
wire  jeb ;
wire  JEB ;
wire  jec ;
wire  JEC ;
wire  jed ;
wire  JED ;
wire  jee ;
wire  JEE ;
wire  jef ;
wire  JEF ;
wire  jeg ;
wire  JEG ;
wire  jfa ;
wire  JFA ;
wire  jfb ;
wire  JFB ;
wire  jfc ;
wire  JFC ;
wire  jfd ;
wire  JFD ;
wire  jfe ;
wire  JFE ;
wire  jff ;
wire  JFF ;
wire  jfg ;
wire  JFG ;
wire  jga ;
wire  JGA ;
wire  jgb ;
wire  JGB ;
wire  jgc ;
wire  JGC ;
wire  jgd ;
wire  JGD ;
wire  jge ;
wire  JGE ;
wire  jgf ;
wire  JGF ;
wire  jgg ;
wire  JGG ;
wire  jha ;
wire  JHA ;
wire  jhb ;
wire  JHB ;
wire  jhc ;
wire  JHC ;
wire  jhd ;
wire  JHD ;
wire  jhe ;
wire  JHE ;
wire  jhf ;
wire  JHF ;
wire  jhg ;
wire  JHG ;
wire  jia ;
wire  JIA ;
wire  jib ;
wire  JIB ;
wire  jic ;
wire  JIC ;
wire  jid ;
wire  JID ;
wire  jie ;
wire  JIE ;
wire  JJA ;
wire  JJB ;
wire  jpa ;
wire  JPA ;
wire  jqa ;
wire  JQA ;
wire  jqb ;
wire  JQB ;
wire  jqc ;
wire  JQC ;
wire  jqd ;
wire  JQD ;
wire  kaa ;
wire  KAA ;
wire  kab ;
wire  KAB ;
wire  kac ;
wire  KAC ;
wire  KAD ;
wire  kad ;
wire  kba ;
wire  KBA ;
wire  kbb ;
wire  KBB ;
wire  kbc ;
wire  KBC ;
wire  KBD ;
wire  kbd ;
wire  kca ;
wire  KCA ;
wire  kcb ;
wire  KCB ;
wire  kcc ;
wire  KCC ;
wire  KCD ;
wire  kcd ;
wire  kda ;
wire  KDA ;
wire  kdb ;
wire  KDB ;
wire  kdc ;
wire  KDC ;
wire  KDD ;
wire  kdd ;
wire  kea ;
wire  KEA ;
wire  keb ;
wire  KEB ;
wire  kec ;
wire  KEC ;
wire  KED ;
wire  ked ;
wire  kfa ;
wire  KFA ;
wire  kfb ;
wire  KFB ;
wire  kfc ;
wire  KFC ;
wire  KFD ;
wire  kfd ;
wire  kga ;
wire  KGA ;
wire  kgb ;
wire  KGB ;
wire  kgc ;
wire  KGC ;
wire  KGD ;
wire  kgd ;
wire  kha ;
wire  KHA ;
wire  khb ;
wire  KHB ;
wire  khc ;
wire  KHC ;
wire  KHD ;
wire  khd ;
wire  laa ;
wire  lab ;
wire  lac ;
wire  LBA ;
wire  LBB ;
wire  LBC ;
wire  maa ;
wire  MAA ;
wire  mab ;
wire  MAB ;
wire  mac ;
wire  MAC ;
wire  naa ;
wire  nab ;
wire  nac ;
wire  nad ;
wire  nae ;
wire  naf ;
wire  nba ;
wire  nbb ;
wire  nbc ;
wire  nbd ;
wire  nbe ;
wire  nbf ;
wire  nca ;
wire  ncb ;
wire  ncc ;
wire  ncd ;
wire  nce ;
wire  ncf ;
wire  nda ;
wire  ndb ;
wire  ndc ;
wire  ndd ;
wire  nde ;
wire  ndf ;
wire  nea ;
wire  neb ;
wire  nec ;
wire  ned ;
wire  nee ;
wire  nef ;
wire  nfa ;
wire  nfb ;
wire  nfc ;
wire  nfd ;
wire  nfe ;
wire  nff ;
wire  nga ;
wire  ngb ;
wire  ngc ;
wire  ngd ;
wire  nge ;
wire  ngf ;
wire  nha ;
wire  nhb ;
wire  nhc ;
wire  nhd ;
wire  nhe ;
wire  nhf ;
wire  nia ;
wire  nib ;
wire  nic ;
wire  nid ;
wire  nie ;
wire  nif ;
wire  nja ;
wire  njb ;
wire  njc ;
wire  njd ;
wire  nje ;
wire  njf ;
wire  nka ;
wire  nkb ;
wire  nkc ;
wire  nkd ;
wire  nke ;
wire  nkf ;
wire  nla ;
wire  nlb ;
wire  nlc ;
wire  nld ;
wire  nle ;
wire  nlf ;
wire  nma ;
wire  nmb ;
wire  nmc ;
wire  nmd ;
wire  nme ;
wire  nmf ;
wire  nna ;
wire  nnb ;
wire  nnc ;
wire  nnd ;
wire  nne ;
wire  nnf ;
wire  noa ;
wire  nob ;
wire  noc ;
wire  nod ;
wire  noe ;
wire  nof ;
wire  npa ;
wire  npb ;
wire  npc ;
wire  npd ;
wire  npe ;
wire  npf ;
wire  nqa ;
wire  nqb ;
wire  nqc ;
wire  nqd ;
wire  nqe ;
wire  nqf ;
wire  nra ;
wire  nrb ;
wire  nrc ;
wire  nrd ;
wire  nre ;
wire  nrf ;
wire  nsa ;
wire  nsb ;
wire  nsc ;
wire  nsd ;
wire  nse ;
wire  nsf ;
wire  oaa ;
wire  oab ;
wire  oac ;
wire  oad ;
wire  oae ;
wire  oaf ;
wire  oag ;
wire  oah ;
wire  oai ;
wire  oaj ;
wire  oak ;
wire  oal ;
wire  oam ;
wire  oan ;
wire  oao ;
wire  oap ;
wire  oba ;
wire  obb ;
wire  obc ;
wire  obd ;
wire  obe ;
wire  obf ;
wire  obg ;
wire  obh ;
wire  obi ;
wire  obj ;
wire  obk ;
wire  obl ;
wire  obm ;
wire  obn ;
wire  obo ;
wire  obp ;
wire  oca ;
wire  ocb ;
wire  occ ;
wire  ocd ;
wire  oce ;
wire  ocf ;
wire  ocg ;
wire  och ;
wire  oci ;
wire  ocj ;
wire  ock ;
wire  ocl ;
wire  ocm ;
wire  ocn ;
wire  oco ;
wire  ocp ;
wire  oda ;
wire  odb ;
wire  odc ;
wire  odd ;
wire  ode ;
wire  odf ;
wire  odg ;
wire  odh ;
wire  odi ;
wire  odj ;
wire  odk ;
wire  odl ;
wire  odm ;
wire  odn ;
wire  odo ;
wire  odp ;
wire  oea ;
wire  oeb ;
wire  oec ;
wire  oed ;
wire  oee ;
wire  oef ;
wire  oeg ;
wire  oeh ;
wire  oei ;
wire  oej ;
wire  oek ;
wire  oel ;
wire  oem ;
wire  oen ;
wire  oeo ;
wire  oep ;
wire  ofa ;
wire  ofb ;
wire  ofc ;
wire  ofd ;
wire  ofe ;
wire  off ;
wire  ofg ;
wire  ofh ;
wire  ofi ;
wire  ofj ;
wire  ofk ;
wire  ofl ;
wire  ofm ;
wire  ofn ;
wire  ofo ;
wire  ofp ;
wire  oga ;
wire  ogb ;
wire  ogc ;
wire  ogd ;
wire  oge ;
wire  ogf ;
wire  ogg ;
wire  ogh ;
wire  ogi ;
wire  ogj ;
wire  ogk ;
wire  ogl ;
wire  ogm ;
wire  ogn ;
wire  ogo ;
wire  ogp ;
wire  oha ;
wire  ohb ;
wire  ohc ;
wire  ohd ;
wire  ohe ;
wire  ohf ;
wire  ohg ;
wire  ohh ;
wire  ohi ;
wire  ohj ;
wire  ohk ;
wire  ohl ;
wire  ohm ;
wire  ohn ;
wire  oho ;
wire  ohp ;
wire  oia ;
wire  oib ;
wire  oic ;
wire  oid ;
wire  oie ;
wire  oif ;
wire  oig ;
wire  oih ;
wire  oja ;
wire  OJB ;
wire  oka ;
wire  okb ;
wire  okc ;
wire  okd ;
wire  oke ;
wire  ola ;
wire  olb ;
wire  olc ;
wire  old ;
wire  ole ;
wire  oma ;
wire  omb ;
wire  omc ;
wire  omd ;
wire  ona ;
wire  onb ;
wire  onc ;
wire  ooa ;
wire  oob ;
wire  ooc ;
wire  opa ;
wire  pad ;
wire  pae ;
wire  paf ;
wire  pca ;
wire  pcb ;
wire  pcc ;
wire  psd ;
wire  pse ;
wire  psf ;
wire  qaa ;
wire  qab ;
wire  qac ;
wire  qad ;
wire  taa ;
wire  tab ;
wire  tac ;
wire  tad ;
wire  tae ;
wire  taf ;
wire  tag ;
wire  tah ;
wire  tai ;
wire  tba ;
wire  tbb ;
wire  tbc ;
wire  tbd ;
wire  tbe ;
wire  tbf ;
wire  tbg ;
wire  tbh ;
wire  tbi ;
wire  tca ;
wire  tcb ;
wire  tcc ;
wire  tcd ;
wire  tce ;
wire  tcf ;
wire  tcg ;
wire  tch ;
wire  tci ;
wire  tda ;
wire  tdb ;
wire  tdc ;
wire  tdd ;
wire  tde ;
wire  tdf ;
wire  tdg ;
wire  tdh ;
wire  tdi ;
wire  ZZI ;
wire  ZZO ;
assign ZZI = 1'b1;
assign ZZO = 1'b0;
assign baa = ~BAA;  //complement 
assign bba = ~BBA;  //complement 
assign bca = ~BCA;  //complement 
assign bda = ~BDA;  //complement 
assign bai = ~BAI;  //complement 
assign bbi = ~BBI;  //complement 
assign bci = ~BCI;  //complement 
assign bdi = ~BDI;  //complement 
assign ega = ~EGA;  //complement 
assign baq = ~BAQ;  //complement 
assign bbq = ~BBQ;  //complement 
assign bcq = ~BCQ;  //complement 
assign bdq = ~BDQ;  //complement 
assign nba = ~NBA;  //complement 
assign nca = ~NCA;  //complement 
assign nea = ~NEA;  //complement 
assign nda = ~NDA;  //complement 
assign nfa = ~NFA;  //complement 
assign nga = ~NGA;  //complement 
assign nha = ~NHA;  //complement 
assign nia = ~NIA;  //complement 
assign nja = ~NJA;  //complement 
assign nka = ~NKA;  //complement 
assign nla = ~NLA;  //complement 
assign nma = ~NMA;  //complement 
assign nna = ~NNA;  //complement 
assign noa = ~NOA;  //complement 
assign npa = ~NPA;  //complement 
assign nqa = ~NQA;  //complement 
assign daa = ~DAA;  //complement 
assign dba = ~DBA;  //complement 
assign eaa = ~EAA;  //complement 
assign eba = ~EBA;  //complement 
assign dca = ~DCA;  //complement 
assign dda = ~DDA;  //complement 
assign eca = ~ECA;  //complement 
assign eda = ~EDA;  //complement 
assign dea = ~DEA;  //complement 
assign dfa = ~DFA;  //complement 
assign eea = ~EEA;  //complement 
assign efa = ~EFA;  //complement 
assign dga = ~DGA;  //complement 
assign dha = ~DHA;  //complement 
assign eha = ~EHA;  //complement 
assign cda = ~CDA;  //complement 
assign cdi = ~CDI;  //complement 
assign JDA =  CDF & cdg & cdh  |  cdf & CDG & cdh  |  cdf & cdg & CDH  |  CDF & CDG & CDH  ; 
assign jda = ~JDA; //complement 
assign dma = ~DMA;  //complement 
assign cea = ~CEA;  //complement 
assign cei = ~CEI;  //complement 
assign JEA =  CEF & ceg & ceh  |  cef & CEG & ceh  |  cef & ceg & CEH  |  CEF & CEG & CEH  ; 
assign jea = ~JEA; //complement 
assign dna = ~DNA;  //complement 
assign cfa = ~CFA;  //complement 
assign cfi = ~CFI;  //complement 
assign JFA =  CFF & cfg & cfh  |  cff & CFG & cfh  |  cff & cfg & CFH  |  CFF & CFG & CFH  ; 
assign jfa = ~JFA; //complement 
assign doa = ~DOA;  //complement 
assign nra = ~NRA;  //complement 
assign nsa = ~NSA;  //complement 
assign KAA =  DJA & dka & dla  |  dja & DKA & dla  |  dja & dka & DLA  |  DJA & DKA & DLA  ; 
assign kaa = ~KAA; //complement 
assign caa = ~CAA;  //complement 
assign cai = ~CAI;  //complement 
assign JAA =  CAF & cag & cah  |  caf & CAG & cah  |  caf & cag & CAH  |  CAF & CAG & CAH  ; 
assign jaa = ~JAA; //complement 
assign dja = ~DJA;  //complement 
assign cba = ~CBA;  //complement 
assign cbi = ~CBI;  //complement 
assign JBA =  CBF & cbg & cbh  |  cbf & CBG & cbh  |  cbf & cbg & CBH  |  CBF & CBG & CBH  ; 
assign jba = ~JBA; //complement 
assign dka = ~DKA;  //complement 
assign cca = ~CCA;  //complement 
assign cci = ~CCI;  //complement 
assign JCA =  CCF & ccg & cch  |  ccf & CCG & cch  |  ccf & ccg & CCH  |  CCF & CCG & CCH  ; 
assign jca = ~JCA; //complement 
assign dla = ~DLA;  //complement 
assign oai = ~OAI;  //complement 
assign JGA =  CGF & cgg & cgh  |  cgf & CGG & cgh  |  cgf & cgg & CGH  |  CGF & CGG & CGH  ; 
assign jga = ~JGA; //complement 
assign cga = ~CGA;  //complement 
assign cgi = ~CGI;  //complement 
assign AAA = ~aaa;  //complement 
assign ABA = ~aba;  //complement 
assign ACA = ~aca;  //complement 
assign ADA = ~ada;  //complement 
assign JHA =  CHF & chg & chh  |  chf & CHG & chh  |  chf & chg & CHH  |  CHF & CHG & CHH  ; 
assign jha = ~JHA; //complement 
assign cha = ~CHA;  //complement 
assign chi = ~CHI;  //complement 
assign AAI = ~aai;  //complement 
assign ABI = ~abi;  //complement 
assign ACI = ~aci;  //complement 
assign ADI = ~adi;  //complement 
assign dpa = ~DPA;  //complement 
assign dqa = ~DQA;  //complement 
assign cia = ~CIA;  //complement 
assign AAQ = ~aaq;  //complement 
assign ABQ = ~abq;  //complement 
assign ACQ = ~acq;  //complement 
assign ADQ = ~adq;  //complement 
assign pcb = ~PCB;  //complement 
assign oma = ~OMA;  //complement 
assign naa = ~NAA;  //complement 
assign hba = ~HBA;  //complement 
assign oia = ~OIA;  //complement 
assign oka = ~OKA;  //complement 
assign ola = ~OLA;  //complement 
assign KAB =  DMA & dne & doe  |  dma & DNE & doe  |  dma & dne & DOE  |  DMA & DNE & DOE  ; 
assign kab = ~KAB; //complement 
assign KAC =  DPE & dia  |  dpe & DIA  ; 
assign kac = ~KAC; //complement 
assign KAD =  DPE & dia  |  dpe & DIA  ; 
assign kad = ~KAD;  //complement 
assign oaa = ~OAA;  //complement 
assign oea = ~OEA;  //complement 
assign oca = ~OCA;  //complement 
assign oga = ~OGA;  //complement 
assign eia = ~EIA;  //complement 
assign FAH =  EID & EIC & EIB & eia & jja  ; 
assign fah = ~FAH;  //complement  
assign fca =  eia  ; 
assign FCA = ~fca;  //complement 
assign oei = ~OEI;  //complement 
assign oci = ~OCI;  //complement 
assign ogi = ~OGI;  //complement 
assign eja = ~EJA;  //complement 
assign dia = ~DIA;  //complement 
assign FBH =  EJD & EJC & EJB & eja & jjb  ; 
assign fbh = ~FBH;  //complement  
assign oba = ~OBA;  //complement 
assign ofa = ~OFA;  //complement 
assign oda = ~ODA;  //complement 
assign oha = ~OHA;  //complement 
assign eka = ~EKA;  //complement 
assign GAA =  ekd & ekc & ekb & eka  ; 
assign gaa = ~GAA;  //complement  
assign GBA =  ekh & ekg & ekf & eke  ; 
assign gba = ~GBA;  //complement 
assign obi = ~OBI;  //complement 
assign ofi = ~OFI;  //complement 
assign odi = ~ODI;  //complement 
assign ohi = ~OHI;  //complement 
assign bab = ~BAB;  //complement 
assign bbb = ~BBB;  //complement 
assign bcb = ~BCB;  //complement 
assign bdb = ~BDB;  //complement 
assign baj = ~BAJ;  //complement 
assign bbj = ~BBJ;  //complement 
assign bcj = ~BCJ;  //complement 
assign bdj = ~BDJ;  //complement 
assign bar = ~BAR;  //complement 
assign bbr = ~BBR;  //complement 
assign bcr = ~BCR;  //complement 
assign bdr = ~BDR;  //complement 
assign ecb = ~ECB;  //complement 
assign edb = ~EDB;  //complement 
assign nbb = ~NBB;  //complement 
assign ncb = ~NCB;  //complement 
assign nfb = ~NFB;  //complement 
assign ngb = ~NGB;  //complement 
assign nhb = ~NHB;  //complement 
assign nib = ~NIB;  //complement 
assign njb = ~NJB;  //complement 
assign nkb = ~NKB;  //complement 
assign nlb = ~NLB;  //complement 
assign nmb = ~NMB;  //complement 
assign nnb = ~NNB;  //complement 
assign nob = ~NOB;  //complement 
assign npb = ~NPB;  //complement 
assign nqb = ~NQB;  //complement 
assign dab = ~DAB;  //complement 
assign dbb = ~DBB;  //complement 
assign eab = ~EAB;  //complement 
assign ebb = ~EBB;  //complement 
assign dcb = ~DCB;  //complement 
assign ddb = ~DDB;  //complement 
assign deb = ~DEB;  //complement 
assign dfb = ~DFB;  //complement 
assign eeb = ~EEB;  //complement 
assign efb = ~EFB;  //complement 
assign ndb = ~NDB;  //complement 
assign neb = ~NEB;  //complement 
assign haa = ~HAA;  //complement 
assign hab = ~HAB;  //complement 
assign dgb = ~DGB;  //complement 
assign dhb = ~DHB;  //complement 
assign egb = ~EGB;  //complement 
assign ehb = ~EHB;  //complement 
assign cdb = ~CDB;  //complement 
assign cdj = ~CDJ;  //complement 
assign JDB =  CDB & cdc & cde  |  cdb & CDC & cde  |  cdb & cdc & CDE  |  CDB & CDC & CDE  ; 
assign jdb = ~JDB; //complement 
assign dmb = ~DMB;  //complement 
assign ceb = ~CEB;  //complement 
assign cej = ~CEJ;  //complement 
assign JEB =  CEB & cec & cee  |  ceb & CEC & cee  |  ceb & cec & CEE  |  CEB & CEC & CEE  ; 
assign jeb = ~JEB; //complement 
assign ACK = ~ack;  //complement 
assign cfb = ~CFB;  //complement 
assign cfj = ~CFJ;  //complement 
assign JFB =  CFB & cfc & cfe  |  cfb & CFC & cfe  |  cfb & cfc & CFE  |  CFB & CFC & CFE  ; 
assign jfb = ~JFB; //complement 
assign dob = ~DOB;  //complement 
assign nrb = ~NRB;  //complement 
assign nsb = ~NSB;  //complement 
assign dnb = ~DNB;  //complement 
assign dkb = ~DKB;  //complement 
assign KBA =  DJB & dkb & dlb  |  djb & DKB & dlb  |  djb & dkb & DLB  |  DJB & DKB & DLB  ; 
assign kba = ~KBA; //complement 
assign cab = ~CAB;  //complement 
assign caj = ~CAJ;  //complement 
assign JAB =  CAB & cac & cae  |  cab & CAC & cae  |  cab & cac & CAE  |  CAB & CAC & CAE  ; 
assign jab = ~JAB; //complement 
assign djb = ~DJB;  //complement 
assign cbb = ~CBB;  //complement 
assign cbj = ~CBJ;  //complement 
assign JBB =  CBB & cbc & cbe  |  cbb & CBC & cbe  |  cbb & cbc & CBE  |  CBB & CBC & CBE  ; 
assign jbb = ~JBB; //complement 
assign ccb = ~CCB;  //complement 
assign ccj = ~CCJ;  //complement 
assign JCB =  CCB & ccc & cce  |  ccb & CCC & cce  |  ccb & ccc & CCE  |  CCB & CCC & CCE  ; 
assign jcb = ~JCB; //complement 
assign dlb = ~DLB;  //complement 
assign dqb = ~DQB;  //complement 
assign JGB =  CGB & cgc & cge  |  cgb & CGC & cge  |  cgb & cgc & CGE  |  CGB & CGC & CGE  ; 
assign jgb = ~JGB; //complement 
assign cgb = ~CGB;  //complement 
assign cgj = ~CGJ;  //complement 
assign AAB = ~aab;  //complement 
assign ABB = ~abb;  //complement 
assign ACB = ~acb;  //complement 
assign ADB = ~adb;  //complement 
assign KBB =  DMB & dne & doe  |  dmb & DNE & doe  |  dmb & dne & DOE  |  DMB & DNE & DOE  ; 
assign kbb = ~KBB; //complement 
assign JHB =  CHB & chc & che  |  chb & CHC & che  |  chb & chc & CHE  |  CHB & CHC & CHE  ; 
assign jhb = ~JHB; //complement 
assign chb = ~CHB;  //complement 
assign chj = ~CHJ;  //complement 
assign AAJ = ~aaj;  //complement 
assign ABJ = ~abj;  //complement 
assign ACJ = ~acj;  //complement 
assign ADJ = ~adj;  //complement 
assign dpb = ~DPB;  //complement 
assign ofj = ~OFJ;  //complement 
assign cib = ~CIB;  //complement 
assign AAR = ~aar;  //complement 
assign ABR = ~abr;  //complement 
assign ACR = ~acr;  //complement 
assign ADR = ~adr;  //complement 
assign omb = ~OMB;  //complement 
assign nab = ~NAB;  //complement 
assign hbb = ~HBB;  //complement 
assign oib = ~OIB;  //complement 
assign okb = ~OKB;  //complement 
assign olb = ~OLB;  //complement 
assign ohb = ~OHB;  //complement 
assign KBC =  DQE & dib  |  dqe & DIB  ; 
assign kbc = ~KBC; //complement 
assign KBC =  DQE & dib  |  dqe & DIB  ; 
assign kbd = ~KBD;  //complement 
assign oab = ~OAB;  //complement 
assign oeb = ~OEB;  //complement 
assign ocb = ~OCB;  //complement 
assign ogb = ~OGB;  //complement 
assign eib = ~EIB;  //complement 
assign FAG =  EID & EIC & eib & EIA & jja  ; 
assign fag = ~FAG;  //complement  
assign fcb =  eib  ; 
assign FCB = ~fcb;  //complement 
assign oaj = ~OAJ;  //complement 
assign oej = ~OEJ;  //complement 
assign ocj = ~OCJ;  //complement 
assign ogj = ~OGJ;  //complement 
assign ejb = ~EJB;  //complement 
assign dib = ~DIB;  //complement 
assign FBG =  EJD & EJC & ejb & EJA & jjb  ; 
assign fbg = ~FBG;  //complement  
assign obb = ~OBB;  //complement 
assign ofb = ~OFB;  //complement 
assign odb = ~ODB;  //complement 
assign ekb = ~EKB;  //complement 
assign GAB =  EKD & ekc & ekb & EKA  ; 
assign gab = ~GAB;  //complement  
assign GBB =  EKH & ekg & ekf & EKE  ; 
assign gbb = ~GBB;  //complement 
assign obj = ~OBJ;  //complement 
assign odj = ~ODJ;  //complement 
assign ohj = ~OHJ;  //complement 
assign bac = ~BAC;  //complement 
assign bbc = ~BBC;  //complement 
assign bcc = ~BCC;  //complement 
assign bdc = ~BDC;  //complement 
assign bak = ~BAK;  //complement 
assign bbk = ~BBK;  //complement 
assign bck = ~BCK;  //complement 
assign bdk = ~BDK;  //complement 
assign bds = ~BDS;  //complement 
assign bas = ~BAS;  //complement 
assign bat = ~BAT;  //complement 
assign bbs = ~BBS;  //complement 
assign bcs = ~BCS;  //complement 
assign nbc = ~NBC;  //complement 
assign ncc = ~NCC;  //complement 
assign nec = ~NEC;  //complement 
assign ndc = ~NDC;  //complement 
assign nfc = ~NFC;  //complement 
assign ngc = ~NGC;  //complement 
assign nhc = ~NHC;  //complement 
assign nic = ~NIC;  //complement 
assign njc = ~NJC;  //complement 
assign nkc = ~NKC;  //complement 
assign nlc = ~NLC;  //complement 
assign nmc = ~NMC;  //complement 
assign nnc = ~NNC;  //complement 
assign noc = ~NOC;  //complement 
assign npc = ~NPC;  //complement 
assign nqc = ~NQC;  //complement 
assign dac = ~DAC;  //complement 
assign dbc = ~DBC;  //complement 
assign dbd = ~DBD;  //complement 
assign eac = ~EAC;  //complement 
assign ead = ~EAD;  //complement 
assign ebc = ~EBC;  //complement 
assign ebd = ~EBD;  //complement 
assign dcd = ~DCD;  //complement 
assign ddc = ~DDC;  //complement 
assign ecc = ~ECC;  //complement 
assign edc = ~EDC;  //complement 
assign efc = ~EFC;  //complement 
assign efd = ~EFD;  //complement 
assign dec = ~DEC;  //complement 
assign dfc = ~DFC;  //complement 
assign dfd = ~DFD;  //complement 
assign eec = ~EEC;  //complement 
assign ehd = ~EHD;  //complement 
assign dcc = ~DCC;  //complement 
assign dgc = ~DGC;  //complement 
assign dhc = ~DHC;  //complement 
assign egc = ~EGC;  //complement 
assign ehc = ~EHC;  //complement 
assign cdc = ~CDC;  //complement 
assign cdk = ~CDK;  //complement 
assign dkc = ~DKC;  //complement 
assign JDC =  CDA & cdd  |  cda & CDD  |  cda & cdd  |  CDA & CDD  ; 
assign jdc = ~JDC; //complement 
assign dmc = ~DMC;  //complement 
assign cec = ~CEC;  //complement 
assign cek = ~CEK;  //complement 
assign JEC =  CEA & ced  |  cea & CED  |  cea & ced  |  CEA & CED  ; 
assign jec = ~JEC; //complement 
assign dnc = ~DNC;  //complement 
assign cfc = ~CFC;  //complement 
assign cfk = ~CFK;  //complement 
assign cfp = ~CFP;  //complement 
assign JFC =  CFA & cfd  |  cfa & CFD  |  cfa & cfd  |  CFA & CFD  ; 
assign jfc = ~JFC; //complement 
assign doc = ~DOC;  //complement 
assign nrc = ~NRC;  //complement 
assign nsc = ~NSC;  //complement 
assign tbc = ~TBC;  //complement 
assign KCA =  DJC & dkc & dlc  |  djc & DKC & dlc  |  djc & dkc & DLC  |  DJC & DKC & DLC  ; 
assign kca = ~KCA; //complement 
assign cac = ~CAC;  //complement 
assign cak = ~CAK;  //complement 
assign JAC =  CAA & cad  |  caa & CAD  |  caa & cad  |  CAA & CAD  ; 
assign jac = ~JAC; //complement 
assign djc = ~DJC;  //complement 
assign cbc = ~CBC;  //complement 
assign cbk = ~CBK;  //complement 
assign JBC =  CBA & cbd  |  cba & CBD  |  cba & cbd  |  CBA & CBD  ; 
assign jbc = ~JBC; //complement 
assign ccc = ~CCC;  //complement 
assign cck = ~CCK;  //complement 
assign JCC =  CCA & ccd  |  cca & CCD  |  cca & ccd  |  CCA & CCD  ; 
assign jcc = ~JCC; //complement 
assign dlc = ~DLC;  //complement 
assign ofk = ~OFK;  //complement 
assign JGC =  CGA & cgd  |  cga & CGD  |  cga & cgd  |  CGA & CGD  ; 
assign jgc = ~JGC; //complement 
assign cgc = ~CGC;  //complement 
assign cgk = ~CGK;  //complement 
assign AAC = ~aac;  //complement 
assign ACC = ~acc;  //complement 
assign ADC = ~adc;  //complement 
assign JHC =  CHA & chd  |  cha & CHD  |  cha & chd  |  CHA & CHD  ; 
assign jhc = ~JHC; //complement 
assign chc = ~CHC;  //complement 
assign chk = ~CHK;  //complement 
assign AAK = ~aak;  //complement 
assign ABK = ~abk;  //complement 
assign ADK = ~adk;  //complement 
assign dpc = ~DPC;  //complement 
assign dqc = ~DQC;  //complement 
assign cic = ~CIC;  //complement 
assign AAS = ~aas;  //complement 
assign ABS = ~abs;  //complement 
assign ACS = ~acs;  //complement 
assign ADS = ~ads;  //complement 
assign KCB =  DMC & dne & dqe  |  dmc & DNE & dqe  |  dmc & dne & DQE  |  DMC & DNE & DQE  ; 
assign kcb = ~KCB; //complement 
assign omc = ~OMC;  //complement 
assign nac = ~NAC;  //complement 
assign hbc = ~HBC;  //complement 
assign oic = ~OIC;  //complement 
assign okc = ~OKC;  //complement 
assign olc = ~OLC;  //complement 
assign ohc = ~OHC;  //complement 
assign KCC =  DPE & dic  |  dpe & DIC  ; 
assign kcc = ~KCC; //complement 
assign KCD =  DPE & dic  |  dpe & DIC  ; 
assign kcd = ~KCD;  //complement 
assign oac = ~OAC;  //complement 
assign oec = ~OEC;  //complement 
assign occ = ~OCC;  //complement 
assign ogc = ~OGC;  //complement 
assign eic = ~EIC;  //complement 
assign hac = ~HAC;  //complement 
assign FAF =  EID & eic & EIB & EIA & jja  ; 
assign faf = ~FAF;  //complement  
assign fcc =  eic  ; 
assign FCC = ~fcc;  //complement 
assign oak = ~OAK;  //complement 
assign oek = ~OEK;  //complement 
assign ock = ~OCK;  //complement 
assign ogk = ~OGK;  //complement 
assign ejc = ~EJC;  //complement 
assign dic = ~DIC;  //complement 
assign FBF =  EJD & ejc & EJB & EJA & jjb  ; 
assign fbf = ~FBF;  //complement  
assign obc = ~OBC;  //complement 
assign ofc = ~OFC;  //complement 
assign odc = ~ODC;  //complement 
assign ekc = ~EKC;  //complement 
assign GAC =  EKD & ekc & EKB & eka  ; 
assign gac = ~GAC;  //complement  
assign GBC =  EKH & ekg & EKF & eke  ; 
assign gbc = ~GBC;  //complement 
assign obk = ~OBK;  //complement 
assign odk = ~ODK;  //complement 
assign ohk = ~OHK;  //complement 
assign bad = ~BAD;  //complement 
assign bbd = ~BBD;  //complement 
assign bcd = ~BCD;  //complement 
assign bdd = ~BDD;  //complement 
assign bal = ~BAL;  //complement 
assign bbl = ~BBL;  //complement 
assign bcl = ~BCL;  //complement 
assign bdl = ~BDL;  //complement 
assign bbt = ~BBT;  //complement 
assign bct = ~BCT;  //complement 
assign bdt = ~BDT;  //complement 
assign nbd = ~NBD;  //complement 
assign ncd = ~NCD;  //complement 
assign ndd = ~NDD;  //complement 
assign ned = ~NED;  //complement 
assign nfd = ~NFD;  //complement 
assign ngd = ~NGD;  //complement 
assign nhd = ~NHD;  //complement 
assign nid = ~NID;  //complement 
assign njd = ~NJD;  //complement 
assign nkd = ~NKD;  //complement 
assign nld = ~NLD;  //complement 
assign nmd = ~NMD;  //complement 
assign nnd = ~NND;  //complement 
assign nod = ~NOD;  //complement 
assign npd = ~NPD;  //complement 
assign nqd = ~NQD;  //complement 
assign dad = ~DAD;  //complement 
assign ddd = ~DDD;  //complement 
assign ecd = ~ECD;  //complement 
assign edd = ~EDD;  //complement 
assign ded = ~DED;  //complement 
assign eed = ~EED;  //complement 
assign dgd = ~DGD;  //complement 
assign dhd = ~DHD;  //complement 
assign egd = ~EGD;  //complement 
assign cdd = ~CDD;  //complement 
assign cdl = ~CDL;  //complement 
assign JDD =  CDB & cdd & cdf  |  cdb & CDD & cdf  |  cdb & cdd & CDF  |  CDB & CDD & CDF  ; 
assign jdd = ~JDD; //complement 
assign dmd = ~DMD;  //complement 
assign ced = ~CED;  //complement 
assign cel = ~CEL;  //complement 
assign JED =  CEB & ced & cef  |  ceb & CED & cef  |  ceb & ced & CEF  |  CEB & CED & CEF  ; 
assign jed = ~JED; //complement 
assign dnd = ~DND;  //complement 
assign cfd = ~CFD;  //complement 
assign cfl = ~CFL;  //complement 
assign JFD =  CFB & cfd & cff  |  cfb & CFD & cff  |  cfb & cfd & CFF  |  CFB & CFD & CFF  ; 
assign jfd = ~JFD; //complement 
assign dod = ~DOD;  //complement 
assign nrd = ~NRD;  //complement 
assign nsd = ~NSD;  //complement 
assign psd = ~PSD;  //complement 
assign KDA =  DJD & dkd & dld  |  djd & DKD & dld  |  djd & dkd & DLD  |  DJD & DKD & DLD  ; 
assign kda = ~KDA; //complement 
assign cad = ~CAD;  //complement 
assign cal = ~CAL;  //complement 
assign JAD =  CAB & cad & caf  |  cab & CAD & caf  |  cab & cad & CAF  |  CAB & CAD & CAF  ; 
assign jad = ~JAD; //complement 
assign djd = ~DJD;  //complement 
assign cbd = ~CBD;  //complement 
assign cbl = ~CBL;  //complement 
assign JBD =  CBB & cbd & cbf  |  cbb & CBD & cbf  |  cbb & cbd & CBF  |  CBB & CBD & CBF  ; 
assign jbd = ~JBD; //complement 
assign dkd = ~DKD;  //complement 
assign ccd = ~CCD;  //complement 
assign ccl = ~CCL;  //complement 
assign JCD =  CCB & ccd & ccf  |  ccb & CCD & ccf  |  ccb & ccd & CCF  |  CCB & CCD & CCF  ; 
assign jcd = ~JCD; //complement 
assign dld = ~DLD;  //complement 
assign JGD =  CGB & cgd & cgf  |  cgb & CGD & cgf  |  cgb & cgd & CGF  |  CGB & CGD & CGF  ; 
assign jgd = ~JGD; //complement 
assign cgd = ~CGD;  //complement 
assign cgl = ~CGL;  //complement 
assign AAD = ~aad;  //complement 
assign ABD = ~abd;  //complement 
assign ACD = ~acd;  //complement 
assign ADD = ~add;  //complement 
assign JHD =  CHB & chd & chf  |  chb & CHD & chf  |  chb & chd & CHF  |  CHB & CHD & CHF  ; 
assign jhd = ~JHD; //complement 
assign chd = ~CHD;  //complement 
assign chl = ~CHL;  //complement 
assign AAL = ~aal;  //complement 
assign ABL = ~abl;  //complement 
assign ACL = ~acl;  //complement 
assign ADL = ~adl;  //complement 
assign dpd = ~DPD;  //complement 
assign dqd = ~DQD;  //complement 
assign cid = ~CID;  //complement 
assign AAT = ~aat;  //complement 
assign ABT = ~abt;  //complement 
assign ACT = ~act;  //complement 
assign ADT = ~adt;  //complement 
assign KDB =  DMD & doe & dpe  |  dmd & DOE & dpe  |  dmd & doe & DPE  |  DMD & DOE & DPE  ; 
assign kdb = ~KDB; //complement 
assign nad = ~NAD;  //complement 
assign pad = ~PAD;  //complement 
assign hbd = ~HBD;  //complement 
assign oid = ~OID;  //complement 
assign okd = ~OKD;  //complement 
assign old = ~OLD;  //complement 
assign ohd = ~OHD;  //complement 
assign KDC =  DQE & did  |  dqe & DID  ; 
assign kdc = ~KDC; //complement 
assign KDD =  DQE & did  |  dqe & DID  ; 
assign kdd = ~KDD;  //complement 
assign oad = ~OAD;  //complement 
assign oed = ~OED;  //complement 
assign ocd = ~OCD;  //complement 
assign ogd = ~OGD;  //complement 
assign eid = ~EID;  //complement 
assign had = ~HAD;  //complement 
assign FAE =  eid & EIC & EIB & EIA & jja  ; 
assign fae = ~FAE;  //complement  
assign fcd =  eid  ; 
assign FCD = ~fcd;  //complement 
assign oal = ~OAL;  //complement 
assign oel = ~OEL;  //complement 
assign ocl = ~OCL;  //complement 
assign ogl = ~OGL;  //complement 
assign ejd = ~EJD;  //complement 
assign did = ~DID;  //complement 
assign FBE =  ejd & EJC & EJB & EJA & jjb  ; 
assign fbe = ~FBE;  //complement  
assign obd = ~OBD;  //complement 
assign ofd = ~OFD;  //complement 
assign odd = ~ODD;  //complement 
assign ekd = ~EKD;  //complement 
assign GAD =  ekd & ekc & EKB & EKA  ; 
assign gad = ~GAD;  //complement  
assign GBD =  ekh & ekg & EKF & EKE  ; 
assign gbd = ~GBD;  //complement 
assign obl = ~OBL;  //complement 
assign ofl = ~OFL;  //complement 
assign odl = ~ODL;  //complement 
assign ohl = ~OHL;  //complement 
assign cdh = ~CDH;  //complement 
assign bae = ~BAE;  //complement 
assign bbe = ~BBE;  //complement 
assign bce = ~BCE;  //complement 
assign bde = ~BDE;  //complement 
assign cem = ~CEM;  //complement 
assign bam = ~BAM;  //complement 
assign bbm = ~BBM;  //complement 
assign bcm = ~BCM;  //complement 
assign bdm = ~BDM;  //complement 
assign bau = ~BAU;  //complement 
assign bbu = ~BBU;  //complement 
assign bcu = ~BCU;  //complement 
assign bdu = ~BDU;  //complement 
assign nbe = ~NBE;  //complement 
assign nce = ~NCE;  //complement 
assign nde = ~NDE;  //complement 
assign nee = ~NEE;  //complement 
assign nfe = ~NFE;  //complement 
assign nge = ~NGE;  //complement 
assign nhe = ~NHE;  //complement 
assign nie = ~NIE;  //complement 
assign nje = ~NJE;  //complement 
assign nke = ~NKE;  //complement 
assign nle = ~NLE;  //complement 
assign nme = ~NME;  //complement 
assign nne = ~NNE;  //complement 
assign noe = ~NOE;  //complement 
assign npe = ~NPE;  //complement 
assign nqe = ~NQE;  //complement 
assign dae = ~DAE;  //complement 
assign dbe = ~DBE;  //complement 
assign eae = ~EAE;  //complement 
assign ebe = ~EBE;  //complement 
assign dce = ~DCE;  //complement 
assign dde = ~DDE;  //complement 
assign ede = ~EDE;  //complement 
assign ece = ~ECE;  //complement 
assign dee = ~DEE;  //complement 
assign dfe = ~DFE;  //complement 
assign eee = ~EEE;  //complement 
assign efe = ~EFE;  //complement 
assign dge = ~DGE;  //complement 
assign dhe = ~DHE;  //complement 
assign ege = ~EGE;  //complement 
assign ehe = ~EHE;  //complement 
assign cde = ~CDE;  //complement 
assign cdm = ~CDM;  //complement 
assign JDE =  CDC & cdd & cdg  |  cdc & CDD & cdg  |  cdc & cdd & CDG  |  CDC & CDD & CDG  ; 
assign jde = ~JDE; //complement 
assign dme = ~DME;  //complement 
assign cee = ~CEE;  //complement 
assign JDG =  CDE  ; 
assign jdg = ~JDG;  //complement 
assign JEE =  CEC & ced & ceg  |  cec & CED & ceg  |  cec & ced & CEG  |  CEC & CED & CEG  ; 
assign jee = ~JEE; //complement 
assign dne = ~DNE;  //complement 
assign cfe = ~CFE;  //complement 
assign cfm = ~CFM;  //complement 
assign JEG =  CEE  ; 
assign jeg = ~JEG;  //complement 
assign JFE =  CFC & cfd & cfg  |  cfc & CFD & cfg  |  cfc & cfd & CFG  |  CFC & CFD & CFG  ; 
assign jfe = ~JFE; //complement 
assign JFG = CFE; 
assign jfg = ~JFG; 
assign doe = ~DOE;  //complement 
assign nre = ~NRE;  //complement 
assign nse = ~NSE;  //complement 
assign pse = ~PSE;  //complement 
assign JAG =  CAE  |  CAE  ; 
assign jag = ~JAG; //complement 
assign KEA =  DOA & dpa & dqa  |  doa & DPA & dqa  |  doa & dpa & DQA  |  DOA & DPA & DQA  ; 
assign kea = ~KEA; //complement 
assign pcc = ~PCC;  //complement 
assign cae = ~CAE;  //complement 
assign cam = ~CAM;  //complement 
assign JAE =  CAC & cad & cag  |  cac & CAD & cag  |  cac & cad & CAG  |  CAC & CAD & CAG  ; 
assign jae = ~JAE; //complement 
assign dje = ~DJE;  //complement 
assign cbe = ~CBE;  //complement 
assign cbm = ~CBM;  //complement 
assign JBE =  CBC & cbd & cbg  |  cbc & CBD & cbg  |  cbc & cbd & CBG  |  CBC & CBD & CBG  ; 
assign jbe = ~JBE; //complement 
assign JBG = CBE; 
assign jbg = ~JBG; 
assign dke = ~DKE;  //complement 
assign cce = ~CCE;  //complement 
assign ccm = ~CCM;  //complement 
assign JCE =  CCC & ccd & ccg  |  ccc & CCD & ccg  |  ccc & ccd & CCG  |  CCC & CCD & CCG  ; 
assign jce = ~JCE; //complement 
assign JCG = CCE; 
assign jcg = ~JCG; 
assign dle = ~DLE;  //complement 
assign JGE =  CGC & cgd & cgg  |  cgc & CGD & cgg  |  cgc & cgd & CGG  |  CGC & CGD & CGG  ; 
assign jge = ~JGE; //complement 
assign JGG = CGE; 
assign jgg = ~JGG; 
assign cge = ~CGE;  //complement 
assign cgm = ~CGM;  //complement 
assign AAE = ~aae;  //complement 
assign ABE = ~abe;  //complement 
assign ACE = ~ace;  //complement 
assign ADE = ~ade;  //complement 
assign KEB =  DNA & dke & dle  |  dna & DKE & dle  |  dna & dke & DLE  |  DNA & DKE & DLE  ; 
assign keb = ~KEB; //complement 
assign JHE =  CHC & chd & chg  |  chc & CHD & chg  |  chc & chd & CHG  |  CHC & CHD & CHG  ; 
assign jhe = ~JHE; //complement 
assign JHG = CHE; 
assign jhg = ~JHG; 
assign che = ~CHE;  //complement 
assign chm = ~CHM;  //complement 
assign AAM = ~aam;  //complement 
assign ABM = ~abm;  //complement 
assign ACM = ~acm;  //complement 
assign ADM = ~adm;  //complement 
assign dpe = ~DPE;  //complement 
assign dqe = ~DQE;  //complement 
assign cie = ~CIE;  //complement 
assign AAU = ~aau;  //complement 
assign ABU = ~abu;  //complement 
assign ACU = ~acu;  //complement 
assign ADU = ~adu;  //complement 
assign JIA =  paf & PAE & PAD  ; 
assign jia = ~JIA;  //complement 
assign JIB =  PSF & pse  ; 
assign jib = ~JIB;  //complement 
assign JIC =  PSF & PSE  ; 
assign jic = ~JIC;  //complement 
assign omd = ~OMD;  //complement 
assign nae = ~NAE;  //complement 
assign pae = ~PAE;  //complement 
assign hbe = ~HBE;  //complement 
assign oie = ~OIE;  //complement 
assign oke = ~OKE;  //complement 
assign ole = ~OLE;  //complement 
assign ode = ~ODE;  //complement 
assign KEC =  DJE & die  |  dje & DIE  ; 
assign kec = ~KEC; //complement 
assign KED =  DJE & die  |  dje & DIE  ; 
assign ked = ~KED;  //complement 
assign oae = ~OAE;  //complement 
assign oee = ~OEE;  //complement 
assign oce = ~OCE;  //complement 
assign oge = ~OGE;  //complement 
assign eie = ~EIE;  //complement 
assign hae = ~HAE;  //complement 
assign FAD =  EIH & EIG & EIF & eie & jja  ; 
assign fad = ~FAD;  //complement  
assign fce =  eie  ; 
assign FCE = ~fce;  //complement 
assign oam = ~OAM;  //complement 
assign oem = ~OEM;  //complement 
assign ocm = ~OCM;  //complement 
assign ogm = ~OGM;  //complement 
assign eje = ~EJE;  //complement 
assign die = ~DIE;  //complement 
assign FBD =  EJH & EJG & EJF & eje & jjb  ; 
assign fbd = ~FBD;  //complement  
assign obe = ~OBE;  //complement 
assign ofe = ~OFE;  //complement 
assign ohe = ~OHE;  //complement 
assign eke = ~EKE;  //complement 
assign GAE =  EKD & EKC & ekb & eka  ; 
assign gae = ~GAE;  //complement  
assign GBE =  EKH & EKG & ekf & eke  ; 
assign gbe = ~GBE;  //complement 
assign obm = ~OBM;  //complement 
assign ofm = ~OFM;  //complement 
assign odm = ~ODM;  //complement 
assign ohm = ~OHM;  //complement 
assign baf = ~BAF;  //complement 
assign bbf = ~BBF;  //complement 
assign bcf = ~BCF;  //complement 
assign bdf = ~BDF;  //complement 
assign dcf = ~DCF;  //complement 
assign ban = ~BAN;  //complement 
assign bbn = ~BBN;  //complement 
assign bcn = ~BCN;  //complement 
assign bdn = ~BDN;  //complement 
assign bav = ~BAV;  //complement 
assign bbv = ~BBV;  //complement 
assign bcv = ~BCV;  //complement 
assign bdv = ~BDV;  //complement 
assign nbf = ~NBF;  //complement 
assign ncf = ~NCF;  //complement 
assign ndf = ~NDF;  //complement 
assign nef = ~NEF;  //complement 
assign nff = ~NFF;  //complement 
assign ngf = ~NGF;  //complement 
assign nhf = ~NHF;  //complement 
assign nif = ~NIF;  //complement 
assign njf = ~NJF;  //complement 
assign nkf = ~NKF;  //complement 
assign nlf = ~NLF;  //complement 
assign nmf = ~NMF;  //complement 
assign nnf = ~NNF;  //complement 
assign nof = ~NOF;  //complement 
assign npf = ~NPF;  //complement 
assign nqf = ~NQF;  //complement 
assign daf = ~DAF;  //complement 
assign dbf = ~DBF;  //complement 
assign eaf = ~EAF;  //complement 
assign ebf = ~EBF;  //complement 
assign ddf = ~DDF;  //complement 
assign ecf = ~ECF;  //complement 
assign edf = ~EDF;  //complement 
assign def = ~DEF;  //complement 
assign dff = ~DFF;  //complement 
assign eef = ~EEF;  //complement 
assign eff = ~EFF;  //complement 
assign dgf = ~DGF;  //complement 
assign dhf = ~DHF;  //complement 
assign egf = ~EGF;  //complement 
assign ehf = ~EHF;  //complement 
assign cdf = ~CDF;  //complement 
assign cdn = ~CDN;  //complement 
assign cef = ~CEF;  //complement 
assign cen = ~CEN;  //complement 
assign cff = ~CFF;  //complement 
assign cfn = ~CFN;  //complement 
assign nrf = ~NRF;  //complement 
assign nsf = ~NSF;  //complement 
assign psf = ~PSF;  //complement 
assign KFA =  DOB & dpb & dqb  |  dob & DPB & dqb  |  dob & dpb & DQB  |  DOB & DPB & DQB  ; 
assign kfa = ~KFA; //complement 
assign caf = ~CAF;  //complement 
assign can = ~CAN;  //complement 
assign cbf = ~CBF;  //complement 
assign cbn = ~CBN;  //complement 
assign jqd =  jqa & jqb & jqc  ; 
assign JQD = ~jqd;  //complement 
assign jqa =  EJA & ejb & eje  |  eja & EJB & eje  |  eja & ejb & EJE  |  eja & ejb & eje  ; 
assign JQA = ~jqa;  //complement 
assign ccf = ~CCF;  //complement 
assign ccn = ~CCN;  //complement 
assign cgf = ~CGF;  //complement 
assign cgn = ~CGN;  //complement 
assign AAF = ~aaf;  //complement 
assign ABF = ~abf;  //complement 
assign ACF = ~acf;  //complement 
assign ADF = ~adf;  //complement 
assign AAN = ~aan;  //complement 
assign ABN = ~abn;  //complement 
assign ACN = ~acn;  //complement 
assign ADN = ~adn;  //complement 
assign chf = ~CHF;  //complement 
assign chn = ~CHN;  //complement 
assign oen = ~OEN;  //complement 
assign dif = ~DIF;  //complement 
assign cif = ~CIF;  //complement 
assign AAV = ~aav;  //complement 
assign ABV = ~abv;  //complement 
assign ACV = ~acv;  //complement 
assign ADV = ~adv;  //complement 
assign JID =  psf & pse & PSD  ; 
assign jid = ~JID;  //complement 
assign JIE =  psf & PSE & psd  ; 
assign jie = ~JIE;  //complement 
assign naf = ~NAF;  //complement 
assign paf = ~PAF;  //complement 
assign hbf = ~HBF;  //complement 
assign oif = ~OIF;  //complement 
assign onc = ~ONC;  //complement 
assign ooc = ~OOC;  //complement 
assign KFB =  DNB & dje & dme  |  dnb & DJE & dme  |  dnb & dje & DME  |  DNB & DJE & DME  ; 
assign kfb = ~KFB; //complement 
assign KFC =  DKE & dif  |  dke & DIF  ; 
assign kfc = ~KFC; //complement 
assign KFD =  DKE & dif  |  dke & DIF  ; 
assign kfd = ~KFD;  //complement 
assign oaf = ~OAF;  //complement 
assign oef = ~OEF;  //complement 
assign ocf = ~OCF;  //complement 
assign ogf = ~OGF;  //complement 
assign eif = ~EIF;  //complement 
assign haf = ~HAF;  //complement 
assign FAC =  EEH & EIG & eif & EIE & jja  ; 
assign fac = ~FAC;  //complement  
assign fcf =  eif  ; 
assign FCF = ~fcf;  //complement 
assign oan = ~OAN;  //complement 
assign ocn = ~OCN;  //complement 
assign ogn = ~OGN;  //complement 
assign ejf = ~EJF;  //complement 
assign FBC =  EJH & EJG & ejf & EJE & jjb  ; 
assign fbc = ~FBC;  //complement  
assign obf = ~OBF;  //complement 
assign off = ~OFF;  //complement 
assign odf = ~ODF;  //complement 
assign ohf = ~OHF;  //complement 
assign ekf = ~EKF;  //complement 
assign GAF =  ekd & EKC & ekb & EKA  ; 
assign gaf = ~GAF;  //complement  
assign GBF =  ekh & EKG & ekf & EKE  ; 
assign gbf = ~GBF;  //complement 
assign obn = ~OBN;  //complement 
assign ofn = ~OFN;  //complement 
assign odn = ~ODN;  //complement 
assign ohn = ~OHN;  //complement 
assign bag = ~BAG;  //complement 
assign bbg = ~BBG;  //complement 
assign bcg = ~BCG;  //complement 
assign bdg = ~BDG;  //complement 
assign bao = ~BAO;  //complement 
assign bbo = ~BBO;  //complement 
assign bco = ~BCO;  //complement 
assign bdo = ~BDO;  //complement 
assign baw = ~BAW;  //complement 
assign bbw = ~BBW;  //complement 
assign bcw = ~BCW;  //complement 
assign bdw = ~BDW;  //complement 
assign dag = ~DAG;  //complement 
assign dbg = ~DBG;  //complement 
assign eag = ~EAG;  //complement 
assign ebg = ~EBG;  //complement 
assign dcg = ~DCG;  //complement 
assign ddg = ~DDG;  //complement 
assign ecg = ~ECG;  //complement 
assign edg = ~EDG;  //complement 
assign deg = ~DEG;  //complement 
assign dfg = ~DFG;  //complement 
assign eeg = ~EEG;  //complement 
assign efg = ~EFG;  //complement 
assign dgg = ~DGG;  //complement 
assign dhg = ~DHG;  //complement 
assign egg = ~EGG;  //complement 
assign ehg = ~EHG;  //complement 
assign cdg = ~CDG;  //complement 
assign cdo = ~CDO;  //complement 
assign ABC = ~abc;  //complement 
assign ceg = ~CEG;  //complement 
assign ceo = ~CEO;  //complement 
assign cfg = ~CFG;  //complement 
assign cfo = ~CFO;  //complement 
assign cbg = ~CBG;  //complement 
assign laa = ~LAA;  //complement 
assign LBA = ~lba;  //complement 
assign KGA =  DOC & dpc & dqc  |  doc & DPC & dqc  |  doc & dpc & DQC  |  DOC & DPC & DQC  ; 
assign kga = ~KGA; //complement 
assign cag = ~CAG;  //complement 
assign cao = ~CAO;  //complement 
assign cbo = ~CBO;  //complement 
assign opa = ~OPA;  //complement 
assign ccg = ~CCG;  //complement 
assign cco = ~CCO;  //complement 
assign cgg = ~CGG;  //complement 
assign cgo = ~CGO;  //complement 
assign AAG = ~aag;  //complement 
assign ABG = ~abg;  //complement 
assign ACG = ~acg;  //complement 
assign ADG = ~adg;  //complement 
assign mac =  lba & lbb & lbc  ; 
assign MAC = ~mac;  //complement 
assign chg = ~CHG;  //complement 
assign cho = ~CHO;  //complement 
assign AAO = ~aao;  //complement 
assign ABO = ~abo;  //complement 
assign ACO = ~aco;  //complement 
assign ADO = ~ado;  //complement 
assign MAA =  LAA & lab & lac  |  laa & LAB & lac  |  laa & lab & LAC  |  LAA & LAB & LAC  ; 
assign maa = ~MAA; //complement 
assign mab =  LAA & lab & lac  |  laa & LAB & lac  |  laa & lab & LAC  |  laa & lab & lac  ; 
assign MAB = ~mab;  //complement 
assign cig = ~CIG;  //complement 
assign AAW = ~aaw;  //complement 
assign ABW = ~abw;  //complement 
assign ACW = ~acw;  //complement 
assign ADW = ~adw;  //complement 
assign lab = ~LAB;  //complement 
assign LBB = ~lbb;  //complement 
assign lac = ~LAC;  //complement 
assign LBC = ~lbc;  //complement 
assign oja = ~OJA;  //complement 
assign OJB = ~ojb;  //complement 
assign hbg = ~HBG;  //complement 
assign oig = ~OIG;  //complement 
assign ona = ~ONA;  //complement 
assign ooa = ~OOA;  //complement 
assign KGB =  DNC & dle & dme  |  dnc & DLE & dme  |  dnc & dle & DME  |  DNC & DLE & DME  ; 
assign kgb = ~KGB; //complement 
assign KGC =  DJE & dig  |  dje & DIG  ; 
assign kgc = ~KGC; //complement 
assign KGD =  DJE & dig  |  dje & DIG  ; 
assign kgd = ~KGD;  //complement 
assign oag = ~OAG;  //complement 
assign oeg = ~OEG;  //complement 
assign ocg = ~OCG;  //complement 
assign ogg = ~OGG;  //complement 
assign eig = ~EIG;  //complement 
assign hag = ~HAG;  //complement 
assign FAB =  EIH & eig & EIF & EIE & jja  ; 
assign fab = ~FAB;  //complement  
assign fcg =  eig  ; 
assign FCG = ~fcg;  //complement 
assign oao = ~OAO;  //complement 
assign oeo = ~OEO;  //complement 
assign oco = ~OCO;  //complement 
assign ogo = ~OGO;  //complement 
assign ejg = ~EJG;  //complement 
assign dig = ~DIG;  //complement 
assign FBB =  EJH & ejg & EJF & EJE & jib  ; 
assign fbb = ~FBB;  //complement  
assign obg = ~OBG;  //complement 
assign ofg = ~OFG;  //complement 
assign odg = ~ODG;  //complement 
assign ohg = ~OHG;  //complement 
assign ekg = ~EKG;  //complement 
assign GAG =  ekd & EKC & EKB & eka  ; 
assign gag = ~GAG;  //complement  
assign GBG =  ekh & EKG & EKF & eke  ; 
assign gbg = ~GBG;  //complement 
assign obo = ~OBO;  //complement 
assign ofo = ~OFO;  //complement 
assign odo = ~ODO;  //complement 
assign oho = ~OHO;  //complement 
assign bah = ~BAH;  //complement 
assign bbh = ~BBH;  //complement 
assign bch = ~BCH;  //complement 
assign bdh = ~BDH;  //complement 
assign bap = ~BAP;  //complement 
assign bbp = ~BBP;  //complement 
assign bcp = ~BCP;  //complement 
assign bdp = ~BDP;  //complement 
assign bax = ~BAX;  //complement 
assign bbx = ~BBX;  //complement 
assign bcx = ~BCX;  //complement 
assign bdx = ~BDX;  //complement 
assign dah = ~DAH;  //complement 
assign dbh = ~DBH;  //complement 
assign eah = ~EAH;  //complement 
assign ebh = ~EBH;  //complement 
assign dch = ~DCH;  //complement 
assign ddh = ~DDH;  //complement 
assign ech = ~ECH;  //complement 
assign edh = ~EDH;  //complement 
assign deh = ~DEH;  //complement 
assign dfh = ~DFH;  //complement 
assign eeh = ~EEH;  //complement 
assign efh = ~EFH;  //complement 
assign dgh = ~DGH;  //complement 
assign dhh = ~DHH;  //complement 
assign egh = ~EGH;  //complement 
assign ehh = ~EHH;  //complement 
assign cdp = ~CDP;  //complement 
assign JDF =  CDH  ; 
assign jdf = ~JDF;  //complement 
assign ceh = ~CEH;  //complement 
assign cep = ~CEP;  //complement 
assign JEF =  CEH  ; 
assign jef = ~JEF;  //complement 
assign cfh = ~CFH;  //complement 
assign cbh = ~CBH;  //complement 
assign tad = ~TAD;  //complement 
assign tbd = ~TBD;  //complement 
assign tcd = ~TCD;  //complement 
assign tdd = ~TDD;  //complement 
assign tae = ~TAE;  //complement 
assign tbe = ~TBE;  //complement 
assign tce = ~TCE;  //complement 
assign tde = ~TDE;  //complement 
assign taf = ~TAF;  //complement 
assign tbf = ~TBF;  //complement 
assign tcf = ~TCF;  //complement 
assign tdf = ~TDF;  //complement 
assign tai = ~TAI;  //complement 
assign tbi = ~TBI;  //complement 
assign tci = ~TCI;  //complement 
assign tdi = ~TDI;  //complement 
assign tac = ~TAC;  //complement 
assign tcc = ~TCC;  //complement 
assign tdc = ~TDC;  //complement 
assign tab = ~TAB;  //complement 
assign tbb = ~TBB;  //complement 
assign tcb = ~TCB;  //complement 
assign tdb = ~TDB;  //complement 
assign taa = ~TAA;  //complement 
assign tba = ~TBA;  //complement 
assign tca = ~TCA;  //complement 
assign tda = ~TDA;  //complement 
assign KHA =  DOD & dpd & dqd  |  dod & DPD & dqd  |  dod & dpd & DQD  |  DOD & DPD & DQD  ; 
assign kha = ~KHA; //complement 
assign cah = ~CAH;  //complement 
assign cap = ~CAP;  //complement 
assign JAF =  CAH  ; 
assign jaf = ~JAF;  //complement 
assign JFF =  CFH  ; 
assign jff = ~JFF;  //complement 
assign cbp = ~CBP;  //complement 
assign jqb =  EJF & ejg & ejh  |  ejf & EJG & ejh  |  ejf & ejg & EJH  |  ejf & ejg & ejh  ; 
assign JQB = ~jqb;  //complement 
assign JBF =  CBH  ; 
assign jbf = ~JBF;  //complement 
assign JQC =  EKC & EKD  |  EKC  ; 
assign jqc = ~JQC; //complement 
assign cch = ~CCH;  //complement 
assign ccp = ~CCP;  //complement 
assign JCF =  CCH  ; 
assign jcf = ~JCF;  //complement 
assign KHB =  DND & dle & dme  |  dnd & DLE & dme  |  dnd & dle & DME  |  DND & DLE & DME  ; 
assign khb = ~KHB; //complement 
assign JGF =  CGH  ; 
assign jgf = ~JGF;  //complement 
assign cgh = ~CGH;  //complement 
assign cgp = ~CGP;  //complement 
assign AAH = ~aah;  //complement 
assign ABH = ~abh;  //complement 
assign ACH = ~ach;  //complement 
assign ADH = ~adh;  //complement 
assign JJA = ~jja;  //complement 
assign JJB = ~jjb;  //complement 
assign JHF =  CHH  ; 
assign jhf = ~JHF;  //complement 
assign chh = ~CHH;  //complement 
assign chp = ~CHP;  //complement 
assign AAP = ~aap;  //complement 
assign ABP = ~abp;  //complement 
assign ACP = ~acp;  //complement 
assign ADP = ~adp;  //complement 
assign JPA =  PCA & pcb & pcc  |  pca & PCB & pcc  |  pca & pcb & PCC  |  PCA & PCB & PCC  ; 
assign jpa = ~JPA; //complement 
assign pca = ~PCA;  //complement 
assign cih = ~CIH;  //complement 
assign AAX = ~aax;  //complement 
assign ABX = ~abx;  //complement 
assign ACX = ~acx;  //complement 
assign ADX = ~adx;  //complement 
assign tah = ~TAH;  //complement 
assign tbh = ~TBH;  //complement 
assign tch = ~TCH;  //complement 
assign tdh = ~TDH;  //complement 
assign tag = ~TAG;  //complement 
assign tbg = ~TBG;  //complement 
assign tcg = ~TCG;  //complement 
assign tdg = ~TDG;  //complement 
assign qaa = ~QAA;  //complement 
assign qab = ~QAB;  //complement 
assign qac = ~QAC;  //complement 
assign qad = ~QAD;  //complement 
assign hbh = ~HBH;  //complement 
assign oih = ~OIH;  //complement 
assign onb = ~ONB;  //complement 
assign oob = ~OOB;  //complement 
assign ohh = ~OHH;  //complement 
assign KHC =  DKE & dih  |  dke & DIH  ; 
assign khc = ~KHC; //complement 
assign KHD =  DKE & dih  |  dke & DIH  ; 
assign khd = ~KHD;  //complement 
assign oah = ~OAH;  //complement 
assign oeh = ~OEH;  //complement 
assign och = ~OCH;  //complement 
assign ogh = ~OGH;  //complement 
assign eih = ~EIH;  //complement 
assign hah = ~HAH;  //complement 
assign FAA =  eih & EIG & EIF & EIE & jja  ; 
assign faa = ~FAA;  //complement  
assign fch =  eih  ; 
assign FCH = ~fch;  //complement 
assign oap = ~OAP;  //complement 
assign oep = ~OEP;  //complement 
assign ocp = ~OCP;  //complement 
assign ogp = ~OGP;  //complement 
assign ejh = ~EJH;  //complement 
assign dih = ~DIH;  //complement 
assign FBA =  ejh & EJG & EJF & EJE & jjb  ; 
assign fba = ~FBA;  //complement  
assign obh = ~OBH;  //complement 
assign ofh = ~OFH;  //complement 
assign odh = ~ODH;  //complement 
assign ekh = ~EKH;  //complement 
assign GAH =  EKD & EKC & EKB & EKA  ; 
assign gah = ~GAH;  //complement  
assign GBH =  EKH & EKG & EKF & EKE  ; 
assign gbh = ~GBH;  //complement 
assign obp = ~OBP;  //complement 
assign ofp = ~OFP;  //complement 
assign odp = ~ODP;  //complement 
assign ohp = ~OHP;  //complement 
assign iaa = ~IAA; //complement 
assign iab = ~IAB; //complement 
assign iac = ~IAC; //complement 
assign iad = ~IAD; //complement 
assign iae = ~IAE; //complement 
assign iaf = ~IAF; //complement 
assign iag = ~IAG; //complement 
assign iah = ~IAH; //complement 
assign iai = ~IAI; //complement 
assign iaj = ~IAJ; //complement 
assign iak = ~IAK; //complement 
assign ial = ~IAL; //complement 
assign iam = ~IAM; //complement 
assign ian = ~IAN; //complement 
assign iao = ~IAO; //complement 
assign iap = ~IAP; //complement 
assign iaq = ~IAQ; //complement 
assign iar = ~IAR; //complement 
assign ias = ~IAS; //complement 
assign iat = ~IAT; //complement 
assign iau = ~IAU; //complement 
assign iav = ~IAV; //complement 
assign iaw = ~IAW; //complement 
assign iax = ~IAX; //complement 
assign iba = ~IBA; //complement 
assign ibb = ~IBB; //complement 
assign ibc = ~IBC; //complement 
assign ibd = ~IBD; //complement 
assign ibe = ~IBE; //complement 
assign ibf = ~IBF; //complement 
assign ibg = ~IBG; //complement 
assign ibh = ~IBH; //complement 
assign ibi = ~IBI; //complement 
assign ibj = ~IBJ; //complement 
assign ibk = ~IBK; //complement 
assign ibl = ~IBL; //complement 
assign ibm = ~IBM; //complement 
assign ibn = ~IBN; //complement 
assign ibo = ~IBO; //complement 
assign ibp = ~IBP; //complement 
assign ibq = ~IBQ; //complement 
assign ibr = ~IBR; //complement 
assign ibs = ~IBS; //complement 
assign ibt = ~IBT; //complement 
assign ibu = ~IBU; //complement 
assign ibv = ~IBV; //complement 
assign ibw = ~IBW; //complement 
assign ibx = ~IBX; //complement 
assign ica = ~ICA; //complement 
assign icb = ~ICB; //complement 
assign icc = ~ICC; //complement 
assign icd = ~ICD; //complement 
assign ice = ~ICE; //complement 
assign icf = ~ICF; //complement 
assign icg = ~ICG; //complement 
assign ich = ~ICH; //complement 
assign ici = ~ICI; //complement 
assign icj = ~ICJ; //complement 
assign ick = ~ICK; //complement 
assign icl = ~ICL; //complement 
assign icm = ~ICM; //complement 
assign icn = ~ICN; //complement 
assign ico = ~ICO; //complement 
assign icp = ~ICP; //complement 
assign icq = ~ICQ; //complement 
assign icr = ~ICR; //complement 
assign ics = ~ICS; //complement 
assign ict = ~ICT; //complement 
assign icu = ~ICU; //complement 
assign icv = ~ICV; //complement 
assign icw = ~ICW; //complement 
assign icx = ~ICX; //complement 
assign ida = ~IDA; //complement 
assign idb = ~IDB; //complement 
assign idc = ~IDC; //complement 
assign idd = ~IDD; //complement 
assign ide = ~IDE; //complement 
assign idf = ~IDF; //complement 
assign idg = ~IDG; //complement 
assign idh = ~IDH; //complement 
assign idi = ~IDI; //complement 
assign idj = ~IDJ; //complement 
assign idk = ~IDK; //complement 
assign idl = ~IDL; //complement 
assign idm = ~IDM; //complement 
assign idn = ~IDN; //complement 
assign ido = ~IDO; //complement 
assign idp = ~IDP; //complement 
assign idq = ~IDQ; //complement 
assign idr = ~IDR; //complement 
assign ids = ~IDS; //complement 
assign idt = ~IDT; //complement 
assign idu = ~IDU; //complement 
assign idv = ~IDV; //complement 
assign idw = ~IDW; //complement 
assign idx = ~IDX; //complement 
assign iea = ~IEA; //complement 
assign ieb = ~IEB; //complement 
assign iec = ~IEC; //complement 
assign ied = ~IED; //complement 
assign iee = ~IEE; //complement 
assign ief = ~IEF; //complement 
assign ifa = ~IFA; //complement 
assign ifb = ~IFB; //complement 
assign ifc = ~IFC; //complement 
assign ifd = ~IFD; //complement 
assign ife = ~IFE; //complement 
assign ifff  = ~IFFF ; //complement 
assign iga = ~IGA; //complement 
assign igb = ~IGB; //complement 
assign igc = ~IGC; //complement 
assign igd = ~IGD; //complement 
assign ige = ~IGE; //complement 
assign igf = ~IGF; //complement 
assign iha = ~IHA; //complement 
assign ihb = ~IHB; //complement 
assign ihc = ~IHC; //complement 
assign ihd = ~IHD; //complement 
assign ihe = ~IHE; //complement 
assign ihf = ~IHF; //complement 
assign iia = ~IIA; //complement 
assign ija = ~IJA; //complement 
always@(posedge IZZ )
   begin 
 BAA <= AAA ; 
 BBA <= ABA ; 
 BCA <= ACA ; 
 BDA <= ADA ; 
 BAI <= AAI ; 
 BBI <= ABI ; 
 BCI <= ACI ; 
 BDI <= ADI ; 
 EGA <= DGA ; 
 BAQ <= AAQ ; 
 BBQ <= ABQ ; 
 BCQ <= ACQ ; 
 BDQ <= ADQ ; 
 NBA <= NAA ; 
 NCA <= NBA ; 
 NEA <= NDA ; 
 NDA <= NCA ; 
 NFA <= NEA ; 
 NGA <= NFA ; 
 NHA <= NGA ; 
 NIA <= NHA ; 
 NJA <= NIA ; 
 NKA <= NJA ; 
 NLA <= NKA ; 
 NMA <= NLA ; 
 NNA <= NMA ; 
 NOA <= NNA ; 
 NPA <= NOA ; 
 NQA <= NPA ; 
 DAA <= CAI ; 
 DBA <= CBI ; 
 EAA <= DAA ; 
 EBA <= DBA ; 
 DCA <= CCI ; 
 DDA <= CDI ; 
 ECA <= DCA ; 
 EDA <= DDA ; 
 DEA <= CEI ; 
 DFA <= CFI ; 
 EEA <= DEA ; 
 EFA <= DFA ; 
 DGA <= CGI ; 
 DHA <= CHI ; 
 EHA <= DHA ; 
 CDA <=  AAA & TAD  |  ABA & TBD  |  ACA & TCD  |  ADA & TDD  ; 
 CDI <=  AAA & TAD  |  ABA & TBD  |  ACA & TCD  |  ADA & TDD  ; 
 DMA <=  JDD & jdf  |  jdd & JDF  |  jdd & jdf  |  JDD & JDF  ;
 CEA <=  AAI & TAE  |  ABI & TBE  |  ACI & TCE  |  ADI & TDE  ; 
 CEI <=  AAI & TAE  |  ABI & TBE  |  ACI & TCE  |  ADI & TDE  ; 
 DNA <=  JED & jef  |  jed & JEF  |  jed & jef  |  JED & JEF  ;
 CFA <=  AAQ & TAF  |  ABQ & TBF  |  ACQ & TCF  |  ADQ & TDF  ; 
 CFI <=  AAQ & TAF  |  ABQ & TBF  |  ACQ & TCF  |  ADQ & TDF  ; 
 DOA <=  JFD & jff  |  jfd & JFF  |  jfd & jff  |  JFD & JFF  ;
 NRA <= NQA ; 
 NSA <= NRA ; 
 CAA <=  BAA & TAA  |  BBA & TBA  |  BCA & TCA  |  BDA & TDA  ; 
 CAI <=  BAA & TAA  |  BBA & TBA  |  BCA & TCA  |  BDA & TDA  ; 
 DJA <=  JAD & jaf  |  jad & JAF  |  jad & jaf  |  JAD & JAF  ;
 CBA <=  BAI & TAB  |  BBI & TBB  |  BCI & TCB  |  BDI & TDB  ; 
 CBI <=  BAI & TAB  |  BBI & TBB  |  BCI & TCB  |  BDI & TDB  ; 
 DKA <=  JBD & jbf  |  jbd & JBF  |  jbd & jbf  |  JBD & JBF  ;
 CCA <=  BAQ & TAC  |  BBQ & TBC  |  BCQ & TCC  |  BDQ & TDC  ; 
 CCI <=  BAQ & TAC  |  BBQ & TBC  |  BCQ & TCC  |  BDQ & TDC  ; 
 DLA <=  JCD & jcf  |  jcd & JCF  |  jcd & jcf  |  JCD & JCF  ;
 OAI <=  FAB & GAA & eba  |  fab & EBA  |  gaa & EBA  ; 
 CGA <=  IAA & TAG  |  IBA & TBG  |  ICA & TCG  |  IDA & TDG  ; 
 CGI <=  IAA & TAG  |  IBA & TBG  |  ICA & TCG  |  IDA & TDG  ; 
 aaa <= iaa ; 
 aba <= iba ; 
 aca <= ica ; 
 ada <= ida ; 
 CHA <=  IAI & TAH  |  IBI & TBH  |  ICI & TCH  |  IDI & TDH  ; 
 CHI <=  IAI & TAH  |  IBI & TBH  |  ICI & TCH  |  IDI & TDH  ; 
 aai <= iai ; 
 abi <= ibi ; 
 aci <= ici ; 
 adi <= idi ; 
 DPA <=  JGD & jgf  |  jgd & JGF  |  jgd & jgf  |  JGD & JGF  ;
 DQA <=  JHD & jhf  |  jhd & JHF  |  jhd & jhf  |  JHD & JHF  ;
 CIA <=  IAQ & TAI  |  IBQ & TBI  |  ICQ & TCI  |  IDQ & TDI  ; 
 aaq <= iaq ; 
 abq <= ibq ; 
 acq <= icq ; 
 adq <= idq ; 
 PCB <=  DNE & dqe & dpe  |  dne & DQE & dpe  |  dne & dqe & DPE  |  DNE & DQE & DPE  ;
 OMA <= NAA ; 
 NAA <=  IEA  |  IFA  |  IGA  |  IHA  ; 
 HBA <= HAA ; 
 OIA <= HBA ; 
 OKA <= NSA ; 
 OLA <= NSA ; 
 OAA <=  FAA & GAA & eaa  |  faa & EAA  |  gaa & EAA  ; 
 OEA <=  FAA & GAA & eaa  |  faa & EAA  |  gaa & EAA  ; 
 OCA <=  FAE & GBA & eea  |  fae & EEA  |  gba & EEA  ; 
 OGA <=  FAE & GBA & eea  |  fae & EEA  |  gba & EEA  ; 
 EIA <=  KAA & kab & kac  |  kaa & KAB & kac  |  kaa & kab & KAC  |  KAA & KAB & KAC  ;
 OEI <=  FAB & GAA & eba  |  fab & EBA  |  gaa & EBA  ; 
 OCI <=  FAF & GBA & efa  |  faf & EFA  |  gba & EFA  ; 
 OGI <=  FAF & GBA & efa  |  faf & EFA  |  gba & EFA  ; 
 EJA <=  KAA & kab & kac  |  kaa & KAB & kac  |  kaa & kab & KAC  |  KAA & KAB & KAC  ;
 DIA <= CIA ; 
 OBA <=  FAC & GAA & eca  |  fac & ECA  |  gaa & ECA  ; 
 OFA <=  FAC & GAA & eca  |  fac & ECA  |  gaa & ECA  ; 
 ODA <=  FAG & GBA & ega  |  fag & EGA  |  gba & EGA  ; 
 OHA <=  FAG & GBA & ega  |  fag & EGA  |  gba & EGA  ; 
 EKA <=  KAA & kab & kad  |  kaa & KAB & kad  |  kaa & kab & KAD  |  KAA & KAB & KAD  ;
 OBI <=  FAD & GAA & eda  |  fad & EDA  |  gaa & EDA  ; 
 OFI <=  FAD & GAA & eda  |  fad & EDA  |  gaa & EDA  ; 
 ODI <=  FAH & GBA & eha  |  fah & EHA  |  gba & EHA  ; 
 OHI <=  FAH & GBA & eha  |  fah & EHA  |  gba & EHA  ; 
 BAB <= AAB ; 
 BBB <= ABB ; 
 BCB <= ACB ; 
 BDB <= ADB ; 
 BAJ <= AAJ ; 
 BBJ <= ABJ ; 
 BCJ <= ACJ ; 
 BDJ <= ADJ ; 
 BAR <= AAR ; 
 BBR <= ABR ; 
 BCR <= ACR ; 
 BDR <= ADR ; 
 ECB <= DCB ; 
 EDB <= DDB ; 
 NBB <= NAB ; 
 NCB <= NBB ; 
 NFB <= NEB ; 
 NGB <= NFB ; 
 NHB <= NGB ; 
 NIB <= NHB ; 
 NJB <= NIB ; 
 NKB <= NJB ; 
 NLB <= NKB ; 
 NMB <= NLB ; 
 NNB <= NMB ; 
 NOB <= NNB ; 
 NPB <= NOB ; 
 NQB <= NPB ; 
 DAB <= CAJ ; 
 DBB <= CBJ ; 
 EAB <= DAB ; 
 EBB <= DBB ; 
 DCB <= CCJ ; 
 DDB <= CDJ ; 
 DEB <= CEJ ; 
 DFB <= CFJ ; 
 EEB <= DEB ; 
 EFB <= DFB ; 
 NDB <= NCB ; 
 NEB <= NDB ; 
 HAA <= FCA ; 
 HAB <= FCB ; 
 DGB <= CGJ ; 
 DHB <= CHJ ; 
 EGB <= DGB ; 
 EHB <= DHB ; 
 CDB <=  AAB & TAD  |  ABB & TBD  |  ACB & TCD  |  ADB & TDD  ; 
 CDJ <=  AAB & TAD  |  ABB & TBD  |  ACB & TCD  |  ADB & TDD  ; 
 DMB <=  JDE & jdf  |  jde & JDF  |  jde & jdf  |  JDE & JDF  ;
 CEB <=  AAJ & TAE  |  ABJ & TBE  |  ACJ & TCE  |  ADJ & TDE  ; 
 CEJ <=  AAJ & TAE  |  ABJ & TBE  |  ACJ & TCE  |  ADJ & TDE  ; 
 ack <= ick ; 
 CFB <=  AAR & TAF  |  ABR & TBF  |  ACR & TCF  |  ADR & TDF  ; 
 CFJ <=  AAR & TAF  |  ABR & TBF  |  ACR & TCF  |  ADR & TDF  ; 
 DOB <=  JFE & jff  |  jfe & JFF  |  jfe & jff  |  JFE & JFF  ;
 NRB <= NQB ; 
 NSB <= NRB ; 
 DNB <=  JEE & jef  |  jee & JEF  |  jee & jef  |  JEE & JEF  ;
 DKB <=  JBE & jbf  |  jbe & JBF  |  jbe & jbf  |  JBE & JBF  ;
 CAB <=  BAB & TAA  |  BBB & TBA  |  BCB & TCA  |  BDB & TDA  ; 
 CAJ <=  BAB & TAA  |  BBB & TBA  |  BCB & TCA  |  BDB & TDA  ; 
 DJB <=  JAE & jaf  |  jae & JAF  |  jae & jaf  |  JAE & JAF  ;
 CBB <=  BAJ & TAB  |  BBJ & TBB  |  BCJ & TCB  |  BDJ & TDB  ; 
 CBJ <=  BAJ & TAB  |  BBJ & TBB  |  BCJ & TCB  |  BDJ & TDB  ; 
 CCB <=  BAR & TAC  |  BBR & TBC  |  BCR & TCC  |  BDR & TDC  ; 
 CCJ <=  BAR & TAC  |  BBR & TBC  |  BCR & TCC  |  BDR & TDC  ; 
 DLB <=  JCE & jcf  |  jce & JCF  |  jce & jcf  |  JCE & JCF  ;
 DQB <=  JHE & jhf  |  jhe & JHF  |  jhe & jhf  |  JHE & JHF  ;
 CGB <=  IAB & TAG  |  IBB & TBG  |  ICB & TCG  |  IDB & TDG  ; 
 CGJ <=  IAB & TAG  |  IBB & TBG  |  ICB & TCG  |  IDB & TDG  ; 
 aab <= iab ; 
 abb <= ibb ; 
 acb <= icb ; 
 adb <= idb ; 
 CHB <=  IAJ & TAH  |  IBJ & TBH  |  ICJ & TCH  |  IDJ & TDH  ; 
 CHJ <=  IAJ & TAH  |  IBJ & TBH  |  ICJ & TCH  |  IDJ & TDH  ; 
 aaj <= iaj ; 
 abj <= ibj ; 
 acj <= icj ; 
 adj <= idj ; 
 DPB <=  JGE & jgf  |  jge & JGF  |  jge & jgf  |  JGE & JGF  ;
 OFJ <=  FAD & GAB & edb  |  fad & EDB  |  gab & EDB  ; 
 CIB <=  IAR & TAI  |  IBR & TBI  |  ICR & TCI  |  IDR & TDI  ; 
 aar <= iar ; 
 abr <= ibr ; 
 acr <= icr ; 
 adr <= idr ; 
 OMB <= NAB ; 
 NAB <=  IEB  |  IFB  |  IGB  |  IHB  ; 
 HBB <= HAB ; 
 OIB <= HBB ; 
 OKB <= NSB ; 
 OLB <= NSB ; 
 OHB <=  FAG & GBB & egb  |  fag & EGB  |  gbb & EGB  ; 
 OAB <=  FAA & GAB & eab  |  faa & EAB  |  gab & EAB  ; 
 OEB <=  FAA & GAB & eab  |  faa & EAB  |  gab & EAB  ; 
 OCB <=  FAE & GBB & eeb  |  fae & EEB  |  gbb & EEB  ; 
 OGB <=  FAE & GBB & eeb  |  fae & EEB  |  gbb & EEB  ; 
 EIB <=  KBA & kbb & kbc  |  kba & KBB & kbc  |  kba & kbb & KBC  |  KBA & KBB & KBC  ;
 OAJ <=  FAB & GAB & ebb  |  fab & EBB  |  gab & EBB  ; 
 OEJ <=  FAB & GAB & ebb  |  fab & EBB  |  gab & EBB  ; 
 OCJ <=  FAF & GBB & efb  |  faf & EFB  |  gbb & EFB  ; 
 OGJ <=  FAF & GBB & efb  |  faf & EFB  |  gbb & EFB  ; 
 EJB <=  KBA & kbb & kbc  |  kba & KBB & kbc  |  kba & kbb & KBC  |  KBA & KBB & KBC  ;
 DIB <= CIB ; 
 OBB <=  FAC & GAB & ecb  |  fac & ECB  |  gab & ECB  ; 
 OFB <=  FAC & GAB & ecb  |  fac & ECB  |  gab & ECB  ; 
 ODB <=  FAG & GBB & egb  |  fag & EGB  |  gbb & EGB  ; 
 EKB <=  KBA & kbb & kbd  |  kba & KBB & kbd  |  kba & kbb & KBD  |  KBA & KBB & KBD  ;
 OBJ <=  FAD & GAB & edb  |  fad & EDB  |  gab & EDB  ; 
 ODJ <=  FAH & GBB & ehb  |  fah & EHB  |  gbb & EHB  ; 
 OHJ <=  FAH & GBB & ehb  |  fah & EHB  |  gbb & EHB  ; 
 BAC <= AAC ; 
 BBC <= ABC ; 
 BCC <= ACC ; 
 BDC <= ADC ; 
 BAK <= AAK ; 
 BBK <= ABK ; 
 BCK <= ACK ; 
 BDK <= ADK ; 
 BDS <= ADS ; 
 BAS <= AAS ; 
 BAT <= AAT ; 
 BBS <= ABS ; 
 BCS <= ACS ; 
 NBC <= NAC ; 
 NCC <= NBC ; 
 NEC <= NDC ; 
 NDC <= NCC ; 
 NFC <= NEC ; 
 NGC <= NFC ; 
 NHC <= NGC ; 
 NIC <= NHC ; 
 NJC <= NIC ; 
 NKC <= NJC ; 
 NLC <= NKC ; 
 NMC <= NLC ; 
 NNC <= NMC ; 
 NOC <= NNC ; 
 NPC <= NOC ; 
 NQC <= NPC ; 
 DAC <= CAK ; 
 DBC <= CBK ; 
 DBD <= CBL ; 
 EAC <= DAC ; 
 EAD <= DAD ; 
 EBC <= DBC ; 
 EBD <= DBD ; 
 DCD <= CCL ; 
 DDC <= CDK ; 
 ECC <= DCC ; 
 EDC <= DDC ; 
 EFC <= DFC ; 
 EFD <= DFD ; 
 DEC <= CEK ; 
 DFC <= CFK ; 
 DFD <= CFL ; 
 EEC <= DEC ; 
 EHD <= DHD ; 
 DCC <= CCK ; 
 DGC <= CGK ; 
 DHC <= CHK ; 
 EGC <= DGC ; 
 EHC <= DHC ; 
 CDC <=  AAC & TAD  |  ABC & TBD  |  ACC & TCD  |  ADC & TDD  ; 
 CDK <=  AAC & TAD  |  ABC & TBD  |  ACC & TCD  |  ADC & TDD  ; 
 DKC <=  JBA & jbg  |  jba & JBG  |  jba & jbg  |  JBA & JBG  ;
 DMC <=  JDA & jdg  |  jda & JDG  |  jda & jdg  |  JDA & JDG  ;
 CEC <=  AAK & TAE  |  ABK & TBE  |  ACK & TCE  |  ADK & TDE  ; 
 CEK <=  AAK & TAE  |  ABK & TBE  |  ACK & TCE  |  ADK & TDE  ; 
 DNC <=  JEA & jeg  |  jea & JEG  |  jea & jeg  |  JEA & JEG  ;
 CFC <=  AAS & TAF  |  ABS & TBF  |  ACS & TCF  |  ADS & TDF  ; 
 CFK <=  AAS & TAF  |  ABS & TBF  |  ACS & TCF  |  ADS & TDF  ; 
 CFP <=  AAX & TAF  |  ABX & TBF  |  ACX & TCF  |  ADX & TDF  ; 
 DOC <=  JFA & jfg  |  jfa & JFG  |  jfa & jfg  |  JFA & JFG  ;
 NRC <= NQC ; 
 NSC <= NRC ; 
 TBC <= QAA ; 
 CAC <=  BAC & TAA  |  BBC & TBA  |  BCC & TCA  |  BDC & TDA  ; 
 CAK <=  BAC & TAA  |  BBC & TBA  |  BCC & TCA  |  BDC & TDA  ; 
 DJC <=  JAA & jag  |  jaa & JAG  |  jaa & jag  |  JAA & JAG  ;
 CBC <=  BAK & TAB  |  BBK & TBB  |  BCK & TCB  |  BDK & TDB  ; 
 CBK <=  BAK & TAB  |  BBK & TBB  |  BCK & TCB  |  BDK & TDB  ; 
 CCC <=  BAS & TAC  |  BBS & TBC  |  BCS & TCC  |  BDS & TDC  ; 
 CCK <=  BAS & TAC  |  BBS & TBC  |  BCS & TCC  |  BDS & TDC  ; 
 DLC <=  JCA & jcg  |  jca & JCG  |  jca & jcg  |  JCA & JCG  ;
 OFK <=  FAD & GAC & edc  |  fad & EDC  |  gac & EDC  ; 
 CGC <=  IAC & TAG  |  IBC & TBG  |  ICC & TCG  |  IDC & TDG  ; 
 CGK <=  IAC & TAG  |  IBC & TBG  |  ICC & TCG  |  IDC & TDG  ; 
 aac <= iac ; 
 acc <= icc ; 
 adc <= idc ; 
 CHC <=  IAK & TAH  |  IBK & TBH  |  ICK & TCH  |  IDK & TDH  ; 
 CHK <=  IAK & TAH  |  IBK & TBH  |  ICK & TCH  |  IDK & TDH  ; 
 aak <= iak ; 
 abk <= ibk ; 
 adk <= idk ; 
 DPC <=  JGA & jgg  |  jga & JGG  |  jga & jgg  |  JGA & JGG  ;
 DQC <=  JHA & jhg  |  jha & JHG  |  jha & jhg  |  JHA & JHG  ;
 CIC <=  IAS & TAI  |  IBS & TBI  |  ICS & TCI  |  IDS & TDI  ; 
 aas <= ias ; 
 abs <= ibs ; 
 acs <= ics ; 
 ads <= ids ; 
 OMC <= NAC ; 
 NAC <=  IEC  |  IFC  |  IGC  |  IHC  ; 
 HBC <= HAC ; 
 OIC <= HBC ; 
 OKC <= NSC ; 
 OLC <= NSC ; 
 OHC <=  FAG & GBC & egc  |  fag & EGC  |  gbc & EGC  ; 
 OAC <=  FAA & GAC & eac  |  faa & EAC  |  gac & EAC  ; 
 OEC <=  FAA & GAC & eac  |  faa & EAC  |  gac & EAC  ; 
 OCC <=  FAE & GBC & eec  |  fae & EEC  |  gbc & EEC  ; 
 OGC <=  FAE & GBC & eec  |  fae & EEC  |  gbc & EEC  ; 
 EIC <=  KCA & kcb & kcc  |  kca & KCB & kcc  |  kca & kcb & KCC  |  KCA & KCB & KCC  ;
 HAC <= FCC ; 
 OAK <=  FAB & GAC & ebc  |  fab & EBC  |  gac & EBC  ; 
 OEK <=  FAB & GAC & ebc  |  fab & EBC  |  gac & EBC  ; 
 OCK <=  FAF & GBC & efc  |  faf & EFC  |  gbc & EFC  ; 
 OGK <=  FAF & GBC & efc  |  faf & EFC  |  gbc & EFC  ; 
 EJC <=  KCA & kcb & kcc  |  kca & KCB & kcc  |  kca & kcb & KCC  |  KCA & KCB & KCC  ;
 DIC <= CIC ; 
 OBC <=  FAC & GAC & ecc  |  fac & ECC  |  gac & ECC  ; 
 OFC <=  FAC & GAC & ecc  |  fac & ECC  |  gac & ECC  ; 
 ODC <=  FAG & GBC & egc  |  fag & EGC  |  gbc & EGC  ; 
 EKC <=  KCA & kcb & kcd  |  kca & KCB & kcd  |  kca & kcb & KCD  |  KCA & KCB & KCD  ;
 OBK <=  FAD & GAC & edc  |  fad & EDC  |  gac & EDC  ; 
 ODK <=  FAH & GBC & ehc  |  fah & EHC  |  gbc & EHC  ; 
 OHK <=  FAH & GBC & ehc  |  fah & EHC  |  gbc & EHC  ; 
 BAD <= AAD ; 
 BBD <= ABD ; 
 BCD <= ACD ; 
 BDD <= ADD ; 
 BAL <= AAL ; 
 BBL <= ABL ; 
 BCL <= ACL ; 
 BDL <= ADL ; 
 BBT <= ABT ; 
 BCT <= ACT ; 
 BDT <= ADT ; 
 NBD <= NAD ; 
 NCD <= NBD ; 
 NDD <= NCD ; 
 NED <= NDD ; 
 NFD <= NED ; 
 NGD <= NFD ; 
 NHD <= NGD ; 
 NID <= NHD ; 
 NJD <= NID ; 
 NKD <= NJD ; 
 NLD <= NKD ; 
 NMD <= NLD ; 
 NND <= NMD ; 
 NOD <= NND ; 
 NPD <= NOD ; 
 NQD <= NPD ; 
 DAD <= CAL ; 
 DDD <= CDL ; 
 ECD <= DCD ; 
 EDD <= DDD ; 
 DED <= CEL ; 
 EED <= DED ; 
 DGD <= CGL ; 
 DHD <= CHL ; 
 EGD <= DGD ; 
 CDD <=  AAD & TAD  |  ABD & TBD  |  ACD & TCD  |  ADD & TDD  ; 
 CDL <=  AAD & TAD  |  ABD & TBD  |  ACD & TCD  |  ADD & TDD  ; 
 DMD <=  JDB & jdf  |  jdb & JDF  |  jdb & jdf  |  JDB & JDF  ;
 CED <=  AAL & TAE  |  ABL & TBE  |  ACL & TCE  |  ADL & TDE  ; 
 CEL <=  AAL & TAE  |  ABL & TBE  |  ACL & TCE  |  ADL & TDE  ; 
 DND <=  JEB & jef  |  jeb & JEF  |  jeb & jef  |  JEB & JEF  ;
 CFD <=  AAT & TAF  |  ABT & TBF  |  ACT & TCF  |  ADT & TDF  ; 
 CFL <=  AAT & TAF  |  ABT & TBF  |  ACT & TCF  |  ADT & TDF  ; 
 DOD <=  JFB & jff  |  jfb & JFF  |  jfb & jff  |  JFB & JFF  ;
 NRD <= NQD ; 
 NSD <= NRD ; 
 PSD <= NRD ; 
 CAD <=  BAD & TAA  |  BBD & TBA  |  BCD & TCA  |  BDD & TDA  ; 
 CAL <=  BAD & TAA  |  BBD & TBA  |  BCD & TCA  |  BDD & TDA  ; 
 DJD <=  JAB & jaf  |  jab & JAF  |  jab & jaf  |  JAB & JAF  ;
 CBD <=  BAL & TAB  |  BBL & TBB  |  BCL & TCB  |  BDL & TDB  ; 
 CBL <=  BAL & TAB  |  BBL & TBB  |  BCL & TCB  |  BDL & TDB  ; 
 DKD <=  JBB & jbf  |  jbb & JBF  |  jbb & jbf  |  JBB & JBF  ;
 CCD <=  BAT & TAC  |  BBT & TBC  |  BCT & TCC  |  BDT & TDC  ; 
 CCL <=  BAT & TAC  |  BBT & TBC  |  BCT & TCC  |  BDT & TDC  ; 
 DLD <=  JCB & jcf  |  jcb & JCF  |  jcb & jcf  |  JCB & JCF  ;
 CGD <=  IAD & TAG  |  IBD & TBG  |  ICD & TCG  |  IDD & TDG  ; 
 CGL <=  IAD & TAG  |  IBD & TBG  |  ICD & TCG  |  IDD & TDG  ; 
 aad <= iad ; 
 abd <= ibd ; 
 acd <= icd ; 
 add <= idd ; 
 CHD <=  IAL & TAH  |  IBL & TBH  |  ICL & TCH  |  IDL & TDH  ; 
 CHL <=  IAL & TAH  |  IBL & TBH  |  ICL & TCH  |  IDL & TDH  ; 
 aal <= ial ; 
 abl <= ibl ; 
 acl <= icl ; 
 adl <= idl ; 
 DPD <=  JGB & jgf  |  jgb & JGF  |  jgb & jgf  |  JGB & JGF  ;
 DQD <=  JHB & jhf  |  jhb & JHF  |  jhb & jhf  |  JHB & JHF  ;
 CID <=  IAT & TAI  |  IBT & TBI  |  ICT & TCI  |  IDT & TDI  ; 
 aat <= iat ; 
 abt <= ibt ; 
 act <= ict ; 
 adt <= idt ; 
 NAD <=  IED  |  IFD  |  IGD  |  IHD  ; 
 PAD <=  IED  |  IFD  |  IGD  |  IHD  ; 
 HBD <= HAD ; 
 OID <= HBD ; 
 OKD <= NSD ; 
 OLD <= NSD ; 
 OHD <=  FAG & GBD & egd  |  fag & EGD  |  gbd & EGD  ; 
 OAD <=  FAA & GAD & ead  |  faa & EAD  |  gad & EAD  ; 
 OED <=  FAA & GAD & ead  |  faa & EAD  |  gad & EAD  ; 
 OCD <=  FAE & GBD & eed  |  fae & EED  |  gbd & EED  ; 
 OGD <=  FAE & GBD & eed  |  fae & EED  |  gbd & EED  ; 
 EID <=  KDA & kdb & kdc  |  kda & KDB & kdc  |  kda & kdb & KDC  |  KDA & KDB & KDC  ;
 HAD <= FCD ; 
 OAL <=  FAB & GAD & ebd  |  fab & EBD  |  gad & EBD  ; 
 OEL <=  FAB & GAD & ebd  |  fab & EBD  |  gad & EBD  ; 
 OCL <=  FAF & GBD & efd  |  faf & EFD  |  gbd & EFD  ; 
 OGL <=  FAF & GBD & efd  |  faf & EFD  |  gbd & EFD  ; 
 EJD <=  KDA & kdb & kdc  |  kda & KDB & kdc  |  kda & kdb & KDC  |  KDA & KDB & KDC  ;
 DID <= CID ; 
 OBD <=  FAC & GAD & ecd  |  fac & ECD  |  gad & ECD  ; 
 OFD <=  FAC & GAD & ecd  |  fac & ECD  |  gad & ECD  ; 
 ODD <=  FAG & GBD & egd  |  fag & EGD  |  gbd & EGD  ; 
 EKD <=  KDA & kdb & kdd  |  kda & KDB & kdd  |  kda & kdb & KDD  |  KDA & KDB & KDD  ;
 OBL <=  FAD & GAD & edd  |  fad & EDD  |  gad & EDD  ; 
 OFL <=  FAD & GAD & edd  |  fad & EDD  |  gad & EDD  ; 
 ODL <=  FAH & GBD & ehd  |  fah & EHD  |  gbd & EHD  ; 
 OHL <=  FAH & GBD & ehd  |  fah & EHD  |  gbd & EHD  ; 
 CDH <=  AAH & TAD  |  ABH & TBD  |  ACH & TCD  |  ADH & TDD  ; 
 BAE <= AAE ; 
 BBE <= ABE ; 
 BCE <= ACE ; 
 BDE <= ADE ; 
 CEM <=  AAM & TAE  |  ABM & TBE  |  ACM & TCE  |  ADM & TDE  ; 
 BAM <= AAM ; 
 BBM <= ABM ; 
 BCM <= ACM ; 
 BDM <= ADM ; 
 BAU <= AAU ; 
 BBU <= ABU ; 
 BCU <= ACU ; 
 BDU <= ADU ; 
 NBE <= NAE ; 
 NCE <= NBE ; 
 NDE <= NCE ; 
 NEE <= NDE ; 
 NFE <= NEE ; 
 NGE <= NFE ; 
 NHE <= NGE ; 
 NIE <= NHE ; 
 NJE <= NIE ; 
 NKE <= NJE ; 
 NLE <= NKE ; 
 NME <= NLE ; 
 NNE <= NME ; 
 NOE <= NNE ; 
 NPE <= NOE ; 
 NQE <= NPE ; 
 DAE <= CAM ; 
 DBE <= CBM ; 
 EAE <= DAE ; 
 EBE <= DBE ; 
 DCE <= CCM ; 
 DDE <= CDM ; 
 EDE <= DDE ; 
 ECE <= DCE ; 
 DEE <= CEM ; 
 DFE <= CFM ; 
 EEE <= DEE ; 
 EFE <= DFE ; 
 DGE <= CGM ; 
 DHE <= CHM ; 
 EGE <= DGE ; 
 EHE <= DHE ; 
 CDE <=  AAE & TAD  |  ABE & TBD  |  ACE & TCD  |  ADE & TDD  ; 
 CDM <=  AAE & TAD  |  ABE & TBD  |  ACE & TCD  |  ADE & TDD  ; 
 DME <=  JDA & jdb & jdc  |  jda & JDB & jdc  |  jda & jdb & JDC  |  JDA & JDB & JDC  ;
 CEE <=  AAM & TAE  |  ABM & TBE  |  ACM & TCE  |  ADM & TDE  ; 
 DNE <=  JEA & jeb & jec  |  jea & JEB & jec  |  jea & jeb & JEC  |  JEA & JEB & JEC  ;
 CFE <=  AAU & TAF  |  ABU & TBF  |  ACU & TCF  |  ADU & TDF  ; 
 CFM <=  AAU & TAF  |  ABU & TBF  |  ACU & TCF  |  ADU & TDF  ; 
 DOE <=  JFA & jfb & jfc  |  jfa & JFB & jfc  |  jfa & jfb & JFC  |  JFA & JFB & JFC  ;
 NRE <= NQE ; 
 NSE <= NRE ; 
 PSE <= NRE ; 
 PCC <=  DOE & dke  |  doe & DKE  ; 
 CAE <=  BAE & TAA  |  BBE & TBA  |  BCE & TCA  |  BDE & TDA  ; 
 CAM <=  BAE & TAA  |  BBE & TBA  |  BCE & TCA  |  BDE & TDA  ; 
 DJE <=  JAA & jab & jac  |  jaa & JAB & jac  |  jaa & jab & JAC  |  JAA & JAB & JAC  ;
 CBE <=  BAM & TAB  |  BBM & TBB  |  BCM & TCB  |  BDM & TDB  ; 
 CBM <=  BAM & TAB  |  BBM & TBB  |  BCM & TCB  |  BDM & TDB  ; 
 DKE <=  JBA & jbb & jbc  |  jba & JBB & jbc  |  jba & jbb & JBC  |  JBA & JBB & JBC  ;
 CCE <=  BAU & TAC  |  BBU & TBC  |  BCU & TCC  |  BDU & TDC  ; 
 CCM <=  BAU & TAC  |  BBU & TBC  |  BCU & TCC  |  BDU & TDC  ; 
 DLE <=  JCA & jcb & jcc  |  jca & JCB & jcc  |  jca & jcb & JCC  |  JCA & JCB & JCC  ;
 CGE <=  IAE & TAG  |  IBE & TBG  |  ICE & TCG  |  IDE & TDG  ; 
 CGM <=  IAE & TAG  |  IBE & TBG  |  ICE & TCG  |  IDE & TDG  ; 
 aae <= iae ; 
 abe <= ibe ; 
 ace <= ice ; 
 ade <= ide ; 
 CHE <=  IAM & TAH  |  IBM & TBH  |  ICM & TCH  |  IDM & TDH  ; 
 CHM <=  IAM & TAH  |  IBM & TBH  |  ICM & TCH  |  IDM & TDH  ; 
 aam <= iam ; 
 abm <= ibm ; 
 acm <= icm ; 
 adm <= idm ; 
 DPE <=  JGA & jgb & jgc  |  jga & JGB & jgc  |  jga & jgb & JGC  |  JGA & JGB & JGC  ;
 DQE <=  JHA & jhb & jhc  |  jha & JHB & jhc  |  jha & jhb & JHC  |  JHA & JHB & JHC  ;
 CIE <=  IAU & TAI  |  IBU & TBI  |  ICU & TCI  |  IDU & TDI  ; 
 aau <= iau ; 
 abu <= ibu ; 
 acu <= icu ; 
 adu <= idu ; 
 OMD <= JIA ; 
 NAE <=  IEE  |  IFE  |  IGE  |  IHE  ; 
 PAE <=  IEE  |  IFE  |  IGE  |  IHE  ; 
 HBE <= HAE ; 
 OIE <= HBE ; 
 OKE <= JIB ; 
 OLE <= JIC ; 
 ODE <=  FBG & GBE & ege  |  fbg & EGE  |  gbe & EGE  ; 
 OAE <=  FBA & GAE & eae  |  fba & EAE  |  gae & EAE  ; 
 OEE <=  FBA & GAE & eae  |  fba & EAE  |  gae & EAE  ; 
 OCE <=  FBE & GBE & eee  |  fbe & EEE  |  gbe & EEE  ; 
 OGE <=  FBE & GBE & eee  |  fbe & EEE  |  gbe & EEE  ; 
 EIE <=  KEA & keb & kec  |  kea & KEB & kec  |  kea & keb & KEC  |  KEA & KEB & KEC  ;
 HAE <= FCE ; 
 OAM <=  FBB & GAE & ebe  |  fbb & EBE  |  gae & EBE  ; 
 OEM <=  FBB & GAE & ebe  |  fbb & EBE  |  gae & EBE  ; 
 OCM <=  FBF & GBE & efe  |  fbf & EFE  |  gbe & EFE  ; 
 OGM <=  FBF & GBE & efe  |  fbf & EFE  |  gbe & EFE  ; 
 EJE <=  KEA & keb & kec  |  kea & KEB & kec  |  kea & keb & KEC  |  KEA & KEB & KEC  ;
 DIE <= CIE ; 
 OBE <=  FBC & GAE & ece  |  fbc & ECE  |  gae & ECE  ; 
 OFE <=  FBC & GAE & ece  |  fbc & ECE  |  gae & ECE  ; 
 OHE <=  FBG & GBE & ege  |  fbg & EGE  |  gbe & EGE  ; 
 EKE <=  KEA & keb & ked  |  kea & KEB & ked  |  kea & keb & KED  |  KEA & KEB & KED  ;
 OBM <=  FBD & GAE & ede  |  fbd & EDE  |  gae & EDE  ; 
 OFM <=  FBD & GAE & ede  |  fbd & EDE  |  gae & EDE  ; 
 ODM <=  FBH & GBE & ehe  |  fbh & EHE  |  gbe & EHE  ; 
 OHM <=  FBH & GBE & ehe  |  fbh & EHE  |  gbe & EHE  ; 
 BAF <= AAF ; 
 BBF <= ABF ; 
 BCF <= ACF ; 
 BDF <= ADF ; 
 DCF <= CCN ; 
 BAN <= AAN ; 
 BBN <= ABN ; 
 BCN <= ACN ; 
 BDN <= ADN ; 
 BAV <= AAV ; 
 BBV <= ABV ; 
 BCV <= ACV ; 
 BDV <= ADV ; 
 NBF <= NAF ; 
 NCF <= NBF ; 
 NDF <= NCF ; 
 NEF <= NDF ; 
 NFF <= NEF ; 
 NGF <= NFF ; 
 NHF <= NGF ; 
 NIF <= NHF ; 
 NJF <= NIF ; 
 NKF <= NJF ; 
 NLF <= NKF ; 
 NMF <= NLF ; 
 NNF <= NMF ; 
 NOF <= NNF ; 
 NPF <= NOF ; 
 NQF <= NPF ; 
 DAF <= CAN ; 
 DBF <= CBN ; 
 EAF <= DAF ; 
 EBF <= DBF ; 
 DDF <= CDN ; 
 ECF <= DCF ; 
 EDF <= DDF ; 
 DEF <= CEN ; 
 DFF <= CFN ; 
 EEF <= DEF ; 
 EFF <= DFF ; 
 DGF <= CGN ; 
 DHF <= CHN ; 
 EGF <= DGF ; 
 EHF <= DHF ; 
 CDF <=  AAF & TAD  |  ABF & TBD  |  ACF & TCD  |  ADF & TDD  ; 
 CDN <=  AAF & TAD  |  ABF & TBD  |  ACF & TCD  |  ADF & TDD  ; 
 CEF <=  AAN & TAE  |  ABN & TBE  |  ACN & TCE  |  ADN & TDE  ; 
 CEN <=  AAN & TAE  |  ABN & TBE  |  ACN & TCE  |  ADN & TDE  ; 
 CFF <=  AAV & TAF  |  ABV & TBF  |  ACV & TCF  |  ADV & TDF  ; 
 CFN <=  AAV & TAF  |  ABV & TBF  |  ACV & TCF  |  ADV & TDF  ; 
 NRF <= NQF ; 
 NSF <= NRF ; 
 PSF <= NRF ; 
 CAF <=  BAF & TAA  |  BBF & TBA  |  BCF & TCA  |  BDF & TDA  ; 
 CAN <=  BAF & TAA  |  BBF & TBA  |  BCF & TCA  |  BDF & TDA  ; 
 CBF <=  BAN & TAB  |  BBN & TBB  |  BCN & TCB  |  BDN & TDB  ; 
 CBN <=  BAN & TAB  |  BBN & TBB  |  BCN & TCB  |  BDN & TDB  ; 
 CCF <=  BAV & TAC  |  BBV & TBC  |  BCV & TCC  |  BDV & TDC  ; 
 CCN <=  BAV & TAC  |  BBV & TBC  |  BCV & TCC  |  BDV & TDC  ; 
 CGF <=  IAF & TAG  |  IBF & TBG  |  ICF & TCG  |  IDF & TDG  ; 
 CGN <=  IAF & TAG  |  IBF & TBG  |  ICF & TCG  |  IDF & TDG  ; 
 aaf <= iaf ; 
 abf <= ibf ; 
 acf <= icf ; 
 adf <= idf ; 
 aan <= ian ; 
 abn <= ibn ; 
 acn <= icn ; 
 adn <= idn ; 
 CHF <=  IAN & TAH  |  IBN & TBH  |  ICN & TCH  |  IDN & TDH  ; 
 CHN <=  IAN & TAH  |  IBN & TBH  |  ICN & TCH  |  IDN & TDH  ; 
 OEN <=  FBB & GAF & ebf  |  fbb & EBF  |  gaf & EBF  ; 
 DIF <=  CIF  |  CIF  ;
 CIF <=  IAV & TAI  |  IBV & TBI  |  ICV & TCI  |  IDV & TDI  ; 
 aav <= iav ; 
 abv <= ibv ; 
 acv <= icv ; 
 adv <= idv ; 
 NAF <=  IEF  |  IFFF   |  IGF  |  IHF  ; 
 PAF <=  IEF  |  IFFF   |  IGF  |  IHF  ; 
 HBF <= HAF ; 
 OIF <= HBF ; 
 ONC <= JIE ; 
 OOC <= JID ; 
 OAF <=  FBA & GAF & eaf  |  fba & EAF  |  gaf & EAF  ; 
 OEF <=  FBA & GAF & eaf  |  fba & EAF  |  gaf & EAF  ; 
 OCF <=  FBE & GBF & eef  |  fbe & EEF  |  gbf & EEF  ; 
 OGF <=  FBE & GBF & eef  |  fbe & EEF  |  gbf & EEF  ; 
 EIF <=  KFA & kfb & kfc  |  kfa & KFB & kfc  |  kfa & kfb & KFC  |  KFA & KFB & KFC  ;
 HAF <= FCF ; 
 OAN <=  FBB & GAF & ebf  |  fbb & EBF  |  gaf & EBF  ; 
 OCN <=  FBF & GBF & eff  |  fbf & EFF  |  gbf & EFF  ; 
 OGN <=  FBF & GBF & eff  |  fbf & EFF  |  gbf & EFF  ; 
 EJF <=  KFA & kfb & kfc  |  kfa & KFB & kfc  |  kfa & kfb & KFC  |  KFA & KFB & KFC  ;
 OBF <=  FBC & GAF & ecf  |  fbc & ECF  |  gaf & ECF  ; 
 OFF <=  FBC & GAF & ecf  |  fbc & ECF  |  gaf & ECF  ; 
 ODF <=  FBG & GBF & egf  |  fbg & EGF  |  gbf & EGF  ; 
 OHF <=  FBG & GBF & egf  |  fbg & EGF  |  gbf & EGF  ; 
 EKF <=  KFA & kfb & kfd  |  kfa & KFB & kfd  |  kfa & kfb & KFD  |  KFA & KFB & KFD  ;
 OBN <=  FBD & GAF & edf  |  fbd & EDF  |  gaf & EDF  ; 
 OFN <=  FBD & GAF & edf  |  fbd & EDF  |  gaf & EDF  ; 
 ODN <=  FBH & GBF & ehf  |  fbh & EHF  |  gbf & EHF  ; 
 OHN <=  FBH & GBF & ehf  |  fbh & EHF  |  gbf & EHF  ; 
 BAG <= AAG ; 
 BBG <= ABG ; 
 BCG <= ACG ; 
 BDG <= ADG ; 
 BAO <= AAO ; 
 BBO <= ABO ; 
 BCO <= ACO ; 
 BDO <= ADO ; 
 BAW <= AAW ; 
 BBW <= ABW ; 
 BCW <= ACW ; 
 BDW <= ADW ; 
 DAG <= CAO ; 
 DBG <= CBO ; 
 EAG <= DAG ; 
 EBG <= DBG ; 
 DCG <= CCO ; 
 DDG <= CDO ; 
 ECG <= DCG ; 
 EDG <= DDG ; 
 DEG <= CEO ; 
 DFG <= CFO ; 
 EEG <= DEG ; 
 EFG <= DFG ; 
 DGG <= CGO ; 
 DHG <= CHO ; 
 EGG <= DGG ; 
 EHG <= DHG ; 
 CDG <=  AAG & TAD  |  ABG & TBD  |  ACG & TCD  |  ADG & TDD  ; 
 CDO <=  AAG & TAD  |  ABG & TBD  |  ACG & TCD  |  ADG & TDD  ; 
 abc <= ibc ; 
 CEG <=  AAO & TAE  |  ABO & TBE  |  ACO & TCE  |  ADO & TDE  ; 
 CEO <=  AAO & TAE  |  ABO & TBE  |  ACO & TCE  |  ADO & TDE  ; 
 CFG <=  AAW & TAF  |  ABW & TBF  |  ACW & TCF  |  ADW & TDF  ; 
 CFO <=  AAW & TAF  |  ABW & TBF  |  ACW & TCF  |  ADW & TDF  ; 
 CBG <=  BAO & TAB  |  BBO & TBB  |  BCO & TCB  |  BDO & TDB  ; 
 LAA <=  FCA & fcb & fcc  |  fca & FCB & fcc  |  fca & fcb & FCC  |  FCA & FCB & FCC  ;
 lba <=  FCA & fcb & fcc  |  fca & FCB & fcc  |  fca & fcb & FCC  |  fca & fcb & fcc  ;
 CAG <=  BAG & TAA  |  BBG & TBA  |  BCG & TCA  |  BDG & TDA  ; 
 CAO <=  BAG & TAA  |  BBG & TBA  |  BCG & TCA  |  BDG & TDA  ; 
 CBO <=  BAO & TAB  |  BBO & TBB  |  BCO & TCB  |  BDO & TDB  ; 
 OPA <=  JPA & jqd  |  jpa & JQA  |  jpa & JQB  |  jpa & JQC  ; 
 CCG <=  BAW & TAC  |  BBW & TBC  |  BCW & TCC  |  BDW & TDC  ; 
 CCO <=  BAW & TAC  |  BBW & TBC  |  BCW & TCC  |  BDW & TDC  ; 
 CGG <=  IAG & TAG  |  IBG & TBG  |  ICG & TCG  |  IDG & TDG  ; 
 CGO <=  IAG & TAG  |  IBG & TBG  |  ICG & TCG  |  IDG & TDG  ; 
 aag <= iag ; 
 abg <= ibg ; 
 acg <= icg ; 
 adg <= idg ; 
 CHG <=  IAO & TAH  |  IBO & TBH  |  ICO & TCH  |  IDO & TDH  ; 
 CHO <=  IAO & TAH  |  IBO & TBH  |  ICO & TCH  |  IDO & TDH  ; 
 aao <= iao ; 
 abo <= ibo ; 
 aco <= ico ; 
 ado <= ido ; 
 CIG <=  IAW & TAI  |  IBW & TBI  |  ICW & TCI  |  IDW & TDI  ; 
 aaw <= iaw ; 
 abw <= ibw ; 
 acw <= icw ; 
 adw <= idw ; 
 LAB <=  FCD & fce & fcf  |  fcd & FCE & fcf  |  fcd & fce & FCF  |  FCD & FCE & FCF  ;
 lbb <=  FCD & fce & fcf  |  fcd & FCE & fcf  |  fcd & fce & FCF  |  fcd & fce & fcf  ;
 LAC <=  FCG & fch  |  fcg & FCH  |  fcg & fch  |  FCG & FCH  ;
 lbc <=  FCG & fch  |  fcg & FCH  |  fcg & fch  |  fcg & fch  ;
 OJA <=  MAA  ; 
 ojb <=  MAA  |  mab & mac  ; 
 HBG <= HAG ; 
 OIG <= HBG ; 
 ONA <= NSA ; 
 OOA <= NSA ; 
 OAG <=  FBA & GAG & eag  |  fba & EAG  |  gag & EAG  ; 
 OEG <=  FBA & GAG & eag  |  fba & EAG  |  gag & EAG  ; 
 OCG <=  FBE & GBG & eeg  |  fbe & EEG  |  gbg & EEG  ; 
 OGG <=  FBE & GBG & eeg  |  fbe & EEG  |  gbg & EEG  ; 
 EIG <=  KGA & kgb & kgc  |  kga & KGB & kgc  |  kga & kgb & KGC  |  KGA & KGB & KGC  ;
 HAG <= FCG ; 
 OAO <=  FBB & GAG & ebg  |  fbb & EBG  |  gag & EBG  ; 
 OEO <=  FBB & GAG & ebg  |  fbb & EBG  |  gag & EBG  ; 
 OCO <=  FBF & GBG & efg  |  fbf & EFG  |  gbg & EFG  ; 
 OGO <=  FBF & GBG & efg  |  fbf & EFG  |  gbg & EFG  ; 
 EJG <=  KGA & kgb & kgc  |  kga & KGB & kgc  |  kga & kgb & KGC  |  KGA & KGB & KGC  ;
 DIG <= CIG ; 
 OBG <=  FBC & GAG & ecg  |  fbc & ECG  |  gag & ECG  ; 
 OFG <=  FBC & GAG & ecg  |  fbc & ECG  |  gag & ECG  ; 
 ODG <=  FBG & GBG & egg  |  fbg & EGG  |  gbg & EGG  ; 
 OHG <=  FBG & GBG & egg  |  fbg & EGG  |  gbg & EGG  ; 
 EKG <=  KGA & kgb & kgd  |  kga & KGB & kgd  |  kga & kgb & KGD  |  KGA & KGB & KGD  ;
 OBO <=  FBD & GAG & edg  |  fbd & EDG  |  gag & EDG  ; 
 OFO <=  FBD & GAG & edg  |  fbd & EDG  |  gag & EDG  ; 
 ODO <=  FBH & GBG & ehg  |  fbh & EHG  |  gbg & EHG  ; 
 OHO <=  FBH & GBG & ehg  |  fbh & EHG  |  gbg & EHG  ; 
 BAH <= AAH ; 
 BBH <= ABH ; 
 BCH <= ACH ; 
 BDH <= ADH ; 
 BAP <= AAP ; 
 BBP <= ABP ; 
 BCP <= ACP ; 
 BDP <= ADP ; 
 BAX <= AAX ; 
 BBX <= ABX ; 
 BCX <= ACX ; 
 BDX <= ADX ; 
 DAH <= CAP ; 
 DBH <= CBP ; 
 EAH <= DAH ; 
 EBH <= DBH ; 
 DCH <= CCP ; 
 DDH <= CDP ; 
 ECH <= DCH ; 
 EDH <= DDH ; 
 DEH <= CEP ; 
 DFH <= CFP ; 
 EEH <= DEH ; 
 EFH <= DFH ; 
 DGH <= CGP ; 
 DHH <= CHP ; 
 EGH <= DGH ; 
 EHH <= DHH ; 
 CDP <=  AAH & TAD  |  ABH & TBD  |  ACH & TCD  |  ADH & TDD  ; 
 CEH <=  AAP & TAE  |  ABP & TBE  |  ACP & TCE  |  ADP & TDE  ; 
 CEP <=  AAP & TAE  |  ABP & TBE  |  ACP & TCE  |  ADP & TDE  ; 
 CFH <=  AAX & TAF  |  ABX & TBF  |  ACX & TCF  |  ADX & TDF  ; 
 CBH <=  AAX & TAF  |  ABX & TBF  |  ACX & TCF  |  ADX & TDF  ; 
 TAD <= QAD ; 
 TBD <= QAA ; 
 TCD <= QAB ; 
 TDD <= QAC ; 
 TAE <= QAD ; 
 TBE <= QAA ; 
 TCE <= QAB ; 
 TDE <= QAC ; 
 TAF <= QAD ; 
 TBF <= QAA ; 
 TCF <= QAB ; 
 TDF <= QAC ; 
 TAI <= QAD ; 
 TBI <= QAA ; 
 TCI <= QAB ; 
 TDI <= QAC ; 
 TAC <= QAD ; 
 TCC <= QAB ; 
 TDC <= QAC ; 
 TAB <= QAD ; 
 TBB <= QAA ; 
 TCB <= QAB ; 
 TDB <= QAC ; 
 TAA <= QAD ; 
 TBA <= QAA ; 
 TCA <= QAB ; 
 TDA <= QAC ; 
 CAH <=  BAH & TAA  |  BBH & TBA  |  BCH & TCA  |  BDH & TDA  ; 
 CAP <=  BAH & TAA  |  BBH & TBA  |  BCH & TCA  |  BDH & TDA  ; 
 CBP <=  BAP & TAB  |  BBP & TBB  |  BCP & TCB  |  BDP & TDB  ; 
 CCH <=  BAX & TAC  |  BBX & TBC  |  BCX & TCC  |  BDX & TDC  ; 
 CCP <=  BAX & TAC  |  BBX & TBC  |  BCX & TCC  |  BDX & TDC  ; 
 CGH <=  IAH & TAG  |  IBH & TBG  |  ICH & TCG  |  IDH & TDG  ; 
 CGP <=  IAH & TAG  |  IBH & TBG  |  ICH & TCG  |  IDH & TDG  ; 
 aah <= iah ; 
 abh <= ibh ; 
 ach <= ich ; 
 adh <= idh ; 
 jja <=  IJA  ; 
 jjb <=  IJA  ; 
 CHH <=  IAP & TAH  |  IBP & TBH  |  ICP & TCH  |  IDP & TDH  ; 
 CHP <=  IAP & TAH  |  IBP & TBH  |  ICP & TCH  |  IDP & TDH  ; 
 aap <= iap ; 
 abp <= ibp ; 
 acp <= icp ; 
 adp <= idp ; 
 PCA <=  DME & dje & dle  |  dme & DJE & dle  |  dme & dje & DLE  |  DME & DJE & DLE  ;
 CIH <=  IAX & TAI  |  IBX & TBI  |  ICX & TCI  |  IDX & TDI  ; 
 aax <= iax ; 
 abx <= ibx ; 
 acx <= icx ; 
 adx <= idx ; 
 TAH <= QAD ; 
 TBH <= QAA ; 
 TCH <= QAB ; 
 TDH <= QAC ; 
 TAG <= QAD ; 
 TBG <= QAA ; 
 TCG <= QAB ; 
 TDG <= QAC ; 
 QAA <= IIA ; 
 QAB <= QAA ; 
 QAC <= QAB ; 
 QAD <= QAC ; 
 HBH <= HAH ; 
 OIH <= HBH ; 
 ONB <= NSB ; 
 OOB <= NSB ; 
 OHH <=  FBG & GBH & egh  |  fbg & EGH  |  gbh & EGH  ; 
 OAH <=  FBA & GAH & eah  |  fba & EAH  |  gah & EAH  ; 
 OEH <=  FBA & GAH & eah  |  fba & EAH  |  gah & EAH  ; 
 OCH <=  FBE & GBH & eeh  |  fbe & EEH  |  gbh & EEH  ; 
 OGH <=  FBE & GBH & eeh  |  fbe & EEH  |  gbh & EEH  ; 
 EIH <=  KHA & khb & khc  |  kha & KHB & khc  |  kha & khb & KHC  |  KHA & KHB & KHC  ;
 HAH <= FCH ; 
 OAP <=  FBB & GAH & ebh  |  fbb & EBH  |  gah & EBH  ; 
 OEP <=  FBB & GAH & ebh  |  fbb & EBH  |  gah & EBH  ; 
 OCP <=  FBF & GBH & efh  |  fbf & EFH  |  gbh & EFH  ; 
 OGP <=  FBF & GBH & efh  |  fbf & EFH  |  gbh & EFH  ; 
 EJH <=  KHA & khb & khc  |  kha & KHB & khc  |  kha & khb & KHC  |  KHA & KHB & KHC  ;
 DIH <= CIH ; 
 OBH <=  FBC & GAH & ech  |  fbc & ECH  |  gah & ECH  ; 
 OFH <=  FBC & GAH & ech  |  fbc & ECH  |  gah & ECH  ; 
 ODH <=  FBG & GBH & egh  |  fbg & EGH  |  gbh & EGH  ; 
 EKH <=  KHA & khb & khd  |  kha & KHB & khd  |  kha & khb & KHD  |  KHA & KHB & KHD  ;
 OBP <=  FBD & GAH & edh  |  fbd & EDH  |  gah & EDH  ; 
 OFP <=  FBD & GAH & edh  |  fbd & EDH  |  gah & EDH  ; 
 ODP <=  FBH & GBH & ehh  |  fbh & EHH  |  gbh & EHH  ; 
 OHP <=  FBH & GBH & ehh  |  fbh & EHH  |  gbh & EHH  ; 
end
endmodule;
