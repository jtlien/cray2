module tf( IZZ,
 IAA, 
 IAB, 
 IAC, 
 IAD, 
 IAE, 
 IAF, 
 IAG, 
 IAH, 
 IAI, 
 IAJ, 
 IAK, 
 IAL, 
 IAM, 
 IAN, 
 IAO, 
 IAP, 
 IBA, 
 IBB, 
 IBC, 
 IBD, 
 IBE, 
 IBF, 
 IBG, 
 IBH, 
 IBI, 
 IBJ, 
 IBK, 
 IBL, 
 IBM, 
 IBN, 
 IBO, 
 IBP, 
 ICA, 
 ICB, 
 ICC, 
 ICD, 
 ICE, 
 ICF, 
 ICG, 
 ICH, 
 ICI, 
 ICJ, 
 ICK, 
 ICL, 
 ICM, 
 ICN, 
 ICO, 
 ICP, 
 IDA, 
 IDB, 
 IDC, 
 IDD, 
 IDE, 
 IDF, 
 IDG, 
 IDH, 
 IDI, 
 IDJ, 
 IDK, 
 IDL, 
 IDM, 
 IDN, 
 IDO, 
 IDP, 
 IEA, 
 IEB, 
 IEC, 
 IED, 
 IEE, 
 IEF, 
 IEG, 
 IEH, 
 IEI, 
 IEJ, 
 IEK, 
 IEL, 
 IEM, 
 IEN, 
 IEO, 
 IEP, 
 IFA, 
 IFB, 
 IFC, 
 IFD, 
 IFE, 
 IFFF , 
 IFG, 
 IFH, 
 IFI, 
 IFJ, 
 IFK, 
 IFL, 
 IFM, 
 IFN, 
 IFO, 
 IFP, 
 IGA, 
 IGB, 
 IGC, 
 IGD, 
 IGE, 
 IGF, 
 IGG, 
 IGH, 
 IGI, 
 IGJ, 
 IGK, 
 IGL, 
 IGM, 
 IGN, 
 IGO, 
 IGP, 
 IHA, 
 IHB, 
 IHC, 
 IHD, 
 IHE, 
 IHF, 
 IHG, 
 IHH, 
 IHI, 
 IHJ, 
 IHK, 
 IHL, 
 IHM, 
 IHN, 
 IHO, 
 IHP, 
 IIA, 
 IIB, 
 IIC, 
 IID, 
 IIE, 
 IIF, 
 IJA, 
 IJB, 
 IJC, 
 IJD, 
 IJE, 
 IJF, 
 IJG, 
 IJH, 
 IKA, 
 IKB, 
 IKC, 
 IKD, 
 IKE, 
 IKF, 
 IKG, 
 IKH, 
 IKI, 
 IKJ, 
 IKK, 
 IKM, 
 IKN, 
 IKO, 
 IKP, 
 IKQ, 
 IKR, 
 IKS, 
 IKT, 
 IKU, 
 ILA, 
 OAA, 
 OAB, 
 OAC, 
 OAD, 
 OAE, 
 OAF, 
 OAG, 
 OAH, 
 OAI, 
 OAJ, 
 OAK, 
 OAL, 
 OAM, 
 OAN, 
 OBA, 
 OBB, 
 OBC, 
 OBD, 
 OBE, 
 OBF, 
 OBG, 
 OBH, 
 OBI, 
 OBJ, 
 OBK, 
 OBL, 
 OBM, 
 OBN, 
 OCA, 
 OCB, 
 OCC, 
 OCD, 
 OCE, 
 OCF, 
 OCG, 
 OCH, 
 OCI, 
 OCJ, 
 OCK, 
 OCL, 
 OCM, 
 OCN, 
 ODA, 
 ODB, 
 ODC, 
 ODD, 
 ODE, 
 ODF, 
 ODG, 
 ODH, 
 ODI, 
 ODJ, 
 ODK, 
 ODL, 
 ODM, 
 ODN, 
 OEA, 
 OEB, 
 OEC, 
 OED, 
 OEE, 
 OEF, 
 OEG, 
 OEH, 
 OEI, 
 OEJ, 
 OEK, 
 OEL, 
 OEM, 
 OEN, 
 OEO, 
 OEP, 
 OEQ, 
 OER, 
 OES, 
 OET, 
 OEU, 
 OEV, 
 OEW, 
 OEX, 
 OFA, 
 OFB, 
 OFC, 
 OFD, 
 OHA, 
 OHB, 
 OHC, 
 OHD, 
 OHE, 
 OIA, 
 OIB, 
 OIC, 
 OID, 
 OIE, 
 OIF, 
 OIG, 
 OIH, 
 OKA, 
 OLA, 
 OLB, 
 OLC, 
OLD ); 
    
 input IZZ; 
 input IAA; 
 input IAB; 
 input IAC; 
 input IAD; 
 input IAE; 
 input IAF; 
 input IAG; 
 input IAH; 
 input IAI; 
 input IAJ; 
 input IAK; 
 input IAL; 
 input IAM; 
 input IAN; 
 input IAO; 
 input IAP; 
 input IBA; 
 input IBB; 
 input IBC; 
 input IBD; 
 input IBE; 
 input IBF; 
 input IBG; 
 input IBH; 
 input IBI; 
 input IBJ; 
 input IBK; 
 input IBL; 
 input IBM; 
 input IBN; 
 input IBO; 
 input IBP; 
 input ICA; 
 input ICB; 
 input ICC; 
 input ICD; 
 input ICE; 
 input ICF; 
 input ICG; 
 input ICH; 
 input ICI; 
 input ICJ; 
 input ICK; 
 input ICL; 
 input ICM; 
 input ICN; 
 input ICO; 
 input ICP; 
 input IDA; 
 input IDB; 
 input IDC; 
 input IDD; 
 input IDE; 
 input IDF; 
 input IDG; 
 input IDH; 
 input IDI; 
 input IDJ; 
 input IDK; 
 input IDL; 
 input IDM; 
 input IDN; 
 input IDO; 
 input IDP; 
 input IEA; 
 input IEB; 
 input IEC; 
 input IED; 
 input IEE; 
 input IEF; 
 input IEG; 
 input IEH; 
 input IEI; 
 input IEJ; 
 input IEK; 
 input IEL; 
 input IEM; 
 input IEN; 
 input IEO; 
 input IEP; 
 input IFA; 
 input IFB; 
 input IFC; 
 input IFD; 
 input IFE; 
 input IFFF ; 
 input IFG; 
 input IFH; 
 input IFI; 
 input IFJ; 
 input IFK; 
 input IFL; 
 input IFM; 
 input IFN; 
 input IFO; 
 input IFP; 
 input IGA; 
 input IGB; 
 input IGC; 
 input IGD; 
 input IGE; 
 input IGF; 
 input IGG; 
 input IGH; 
 input IGI; 
 input IGJ; 
 input IGK; 
 input IGL; 
 input IGM; 
 input IGN; 
 input IGO; 
 input IGP; 
 input IHA; 
 input IHB; 
 input IHC; 
 input IHD; 
 input IHE; 
 input IHF; 
 input IHG; 
 input IHH; 
 input IHI; 
 input IHJ; 
 input IHK; 
 input IHL; 
 input IHM; 
 input IHN; 
 input IHO; 
 input IHP; 
 input IIA; 
 input IIB; 
 input IIC; 
 input IID; 
 input IIE; 
 input IIF; 
 input IJA; 
 input IJB; 
 input IJC; 
 input IJD; 
 input IJE; 
 input IJF; 
 input IJG; 
 input IJH; 
 input IKA; 
 input IKB; 
 input IKC; 
 input IKD; 
 input IKE; 
 input IKF; 
 input IKG; 
 input IKH; 
 input IKI; 
 input IKJ; 
 input IKK; 
 input IKM; 
 input IKN; 
 input IKO; 
 input IKP; 
 input IKQ; 
 input IKR; 
 input IKS; 
 input IKT; 
 input IKU; 
 input ILA; 
 output OAA; 
 output OAB; 
 output OAC; 
 output OAD; 
 output OAE; 
 output OAF; 
 output OAG; 
 output OAH; 
 output OAI; 
 output OAJ; 
 output OAK; 
 output OAL; 
 output OAM; 
 output OAN; 
 output OBA; 
 output OBB; 
 output OBC; 
 output OBD; 
 output OBE; 
 output OBF; 
 output OBG; 
 output OBH; 
 output OBI; 
 output OBJ; 
 output OBK; 
 output OBL; 
 output OBM; 
 output OBN; 
 output OCA; 
 output OCB; 
 output OCC; 
 output OCD; 
 output OCE; 
 output OCF; 
 output OCG; 
 output OCH; 
 output OCI; 
 output OCJ; 
 output OCK; 
 output OCL; 
 output OCM; 
 output OCN; 
 output ODA; 
 output ODB; 
 output ODC; 
 output ODD; 
 output ODE; 
 output ODF; 
 output ODG; 
 output ODH; 
 output ODI; 
 output ODJ; 
 output ODK; 
 output ODL; 
 output ODM; 
 output ODN; 
 output OEA; 
 output OEB; 
 output OEC; 
 output OED; 
 output OEE; 
 output OEF; 
 output OEG; 
 output OEH; 
 output OEI; 
 output OEJ; 
 output OEK; 
 output OEL; 
 output OEM; 
 output OEN; 
 output OEO; 
 output OEP; 
 output OEQ; 
 output OER; 
 output OES; 
 output OET; 
 output OEU; 
 output OEV; 
 output OEW; 
 output OEX; 
 output OFA; 
 output OFB; 
 output OFC; 
 output OFD; 
 output OHA; 
 output OHB; 
 output OHC; 
 output OHD; 
 output OHE; 
 output OIA; 
 output OIB; 
 output OIC; 
 output OID; 
 output OIE; 
 output OIF; 
 output OIG; 
 output OIH; 
 output OKA; 
 output OLA; 
 output OLB; 
 output OLC; 
 output OLD; 
  
  
reg  AAA ;
reg  AAB ;
reg  AAC ;
reg  AAD ;
reg  AAE ;
reg  AAF ;
reg  AAG ;
reg  AAH ;
reg  AAI ;
reg  AAJ ;
reg  AAK ;
reg  AAL ;
reg  AAM ;
reg  AAN ;
reg  AAO ;
reg  AAP ;
reg  ABA ;
reg  ABB ;
reg  ABC ;
reg  ABD ;
reg  ABE ;
reg  ABF ;
reg  ABG ;
reg  ABH ;
reg  ABI ;
reg  ABJ ;
reg  ABK ;
reg  ABL ;
reg  ABM ;
reg  ABN ;
reg  ABO ;
reg  ABP ;
reg  ACA ;
reg  ACB ;
reg  ACC ;
reg  ACD ;
reg  ACE ;
reg  ACF ;
reg  ACG ;
reg  ACH ;
reg  ACI ;
reg  ACJ ;
reg  ACK ;
reg  ACL ;
reg  ACM ;
reg  ACN ;
reg  ACO ;
reg  ACP ;
reg  ADA ;
reg  ADB ;
reg  ADC ;
reg  ADD ;
reg  ADE ;
reg  ADF ;
reg  ADG ;
reg  ADH ;
reg  ADI ;
reg  ADJ ;
reg  ADK ;
reg  ADL ;
reg  ADM ;
reg  ADN ;
reg  ADO ;
reg  ADP ;
reg  AEA ;
reg  AEB ;
reg  AEC ;
reg  AED ;
reg  AEE ;
reg  AEF ;
reg  AEG ;
reg  AEH ;
reg  AEI ;
reg  AEJ ;
reg  AEK ;
reg  AEL ;
reg  AEM ;
reg  AEN ;
reg  AEO ;
reg  AEP ;
reg  AFA ;
reg  AFB ;
reg  AFC ;
reg  AFD ;
reg  AFE ;
reg  AFF ;
reg  AFG ;
reg  AFH ;
reg  AFI ;
reg  AFJ ;
reg  AFK ;
reg  AFL ;
reg  AFM ;
reg  AFN ;
reg  AFO ;
reg  AFP ;
reg  AGA ;
reg  AGB ;
reg  AGC ;
reg  AGD ;
reg  AGE ;
reg  AGF ;
reg  AGG ;
reg  AGH ;
reg  AGI ;
reg  AGJ ;
reg  AGK ;
reg  AGL ;
reg  AGM ;
reg  AGN ;
reg  AGO ;
reg  AGP ;
reg  AHA ;
reg  AHB ;
reg  AHC ;
reg  AHD ;
reg  AHE ;
reg  AHF ;
reg  AHG ;
reg  AHH ;
reg  AHI ;
reg  AHJ ;
reg  AHK ;
reg  AHL ;
reg  AHM ;
reg  AHN ;
reg  AHO ;
reg  AHP ;
reg  aia ;
reg  aib ;
reg  aic ;
reg  aid ;
reg  aie ;
reg  aif ;
reg  aig ;
reg  aih ;
reg  aii ;
reg  aij ;
reg  aik ;
reg  ail ;
reg  aim ;
reg  ain ;
reg  aio ;
reg  aip ;
reg  aja ;
reg  ajb ;
reg  ajc ;
reg  ajd ;
reg  aje ;
reg  ajf ;
reg  ajg ;
reg  ajh ;
reg  aji ;
reg  ajj ;
reg  ajk ;
reg  ajl ;
reg  ajm ;
reg  ajn ;
reg  ajo ;
reg  ajp ;
reg  aka ;
reg  akb ;
reg  akc ;
reg  akd ;
reg  ake ;
reg  akf ;
reg  akg ;
reg  akh ;
reg  aki ;
reg  akj ;
reg  akk ;
reg  akl ;
reg  akm ;
reg  akn ;
reg  ako ;
reg  akp ;
reg  ala ;
reg  alb ;
reg  alc ;
reg  ald ;
reg  ale ;
reg  alf ;
reg  alg ;
reg  alh ;
reg  ali ;
reg  alj ;
reg  alk ;
reg  all ;
reg  alm ;
reg  aln ;
reg  alo ;
reg  alp ;
reg  CAA ;
reg  CAB ;
reg  CAC ;
reg  CAD ;
reg  CAE ;
reg  CAF ;
reg  CAG ;
reg  CAH ;
reg  CAI ;
reg  CAJ ;
reg  CAK ;
reg  CAL ;
reg  CAM ;
reg  CAN ;
reg  CAO ;
reg  CAP ;
reg  CBA ;
reg  CBB ;
reg  CBC ;
reg  CBD ;
reg  CBE ;
reg  CBF ;
reg  CBG ;
reg  CBH ;
reg  CBI ;
reg  CBJ ;
reg  CBK ;
reg  CBL ;
reg  CBM ;
reg  CBN ;
reg  CBO ;
reg  CBP ;
reg  ccb ;
reg  ccc ;
reg  ccd ;
reg  cce ;
reg  ccf ;
reg  ccg ;
reg  cch ;
reg  cci ;
reg  ccj ;
reg  cck ;
reg  ccl ;
reg  ccm ;
reg  ccn ;
reg  cco ;
reg  ccp ;
reg  cda ;
reg  cdb ;
reg  cdc ;
reg  cdd ;
reg  cde ;
reg  cdf ;
reg  cdg ;
reg  cdh ;
reg  cdi ;
reg  cdj ;
reg  cdk ;
reg  cdl ;
reg  cdm ;
reg  cdn ;
reg  cdo ;
reg  cdp ;
reg  CEA ;
reg  CEB ;
reg  CEC ;
reg  CED ;
reg  CEE ;
reg  CEF ;
reg  CEG ;
reg  CEH ;
reg  CEI ;
reg  CEJ ;
reg  CEK ;
reg  CEL ;
reg  CEM ;
reg  CEN ;
reg  CEO ;
reg  CEP ;
reg  CFA ;
reg  CFB ;
reg  CFC ;
reg  CFD ;
reg  CFE ;
reg  CFF ;
reg  CFG ;
reg  CFH ;
reg  CFI ;
reg  CFJ ;
reg  CFK ;
reg  CFL ;
reg  CFM ;
reg  CFN ;
reg  CFO ;
reg  CFP ;
reg  cgb ;
reg  cgc ;
reg  cgd ;
reg  cge ;
reg  cgf ;
reg  cgg ;
reg  cgh ;
reg  cgi ;
reg  cgj ;
reg  cgk ;
reg  cgl ;
reg  cgm ;
reg  cgn ;
reg  cgo ;
reg  cgp ;
reg  cha ;
reg  chb ;
reg  chc ;
reg  chd ;
reg  che ;
reg  chf ;
reg  chg ;
reg  chh ;
reg  chi ;
reg  chj ;
reg  chk ;
reg  chl ;
reg  chm ;
reg  chn ;
reg  cho ;
reg  chp ;
reg  dab ;
reg  dac ;
reg  dad ;
reg  dae ;
reg  daf ;
reg  dag ;
reg  dah ;
reg  dai ;
reg  daj ;
reg  dak ;
reg  dal ;
reg  dam ;
reg  dan ;
reg  dao ;
reg  dap ;
reg  dba ;
reg  dbb ;
reg  dbc ;
reg  dbd ;
reg  dbe ;
reg  dbf ;
reg  dbg ;
reg  dbh ;
reg  dbi ;
reg  dbj ;
reg  dbk ;
reg  dbl ;
reg  dbm ;
reg  dbn ;
reg  dbo ;
reg  dbp ;
reg  EAB ;
reg  EAC ;
reg  EAD ;
reg  EAE ;
reg  EAF ;
reg  EAG ;
reg  EAH ;
reg  EAI ;
reg  EAJ ;
reg  EAK ;
reg  EAL ;
reg  EAM ;
reg  EAN ;
reg  EAO ;
reg  EAP ;
reg  EBB ;
reg  EBC ;
reg  EBD ;
reg  EBE ;
reg  EBF ;
reg  EBG ;
reg  EBH ;
reg  EDA ;
reg  EDB ;
reg  EDC ;
reg  EDD ;
reg  EDE ;
reg  EDF ;
reg  EDG ;
reg  EDH ;
reg  EDI ;
reg  EDJ ;
reg  EDK ;
reg  EDL ;
reg  EDM ;
reg  EDN ;
reg  EDO ;
reg  EDP ;
reg  FAA ;
reg  FAB ;
reg  FAC ;
reg  FAD ;
reg  FAE ;
reg  FAF ;
reg  FAG ;
reg  FAH ;
reg  FAI ;
reg  FAJ ;
reg  FAK ;
reg  FAL ;
reg  FAM ;
reg  FAN ;
reg  FCA ;
reg  FCB ;
reg  FCC ;
reg  FCD ;
reg  FCE ;
reg  FCF ;
reg  FCG ;
reg  FCH ;
reg  FCI ;
reg  FCJ ;
reg  FCK ;
reg  FCL ;
reg  FCM ;
reg  FCN ;
reg  FCO ;
reg  FCP ;
reg  FCQ ;
reg  FCR ;
reg  FCS ;
reg  FCT ;
reg  FCU ;
reg  FCV ;
reg  FDA ;
reg  FDB ;
reg  FDC ;
reg  FDD ;
reg  FDE ;
reg  FDF ;
reg  FDG ;
reg  FDH ;
reg  FDI ;
reg  FDJ ;
reg  FDK ;
reg  FDL ;
reg  FDM ;
reg  FDN ;
reg  FDO ;
reg  FDP ;
reg  FDQ ;
reg  FDR ;
reg  FDS ;
reg  FDT ;
reg  FDU ;
reg  FDV ;
reg  FEA ;
reg  FEB ;
reg  FEC ;
reg  FED ;
reg  FEE ;
reg  FEF ;
reg  FEI ;
reg  FEJ ;
reg  FEK ;
reg  FEL ;
reg  FEM ;
reg  FEN ;
reg  ffb ;
reg  ffc ;
reg  ffd ;
reg  ffe ;
reg  fff ;
reg  ffj ;
reg  ffk ;
reg  ffl ;
reg  ffm ;
reg  HAA ;
reg  HAB ;
reg  HAC ;
reg  HAD ;
reg  HAE ;
reg  HAF ;
reg  HAG ;
reg  HAH ;
reg  HAI ;
reg  HAJ ;
reg  HAK ;
reg  HAL ;
reg  HAM ;
reg  HAN ;
reg  HAO ;
reg  HAP ;
reg  HAQ ;
reg  HAR ;
reg  HAS ;
reg  HAT ;
reg  HAU ;
reg  HAV ;
reg  HAW ;
reg  HAX ;
reg  MAA ;
reg  MAB ;
reg  MAC ;
reg  MAD ;
reg  MBA ;
reg  MBB ;
reg  MBC ;
reg  MBD ;
reg  nab ;
reg  nac ;
reg  nad ;
reg  nbb ;
reg  nbc ;
reg  nbd ;
reg  OAA ;
reg  OAB ;
reg  OAC ;
reg  OAD ;
reg  OAE ;
reg  OAF ;
reg  OAG ;
reg  OAH ;
reg  OAI ;
reg  OAJ ;
reg  OAK ;
reg  OAL ;
reg  OAM ;
reg  OAN ;
reg  OBA ;
reg  OBB ;
reg  OBC ;
reg  OBD ;
reg  OBE ;
reg  OBF ;
reg  OBG ;
reg  OBH ;
reg  OBI ;
reg  OBJ ;
reg  OBK ;
reg  OBL ;
reg  OBM ;
reg  OBN ;
reg  OCA ;
reg  OCB ;
reg  OCC ;
reg  OCD ;
reg  OCE ;
reg  OCF ;
reg  OCG ;
reg  OCH ;
reg  OCI ;
reg  OCJ ;
reg  OCK ;
reg  OCL ;
reg  OCM ;
reg  OCN ;
reg  ODA ;
reg  ODB ;
reg  ODC ;
reg  ODD ;
reg  ODE ;
reg  ODF ;
reg  ODG ;
reg  ODH ;
reg  ODI ;
reg  ODJ ;
reg  ODK ;
reg  ODL ;
reg  ODM ;
reg  ODN ;
reg  OEA ;
reg  OEB ;
reg  OEC ;
reg  OED ;
reg  OEE ;
reg  OEF ;
reg  OEG ;
reg  OEH ;
reg  OEI ;
reg  OEJ ;
reg  OEK ;
reg  OEL ;
reg  OEM ;
reg  OEN ;
reg  OEO ;
reg  OEP ;
reg  OEQ ;
reg  OER ;
reg  OES ;
reg  OET ;
reg  OEU ;
reg  OEV ;
reg  oew ;
reg  oex ;
reg  ofa ;
reg  ofb ;
reg  ofc ;
reg  ofd ;
reg  oha ;
reg  ohb ;
reg  ohc ;
reg  ohd ;
reg  OHE ;
reg  OIA ;
reg  OIB ;
reg  OIC ;
reg  OID ;
reg  OIE ;
reg  OIF ;
reg  OIG ;
reg  OIH ;
reg  OKA ;
reg  OLA ;
reg  OLB ;
reg  OLC ;
reg  OLD ;
reg  paa ;
reg  pab ;
reg  pac ;
reg  pad ;
reg  pae ;
reg  paf ;
reg  pag ;
reg  pah ;
reg  pai ;
reg  paj ;
reg  pak ;
reg  pam ;
reg  pan ;
reg  pao ;
reg  pap ;
reg  paq ;
reg  par ;
reg  pba ;
reg  pbb ;
reg  pbc ;
reg  pbd ;
reg  pbe ;
reg  pbf ;
reg  pbg ;
reg  pbh ;
reg  pbi ;
reg  pbj ;
reg  pbk ;
reg  pbm ;
reg  pbn ;
reg  pbo ;
reg  pbp ;
reg  pbq ;
reg  pbr ;
reg  pca ;
reg  pcb ;
reg  pcc ;
reg  pcd ;
reg  pce ;
reg  pcf ;
reg  pcg ;
reg  pch ;
reg  pci ;
reg  pcj ;
reg  pck ;
reg  pcm ;
reg  pcn ;
reg  pco ;
reg  pcp ;
reg  pcq ;
reg  pcr ;
reg  pda ;
reg  pdb ;
reg  pdc ;
reg  pdd ;
reg  pde ;
reg  pdf ;
reg  pdg ;
reg  pdh ;
reg  pdi ;
reg  pdj ;
reg  pdk ;
reg  pdm ;
reg  pdn ;
reg  pdo ;
reg  pdp ;
reg  pdq ;
reg  pdr ;
reg  pea ;
reg  peb ;
reg  pec ;
reg  ped ;
reg  pee ;
reg  pef ;
reg  peg ;
reg  peh ;
reg  pei ;
reg  pej ;
reg  pek ;
reg  pem ;
reg  pen ;
reg  peo ;
reg  pep ;
reg  peq ;
reg  per ;
reg  pfa ;
reg  pfb ;
reg  pfc ;
reg  pfd ;
reg  pfe ;
reg  pff ;
reg  pfg ;
reg  pfh ;
reg  pfi ;
reg  pfj ;
reg  pfk ;
reg  pfm ;
reg  pfn ;
reg  pfo ;
reg  pfp ;
reg  pfq ;
reg  pfr ;
reg  pga ;
reg  pgb ;
reg  pgc ;
reg  pgd ;
reg  pge ;
reg  pgf ;
reg  pgg ;
reg  pgh ;
reg  pgi ;
reg  pgj ;
reg  pgk ;
reg  pgm ;
reg  pgn ;
reg  pgo ;
reg  pgp ;
reg  pgq ;
reg  pgr ;
reg  pha ;
reg  phb ;
reg  phc ;
reg  phd ;
reg  phe ;
reg  phf ;
reg  phg ;
reg  phh ;
reg  phi ;
reg  phj ;
reg  phk ;
reg  phm ;
reg  phn ;
reg  pho ;
reg  php ;
reg  phq ;
reg  phr ;
reg  pia ;
reg  pib ;
reg  pic ;
reg  pid ;
reg  pie ;
reg  pif ;
reg  pig ;
reg  pih ;
reg  pii ;
reg  pij ;
reg  pik ;
reg  pim ;
reg  pin ;
reg  pio ;
reg  pip ;
reg  piq ;
reg  pir ;
reg  pja ;
reg  pjb ;
reg  pjc ;
reg  pjd ;
reg  pje ;
reg  pjf ;
reg  pjg ;
reg  pjh ;
reg  pji ;
reg  pjj ;
reg  pjk ;
reg  pjm ;
reg  pjn ;
reg  pjo ;
reg  pjp ;
reg  pjq ;
reg  pjr ;
reg  qaa ;
reg  qab ;
reg  QAC ;
reg  QBA ;
reg  QBB ;
reg  QBC ;
reg  QBD ;
reg  QBE ;
reg  QBF ;
reg  QBG ;
reg  QBH ;
reg  QCA ;
reg  QCB ;
reg  QCC ;
reg  QCD ;
reg  qda ;
reg  qdb ;
reg  qdc ;
reg  qdd ;
reg  qde ;
reg  qdf ;
reg  qdg ;
reg  qdh ;
reg  QEA ;
reg  QEB ;
reg  QEC ;
reg  QFA ;
reg  QFB ;
reg  QFC ;
reg  QFD ;
reg  QGA ;
reg  QGB ;
reg  QGC ;
reg  QGD ;
reg  QMA ;
reg  QMB ;
reg  QMC ;
reg  QMD ;
reg  QME ;
reg  QMF ;
reg  QMG ;
reg  QMH ;
reg  QNA ;
reg  QNB ;
reg  QNC ;
reg  QND ;
reg  QNE ;
reg  QNF ;
reg  QNG ;
reg  QNH ;
reg  QNI ;
reg  QNJ ;
reg  QRA ;
reg  QRB ;
reg  qta ;
reg  qtb ;
reg  qtc ;
reg  qtd ;
reg  saa ;
reg  sab ;
reg  sac ;
reg  sad ;
reg  sae ;
reg  saf ;
reg  sag ;
reg  sah ;
reg  sai ;
reg  saj ;
reg  sak ;
reg  sal ;
reg  sam ;
reg  san ;
reg  sao ;
reg  sap ;
reg  saq ;
reg  sar ;
reg  sas ;
reg  sat ;
reg  sau ;
reg  sav ;
reg  saw ;
reg  sax ;
reg  sba ;
reg  sbb ;
reg  sbc ;
reg  sbd ;
reg  sbe ;
reg  sbf ;
reg  sbg ;
reg  sbh ;
reg  sbi ;
reg  sbj ;
reg  sbk ;
reg  sbl ;
reg  sbm ;
reg  sbn ;
reg  sbo ;
reg  sbp ;
reg  sbq ;
reg  sbr ;
reg  sbs ;
reg  sbt ;
reg  sbu ;
reg  sbv ;
reg  sbw ;
reg  sbx ;
reg  sca ;
reg  scb ;
reg  scc ;
reg  scd ;
reg  sce ;
reg  scf ;
reg  scg ;
reg  sch ;
reg  sci ;
reg  scj ;
reg  sck ;
reg  scl ;
reg  scm ;
reg  scn ;
reg  sco ;
reg  scp ;
reg  scq ;
reg  scr ;
reg  scs ;
reg  sct ;
reg  scu ;
reg  scv ;
reg  scw ;
reg  scx ;
reg  sda ;
reg  sdb ;
reg  sdc ;
reg  sdd ;
reg  sde ;
reg  sdf ;
reg  sdg ;
reg  sdh ;
reg  sdi ;
reg  sdj ;
reg  sdk ;
reg  sdl ;
reg  sdm ;
reg  sdn ;
reg  sdo ;
reg  sdp ;
reg  sdq ;
reg  sdr ;
reg  sds ;
reg  sdt ;
reg  sdu ;
reg  sdv ;
reg  sdw ;
reg  sdx ;
reg  sea ;
reg  seb ;
reg  sec ;
reg  sed ;
reg  see ;
reg  sef ;
reg  seg ;
reg  seh ;
reg  sei ;
reg  sej ;
reg  sek ;
reg  sel ;
reg  sem ;
reg  sen ;
reg  seo ;
reg  sep ;
reg  seq ;
reg  ser ;
reg  ses ;
reg  set ;
reg  seu ;
reg  sev ;
reg  sew ;
reg  sex ;
reg  sfa ;
reg  sfb ;
reg  sfc ;
reg  sfd ;
reg  sfe ;
reg  sff ;
reg  sfg ;
reg  sfh ;
reg  sfi ;
reg  sfj ;
reg  sfk ;
reg  sfl ;
reg  sfm ;
reg  sfn ;
reg  sfo ;
reg  sfp ;
reg  sfq ;
reg  sfr ;
reg  sfs ;
reg  sft ;
reg  sfu ;
reg  sfv ;
reg  sfw ;
reg  sfx ;
reg  sga ;
reg  sgb ;
reg  sgc ;
reg  sgd ;
reg  sge ;
reg  sgf ;
reg  sgg ;
reg  sgh ;
reg  sgi ;
reg  sgj ;
reg  sgk ;
reg  sgl ;
reg  sgm ;
reg  sgn ;
reg  sgo ;
reg  sgp ;
reg  sgq ;
reg  sgr ;
reg  sgs ;
reg  sgt ;
reg  sgu ;
reg  sgv ;
reg  sgw ;
reg  sgx ;
reg  sha ;
reg  shb ;
reg  shc ;
reg  shd ;
reg  she ;
reg  shf ;
reg  shg ;
reg  shh ;
reg  shi ;
reg  shj ;
reg  shk ;
reg  shl ;
reg  shm ;
reg  shn ;
reg  sho ;
reg  shp ;
reg  shq ;
reg  shr ;
reg  shs ;
reg  sht ;
reg  shu ;
reg  shv ;
reg  shw ;
reg  shx ;
reg  sia ;
reg  sib ;
reg  sic ;
reg  sid ;
reg  sie ;
reg  sif ;
reg  sig ;
reg  sih ;
reg  sii ;
reg  sij ;
reg  sik ;
reg  sil ;
reg  sim ;
reg  sin ;
reg  sio ;
reg  sip ;
reg  siq ;
reg  sir ;
reg  sis ;
reg  sit ;
reg  siu ;
reg  siv ;
reg  siw ;
reg  six ;
reg  sja ;
reg  sjb ;
reg  sjc ;
reg  sjd ;
reg  sje ;
reg  sjf ;
reg  sjg ;
reg  sjh ;
reg  sji ;
reg  sjj ;
reg  sjk ;
reg  sjl ;
reg  sjm ;
reg  sjn ;
reg  sjo ;
reg  sjp ;
reg  sjq ;
reg  sjr ;
reg  sjs ;
reg  sjt ;
reg  sju ;
reg  sjv ;
reg  sjw ;
reg  sjx ;
reg  TAA ;
reg  TAB ;
reg  TAC ;
reg  TAD ;
reg  TAE ;
reg  TAF ;
reg  TAG ;
reg  TBA ;
reg  TBB ;
reg  TBC ;
reg  TBD ;
reg  TBE ;
reg  TBF ;
reg  TCA ;
reg  TCB ;
reg  TCC ;
reg  TCD ;
reg  TCE ;
reg  TCF ;
reg  TCG ;
reg  TDA ;
reg  TDB ;
reg  TDC ;
reg  TDD ;
reg  TDE ;
reg  TDF ;
reg  TEA ;
reg  TEB ;
reg  TFA ;
reg  TFB ;
reg  TGA ;
reg  TGB ;
reg  tha ;
reg  thb ;
reg  thc ;
reg  thd ;
reg  TIC ;
reg  TID ;
reg  TJC ;
reg  TJD ;
reg  TKC ;
reg  TKD ;
reg  TLC ;
reg  TLD ;
reg  TMA ;
reg  TMB ;
reg  TMC ;
reg  TMD ;
reg  TNA ;
reg  TNB ;
reg  TNC ;
reg  TND ;
reg  WAA ;
reg  WAB ;
reg  WAC ;
reg  WAD ;
reg  WAE ;
reg  WAF ;
reg  WAG ;
reg  WAH ;
reg  WAI ;
reg  WAJ ;
reg  WAK ;
reg  WAL ;
reg  WAM ;
reg  WAN ;
reg  WBA ;
reg  WBB ;
reg  WBC ;
reg  WBD ;
reg  WBE ;
reg  WBF ;
reg  WBG ;
reg  WBH ;
reg  WBI ;
reg  WBJ ;
reg  WBK ;
reg  WBL ;
reg  WBM ;
reg  WBN ;
reg  WCA ;
reg  WCB ;
reg  WCC ;
reg  WCD ;
reg  WCE ;
reg  WCF ;
reg  WCG ;
reg  WCH ;
reg  WCI ;
reg  WCJ ;
reg  WCK ;
reg  WCL ;
reg  WCM ;
reg  WCN ;
reg  WDA ;
reg  WDB ;
reg  WDC ;
reg  WDD ;
reg  WDE ;
reg  WDF ;
reg  WDG ;
reg  WDH ;
reg  WDI ;
reg  WDJ ;
reg  WDK ;
reg  WDL ;
reg  WDM ;
reg  WDN ;
wire  aaa ;
wire  aab ;
wire  aac ;
wire  aad ;
wire  aae ;
wire  aaf ;
wire  aag ;
wire  aah ;
wire  aai ;
wire  aaj ;
wire  aak ;
wire  aal ;
wire  aam ;
wire  aan ;
wire  aao ;
wire  aap ;
wire  aba ;
wire  abb ;
wire  abc ;
wire  abd ;
wire  abe ;
wire  abf ;
wire  abg ;
wire  abh ;
wire  abi ;
wire  abj ;
wire  abk ;
wire  abl ;
wire  abm ;
wire  abn ;
wire  abo ;
wire  abp ;
wire  aca ;
wire  acb ;
wire  acc ;
wire  acd ;
wire  ace ;
wire  acf ;
wire  acg ;
wire  ach ;
wire  aci ;
wire  acj ;
wire  ack ;
wire  acl ;
wire  acm ;
wire  acn ;
wire  aco ;
wire  acp ;
wire  ada ;
wire  adb ;
wire  adc ;
wire  add ;
wire  ade ;
wire  adf ;
wire  adg ;
wire  adh ;
wire  adi ;
wire  adj ;
wire  adk ;
wire  adl ;
wire  adm ;
wire  adn ;
wire  ado ;
wire  adp ;
wire  aea ;
wire  aeb ;
wire  aec ;
wire  aed ;
wire  aee ;
wire  aef ;
wire  aeg ;
wire  aeh ;
wire  aei ;
wire  aej ;
wire  aek ;
wire  ael ;
wire  aem ;
wire  aen ;
wire  aeo ;
wire  aep ;
wire  afa ;
wire  afb ;
wire  afc ;
wire  afd ;
wire  afe ;
wire  aff ;
wire  afg ;
wire  afh ;
wire  afi ;
wire  afj ;
wire  afk ;
wire  afl ;
wire  afm ;
wire  afn ;
wire  afo ;
wire  afp ;
wire  aga ;
wire  agb ;
wire  agc ;
wire  agd ;
wire  age ;
wire  agf ;
wire  agg ;
wire  agh ;
wire  agi ;
wire  agj ;
wire  agk ;
wire  agl ;
wire  agm ;
wire  agn ;
wire  ago ;
wire  agp ;
wire  aha ;
wire  ahb ;
wire  ahc ;
wire  ahd ;
wire  ahe ;
wire  ahf ;
wire  ahg ;
wire  ahh ;
wire  ahi ;
wire  ahj ;
wire  ahk ;
wire  ahl ;
wire  ahm ;
wire  ahn ;
wire  aho ;
wire  ahp ;
wire  AIA ;
wire  AIB ;
wire  AIC ;
wire  AID ;
wire  AIE ;
wire  AIF ;
wire  AIG ;
wire  AIH ;
wire  AII ;
wire  AIJ ;
wire  AIK ;
wire  AIL ;
wire  AIM ;
wire  AIN ;
wire  AIO ;
wire  AIP ;
wire  AJA ;
wire  AJB ;
wire  AJC ;
wire  AJD ;
wire  AJE ;
wire  AJF ;
wire  AJG ;
wire  AJH ;
wire  AJI ;
wire  AJJ ;
wire  AJK ;
wire  AJL ;
wire  AJM ;
wire  AJN ;
wire  AJO ;
wire  AJP ;
wire  AKA ;
wire  AKB ;
wire  AKC ;
wire  AKD ;
wire  AKE ;
wire  AKF ;
wire  AKG ;
wire  AKH ;
wire  AKI ;
wire  AKJ ;
wire  AKK ;
wire  AKL ;
wire  AKM ;
wire  AKN ;
wire  AKO ;
wire  AKP ;
wire  ALA ;
wire  ALB ;
wire  ALC ;
wire  ALD ;
wire  ALE ;
wire  ALF ;
wire  ALG ;
wire  ALH ;
wire  ALI ;
wire  ALJ ;
wire  ALK ;
wire  ALL ;
wire  ALM ;
wire  ALN ;
wire  ALO ;
wire  ALP ;
wire  baa ;
wire  BAA ;
wire  bab ;
wire  BAB ;
wire  bac ;
wire  BAC ;
wire  bad ;
wire  BAD ;
wire  bae ;
wire  BAE ;
wire  baf ;
wire  BAF ;
wire  bag ;
wire  BAG ;
wire  bah ;
wire  BAH ;
wire  bai ;
wire  BAI ;
wire  baj ;
wire  BAJ ;
wire  bak ;
wire  BAK ;
wire  bal ;
wire  BAL ;
wire  bam ;
wire  BAM ;
wire  ban ;
wire  BAN ;
wire  bao ;
wire  BAO ;
wire  bap ;
wire  BAP ;
wire  bba ;
wire  BBA ;
wire  bbb ;
wire  BBB ;
wire  bbc ;
wire  BBC ;
wire  bbd ;
wire  BBD ;
wire  bbe ;
wire  BBE ;
wire  bbf ;
wire  BBF ;
wire  bbg ;
wire  BBG ;
wire  bbh ;
wire  BBH ;
wire  bbi ;
wire  BBI ;
wire  bbj ;
wire  BBJ ;
wire  bbk ;
wire  BBK ;
wire  bbl ;
wire  BBL ;
wire  bbm ;
wire  BBM ;
wire  bbn ;
wire  BBN ;
wire  bbo ;
wire  BBO ;
wire  bbp ;
wire  BBP ;
wire  bcb ;
wire  BCB ;
wire  bcc ;
wire  BCC ;
wire  bcd ;
wire  BCD ;
wire  bce ;
wire  BCE ;
wire  bcf ;
wire  BCF ;
wire  bcg ;
wire  BCG ;
wire  bch ;
wire  BCH ;
wire  bci ;
wire  BCI ;
wire  bcj ;
wire  BCJ ;
wire  bck ;
wire  BCK ;
wire  bcl ;
wire  BCL ;
wire  bcm ;
wire  BCM ;
wire  bcn ;
wire  BCN ;
wire  bco ;
wire  BCO ;
wire  bcp ;
wire  BCP ;
wire  bda ;
wire  BDA ;
wire  bdb ;
wire  BDB ;
wire  bdc ;
wire  BDC ;
wire  bdd ;
wire  BDD ;
wire  bde ;
wire  BDE ;
wire  bdf ;
wire  BDF ;
wire  bdg ;
wire  BDG ;
wire  bdh ;
wire  BDH ;
wire  bdi ;
wire  BDI ;
wire  bdj ;
wire  BDJ ;
wire  bdk ;
wire  BDK ;
wire  bdl ;
wire  BDL ;
wire  bdm ;
wire  BDM ;
wire  bdn ;
wire  BDN ;
wire  bdo ;
wire  BDO ;
wire  bdp ;
wire  BDP ;
wire  bee ;
wire  BEE ;
wire  bei ;
wire  BEI ;
wire  bem ;
wire  BEM ;
wire  bfa ;
wire  BFA ;
wire  bfe ;
wire  BFE ;
wire  bfi ;
wire  BFI ;
wire  bfm ;
wire  BFM ;
wire  caa ;
wire  cab ;
wire  cac ;
wire  cad ;
wire  cae ;
wire  caf ;
wire  cag ;
wire  cah ;
wire  cai ;
wire  caj ;
wire  cak ;
wire  cal ;
wire  cam ;
wire  can ;
wire  cao ;
wire  cap ;
wire  cba ;
wire  cbb ;
wire  cbc ;
wire  cbd ;
wire  cbe ;
wire  cbf ;
wire  cbg ;
wire  cbh ;
wire  cbi ;
wire  cbj ;
wire  cbk ;
wire  cbl ;
wire  cbm ;
wire  cbn ;
wire  cbo ;
wire  cbp ;
wire  CCB ;
wire  CCC ;
wire  CCD ;
wire  CCE ;
wire  CCF ;
wire  CCG ;
wire  CCH ;
wire  CCI ;
wire  CCJ ;
wire  CCK ;
wire  CCL ;
wire  CCM ;
wire  CCN ;
wire  CCO ;
wire  CCP ;
wire  CDA ;
wire  CDB ;
wire  CDC ;
wire  CDD ;
wire  CDE ;
wire  CDF ;
wire  CDG ;
wire  CDH ;
wire  CDI ;
wire  CDJ ;
wire  CDK ;
wire  CDL ;
wire  CDM ;
wire  CDN ;
wire  CDO ;
wire  CDP ;
wire  cea ;
wire  ceb ;
wire  cec ;
wire  ced ;
wire  cee ;
wire  cef ;
wire  ceg ;
wire  ceh ;
wire  cei ;
wire  cej ;
wire  cek ;
wire  cel ;
wire  cem ;
wire  cen ;
wire  ceo ;
wire  cep ;
wire  cfa ;
wire  cfb ;
wire  cfc ;
wire  cfd ;
wire  cfe ;
wire  cff ;
wire  cfg ;
wire  cfh ;
wire  cfi ;
wire  cfj ;
wire  cfk ;
wire  cfl ;
wire  cfm ;
wire  cfn ;
wire  cfo ;
wire  cfp ;
wire  CGB ;
wire  CGC ;
wire  CGD ;
wire  CGE ;
wire  CGF ;
wire  CGG ;
wire  CGH ;
wire  CGI ;
wire  CGJ ;
wire  CGK ;
wire  CGL ;
wire  CGM ;
wire  CGN ;
wire  CGO ;
wire  CGP ;
wire  CHA ;
wire  CHB ;
wire  CHC ;
wire  CHD ;
wire  CHE ;
wire  CHF ;
wire  CHG ;
wire  CHH ;
wire  CHI ;
wire  CHJ ;
wire  CHK ;
wire  CHL ;
wire  CHM ;
wire  CHN ;
wire  CHO ;
wire  CHP ;
wire  DAB ;
wire  DAC ;
wire  DAD ;
wire  DAE ;
wire  DAF ;
wire  DAG ;
wire  DAH ;
wire  DAI ;
wire  DAJ ;
wire  DAK ;
wire  DAL ;
wire  DAM ;
wire  DAN ;
wire  DAO ;
wire  DAP ;
wire  DBA ;
wire  DBB ;
wire  DBC ;
wire  DBD ;
wire  DBE ;
wire  DBF ;
wire  DBG ;
wire  DBH ;
wire  DBI ;
wire  DBJ ;
wire  DBK ;
wire  DBL ;
wire  DBM ;
wire  DBN ;
wire  DBO ;
wire  DBP ;
wire  eab ;
wire  eac ;
wire  ead ;
wire  eae ;
wire  eaf ;
wire  eag ;
wire  eah ;
wire  eai ;
wire  eaj ;
wire  eak ;
wire  eal ;
wire  eam ;
wire  ean ;
wire  eao ;
wire  eap ;
wire  ebb ;
wire  ebc ;
wire  ebd ;
wire  ebe ;
wire  ebf ;
wire  ebg ;
wire  ebh ;
wire  eda ;
wire  edb ;
wire  edc ;
wire  edd ;
wire  ede ;
wire  edf ;
wire  edg ;
wire  edh ;
wire  edi ;
wire  edj ;
wire  edk ;
wire  edl ;
wire  edm ;
wire  edn ;
wire  edo ;
wire  edp ;
wire  faa ;
wire  fab ;
wire  fac ;
wire  fad ;
wire  fae ;
wire  faf ;
wire  fag ;
wire  fah ;
wire  fai ;
wire  faj ;
wire  fak ;
wire  fal ;
wire  fam ;
wire  fan ;
wire  fca ;
wire  fcb ;
wire  fcc ;
wire  fcd ;
wire  fce ;
wire  fcf ;
wire  fcg ;
wire  fch ;
wire  fci ;
wire  fcj ;
wire  fck ;
wire  fcl ;
wire  fcm ;
wire  fcn ;
wire  fco ;
wire  fcp ;
wire  fcq ;
wire  fcr ;
wire  fcs ;
wire  fct ;
wire  fcu ;
wire  fcv ;
wire  fda ;
wire  fdb ;
wire  fdc ;
wire  fdd ;
wire  fde ;
wire  fdf ;
wire  fdg ;
wire  fdh ;
wire  fdi ;
wire  fdj ;
wire  fdk ;
wire  fdl ;
wire  fdm ;
wire  fdn ;
wire  fdo ;
wire  fdp ;
wire  fdq ;
wire  fdr ;
wire  fds ;
wire  fdt ;
wire  fdu ;
wire  fdv ;
wire  fea ;
wire  feb ;
wire  fec ;
wire  fed ;
wire  fee ;
wire  fef ;
wire  fei ;
wire  fej ;
wire  fek ;
wire  fel ;
wire  fem ;
wire  fen ;
wire  FFB ;
wire  FFC ;
wire  FFD ;
wire  FFE ;
wire  FFF ;
wire  FFJ ;
wire  FFK ;
wire  FFL ;
wire  FFM ;
wire  gaa ;
wire  GAA ;
wire  gab ;
wire  GAB ;
wire  gac ;
wire  GAC ;
wire  gad ;
wire  GAD ;
wire  gae ;
wire  GAE ;
wire  gaf ;
wire  GAF ;
wire  haa ;
wire  hab ;
wire  hac ;
wire  had ;
wire  hae ;
wire  haf ;
wire  hag ;
wire  hah ;
wire  hai ;
wire  haj ;
wire  hak ;
wire  hal ;
wire  ham ;
wire  han ;
wire  hao ;
wire  hap ;
wire  haq ;
wire  har ;
wire  has ;
wire  hat ;
wire  hau ;
wire  hav ;
wire  haw ;
wire  hax ;
wire  iaa ;
wire  iab ;
wire  iac ;
wire  iad ;
wire  iae ;
wire  iaf ;
wire  iag ;
wire  iah ;
wire  iai ;
wire  iaj ;
wire  iak ;
wire  ial ;
wire  iam ;
wire  ian ;
wire  iao ;
wire  iap ;
wire  iba ;
wire  ibb ;
wire  ibc ;
wire  ibd ;
wire  ibe ;
wire  ibf ;
wire  ibg ;
wire  ibh ;
wire  ibi ;
wire  ibj ;
wire  ibk ;
wire  ibl ;
wire  ibm ;
wire  ibn ;
wire  ibo ;
wire  ibp ;
wire  ica ;
wire  icb ;
wire  icc ;
wire  icd ;
wire  ice ;
wire  icf ;
wire  icg ;
wire  ich ;
wire  ici ;
wire  icj ;
wire  ick ;
wire  icl ;
wire  icm ;
wire  icn ;
wire  ico ;
wire  icp ;
wire  ida ;
wire  idb ;
wire  idc ;
wire  idd ;
wire  ide ;
wire  idf ;
wire  idg ;
wire  idh ;
wire  idi ;
wire  idj ;
wire  idk ;
wire  idl ;
wire  idm ;
wire  idn ;
wire  ido ;
wire  idp ;
wire  iea ;
wire  ieb ;
wire  iec ;
wire  ied ;
wire  iee ;
wire  ief ;
wire  ieg ;
wire  ieh ;
wire  iei ;
wire  iej ;
wire  iek ;
wire  iel ;
wire  iem ;
wire  ien ;
wire  ieo ;
wire  iep ;
wire  ifa ;
wire  ifb ;
wire  ifc ;
wire  ifd ;
wire  ife ;
wire  ifff  ;
wire  ifg ;
wire  ifh ;
wire  ifi ;
wire  ifj ;
wire  ifk ;
wire  ifl ;
wire  ifm ;
wire  ifn ;
wire  ifo ;
wire  ifp ;
wire  iga ;
wire  igb ;
wire  igc ;
wire  igd ;
wire  ige ;
wire  igf ;
wire  igg ;
wire  igh ;
wire  igi ;
wire  igj ;
wire  igk ;
wire  igl ;
wire  igm ;
wire  ign ;
wire  igo ;
wire  igp ;
wire  iha ;
wire  ihb ;
wire  ihc ;
wire  ihd ;
wire  ihe ;
wire  ihf ;
wire  ihg ;
wire  ihh ;
wire  ihi ;
wire  ihj ;
wire  ihk ;
wire  ihl ;
wire  ihm ;
wire  ihn ;
wire  iho ;
wire  ihp ;
wire  iia ;
wire  iib ;
wire  iic ;
wire  iid ;
wire  iie ;
wire  iif ;
wire  ija ;
wire  ijb ;
wire  ijc ;
wire  ijd ;
wire  ije ;
wire  ijf ;
wire  ijg ;
wire  ijh ;
wire  ika ;
wire  ikb ;
wire  ikc ;
wire  ikd ;
wire  ike ;
wire  ikf ;
wire  ikg ;
wire  ikh ;
wire  iki ;
wire  ikj ;
wire  ikk ;
wire  ikm ;
wire  ikn ;
wire  iko ;
wire  ikp ;
wire  ikq ;
wire  ikr ;
wire  iks ;
wire  ikt ;
wire  iku ;
wire  ila ;
wire  jac ;
wire  JAC ;
wire  jad ;
wire  JAD ;
wire  jae ;
wire  JAE ;
wire  jaf ;
wire  JAF ;
wire  jag ;
wire  JAG ;
wire  jdb ;
wire  JDB ;
wire  jdc ;
wire  JDC ;
wire  jdd ;
wire  JDD ;
wire  jdf ;
wire  JDF ;
wire  jdg ;
wire  JDG ;
wire  jdh ;
wire  JDH ;
wire  jdj ;
wire  JDJ ;
wire  jdk ;
wire  JDK ;
wire  jdl ;
wire  JDL ;
wire  jdn ;
wire  JDN ;
wire  jdo ;
wire  JDO ;
wire  jdp ;
wire  JDP ;
wire  jdr ;
wire  JDR ;
wire  jds ;
wire  JDS ;
wire  jdt ;
wire  JDT ;
wire  jdv ;
wire  JDV ;
wire  jeb ;
wire  JEB ;
wire  jec ;
wire  JEC ;
wire  jed ;
wire  JED ;
wire  jef ;
wire  JEF ;
wire  jeg ;
wire  JEG ;
wire  jeh ;
wire  JEH ;
wire  jej ;
wire  JEJ ;
wire  jek ;
wire  JEK ;
wire  jel ;
wire  JEL ;
wire  jen ;
wire  JEN ;
wire  jeo ;
wire  JEO ;
wire  jep ;
wire  JEP ;
wire  jer ;
wire  JER ;
wire  jes ;
wire  JES ;
wire  jet ;
wire  JET ;
wire  jev ;
wire  JEV ;
wire  jfa ;
wire  JFA ;
wire  jfb ;
wire  JFB ;
wire  kaa ;
wire  KAA ;
wire  kab ;
wire  KAB ;
wire  kba ;
wire  KBA ;
wire  kbb ;
wire  KBB ;
wire  kbc ;
wire  KBC ;
wire  kbd ;
wire  KBD ;
wire  kbe ;
wire  KBE ;
wire  kbf ;
wire  KBF ;
wire  kbg ;
wire  KBG ;
wire  kbh ;
wire  KBH ;
wire  kca ;
wire  KCA ;
wire  kcb ;
wire  KCB ;
wire  kcc ;
wire  KCC ;
wire  kcd ;
wire  KCD ;
wire  laa ;
wire  LAA ;
wire  lab ;
wire  LAB ;
wire  lac ;
wire  LAC ;
wire  lad ;
wire  LAD ;
wire  lae ;
wire  LAE ;
wire  laf ;
wire  LAF ;
wire  lag ;
wire  LAG ;
wire  lah ;
wire  LAH ;
wire  lai ;
wire  LAI ;
wire  laj ;
wire  LAJ ;
wire  lak ;
wire  LAK ;
wire  lal ;
wire  LAL ;
wire  lam ;
wire  LAM ;
wire  lan ;
wire  LAN ;
wire  lao ;
wire  LAO ;
wire  lap ;
wire  LAP ;
wire  lbb ;
wire  LBB ;
wire  lbc ;
wire  LBC ;
wire  lbd ;
wire  LBD ;
wire  lbe ;
wire  LBE ;
wire  lbf ;
wire  LBF ;
wire  lbg ;
wire  LBG ;
wire  lbh ;
wire  LBH ;
wire  lbi ;
wire  LBI ;
wire  lbj ;
wire  LBJ ;
wire  lbk ;
wire  LBK ;
wire  lbl ;
wire  LBL ;
wire  lbm ;
wire  LBM ;
wire  lbn ;
wire  LBN ;
wire  lbo ;
wire  LBO ;
wire  lbp ;
wire  LBP ;
wire  lca ;
wire  LCA ;
wire  lcb ;
wire  LCB ;
wire  lcc ;
wire  LCC ;
wire  lcd ;
wire  LCD ;
wire  lce ;
wire  LCE ;
wire  lcf ;
wire  LCF ;
wire  lcg ;
wire  LCG ;
wire  lch ;
wire  LCH ;
wire  lci ;
wire  LCI ;
wire  lcj ;
wire  LCJ ;
wire  lck ;
wire  LCK ;
wire  lcl ;
wire  LCL ;
wire  lcm ;
wire  LCM ;
wire  lcn ;
wire  LCN ;
wire  lco ;
wire  LCO ;
wire  lcp ;
wire  LCP ;
wire  ldb ;
wire  LDB ;
wire  ldc ;
wire  LDC ;
wire  ldd ;
wire  LDD ;
wire  lde ;
wire  LDE ;
wire  ldf ;
wire  LDF ;
wire  ldg ;
wire  LDG ;
wire  ldh ;
wire  LDH ;
wire  ldi ;
wire  LDI ;
wire  ldj ;
wire  LDJ ;
wire  ldk ;
wire  LDK ;
wire  ldl ;
wire  LDL ;
wire  ldm ;
wire  LDM ;
wire  ldn ;
wire  LDN ;
wire  ldo ;
wire  LDO ;
wire  ldp ;
wire  LDP ;
wire  maa ;
wire  mab ;
wire  mac ;
wire  mad ;
wire  mba ;
wire  mbb ;
wire  mbc ;
wire  mbd ;
wire  NAB ;
wire  NAC ;
wire  NAD ;
wire  NBB ;
wire  NBC ;
wire  NBD ;
wire  oaa ;
wire  oab ;
wire  oac ;
wire  oad ;
wire  oae ;
wire  oaf ;
wire  oag ;
wire  oah ;
wire  oai ;
wire  oaj ;
wire  oak ;
wire  oal ;
wire  oam ;
wire  oan ;
wire  oba ;
wire  obb ;
wire  obc ;
wire  obd ;
wire  obe ;
wire  obf ;
wire  obg ;
wire  obh ;
wire  obi ;
wire  obj ;
wire  obk ;
wire  obl ;
wire  obm ;
wire  obn ;
wire  oca ;
wire  ocb ;
wire  occ ;
wire  ocd ;
wire  oce ;
wire  ocf ;
wire  ocg ;
wire  och ;
wire  oci ;
wire  ocj ;
wire  ock ;
wire  ocl ;
wire  ocm ;
wire  ocn ;
wire  oda ;
wire  odb ;
wire  odc ;
wire  odd ;
wire  ode ;
wire  odf ;
wire  odg ;
wire  odh ;
wire  odi ;
wire  odj ;
wire  odk ;
wire  odl ;
wire  odm ;
wire  odn ;
wire  oea ;
wire  oeb ;
wire  oec ;
wire  oed ;
wire  oee ;
wire  oef ;
wire  oeg ;
wire  oeh ;
wire  oei ;
wire  oej ;
wire  oek ;
wire  oel ;
wire  oem ;
wire  oen ;
wire  oeo ;
wire  oep ;
wire  oeq ;
wire  oer ;
wire  oes ;
wire  oet ;
wire  oeu ;
wire  oev ;
wire  OEW ;
wire  OEX ;
wire  OFA ;
wire  OFB ;
wire  OFC ;
wire  OFD ;
wire  OHA ;
wire  OHB ;
wire  OHC ;
wire  OHD ;
wire  ohe ;
wire  oia ;
wire  oib ;
wire  oic ;
wire  oid ;
wire  oie ;
wire  oif ;
wire  oig ;
wire  oih ;
wire  oka ;
wire  ola ;
wire  olb ;
wire  olc ;
wire  old ;
wire  PAA ;
wire  PAB ;
wire  PAC ;
wire  PAD ;
wire  PAE ;
wire  PAF ;
wire  PAG ;
wire  PAH ;
wire  PAI ;
wire  PAJ ;
wire  PAK ;
wire  PAM ;
wire  PAN ;
wire  PAO ;
wire  PAP ;
wire  PAQ ;
wire  PAR ;
wire  PBA ;
wire  PBB ;
wire  PBC ;
wire  PBD ;
wire  PBE ;
wire  PBF ;
wire  PBG ;
wire  PBH ;
wire  PBI ;
wire  PBJ ;
wire  PBK ;
wire  PBM ;
wire  PBN ;
wire  PBO ;
wire  PBP ;
wire  PBQ ;
wire  PBR ;
wire  PCA ;
wire  PCB ;
wire  PCC ;
wire  PCD ;
wire  PCE ;
wire  PCF ;
wire  PCG ;
wire  PCH ;
wire  PCI ;
wire  PCJ ;
wire  PCK ;
wire  PCM ;
wire  PCN ;
wire  PCO ;
wire  PCP ;
wire  PCQ ;
wire  PCR ;
wire  PDA ;
wire  PDB ;
wire  PDC ;
wire  PDD ;
wire  PDE ;
wire  PDF ;
wire  PDG ;
wire  PDH ;
wire  PDI ;
wire  PDJ ;
wire  PDK ;
wire  PDM ;
wire  PDN ;
wire  PDO ;
wire  PDP ;
wire  PDQ ;
wire  PDR ;
wire  PEA ;
wire  PEB ;
wire  PEC ;
wire  PED ;
wire  PEE ;
wire  PEF ;
wire  PEG ;
wire  PEH ;
wire  PEI ;
wire  PEJ ;
wire  PEK ;
wire  PEM ;
wire  PEN ;
wire  PEO ;
wire  PEP ;
wire  PEQ ;
wire  PER ;
wire  PFA ;
wire  PFB ;
wire  PFC ;
wire  PFD ;
wire  PFE ;
wire  PFF ;
wire  PFG ;
wire  PFH ;
wire  PFI ;
wire  PFJ ;
wire  PFK ;
wire  PFM ;
wire  PFN ;
wire  PFO ;
wire  PFP ;
wire  PFQ ;
wire  PFR ;
wire  PGA ;
wire  PGB ;
wire  PGC ;
wire  PGD ;
wire  PGE ;
wire  PGF ;
wire  PGG ;
wire  PGH ;
wire  PGI ;
wire  PGJ ;
wire  PGK ;
wire  PGM ;
wire  PGN ;
wire  PGO ;
wire  PGP ;
wire  PGQ ;
wire  PGR ;
wire  PHA ;
wire  PHB ;
wire  PHC ;
wire  PHD ;
wire  PHE ;
wire  PHF ;
wire  PHG ;
wire  PHH ;
wire  PHI ;
wire  PHJ ;
wire  PHK ;
wire  PHM ;
wire  PHN ;
wire  PHO ;
wire  PHP ;
wire  PHQ ;
wire  PHR ;
wire  PIA ;
wire  PIB ;
wire  PIC ;
wire  PID ;
wire  PIE ;
wire  PIF ;
wire  PIG ;
wire  PIH ;
wire  PII ;
wire  PIJ ;
wire  PIK ;
wire  PIM ;
wire  PIN ;
wire  PIO ;
wire  PIP ;
wire  PIQ ;
wire  PIR ;
wire  PJA ;
wire  PJB ;
wire  PJC ;
wire  PJD ;
wire  PJE ;
wire  PJF ;
wire  PJG ;
wire  PJH ;
wire  PJI ;
wire  PJJ ;
wire  PJK ;
wire  PJM ;
wire  PJN ;
wire  PJO ;
wire  PJP ;
wire  PJQ ;
wire  PJR ;
wire  QAA ;
wire  QAB ;
wire  qac ;
wire  qba ;
wire  qbb ;
wire  qbc ;
wire  qbd ;
wire  qbe ;
wire  qbf ;
wire  qbg ;
wire  qbh ;
wire  qca ;
wire  qcb ;
wire  qcc ;
wire  qcd ;
wire  QDA ;
wire  QDB ;
wire  QDC ;
wire  QDD ;
wire  QDE ;
wire  QDF ;
wire  QDG ;
wire  QDH ;
wire  qea ;
wire  qeb ;
wire  qec ;
wire  qfa ;
wire  qfb ;
wire  qfc ;
wire  qfd ;
wire  qga ;
wire  qgb ;
wire  qgc ;
wire  qgd ;
wire  qma ;
wire  qmb ;
wire  qmc ;
wire  qmd ;
wire  qme ;
wire  qmf ;
wire  qmg ;
wire  qmh ;
wire  qna ;
wire  qnb ;
wire  qnc ;
wire  qnd ;
wire  qne ;
wire  qnf ;
wire  qng ;
wire  qnh ;
wire  qni ;
wire  qnj ;
wire  qra ;
wire  qrb ;
wire  QTA ;
wire  QTB ;
wire  QTC ;
wire  QTD ;
wire  SAA ;
wire  SAB ;
wire  SAC ;
wire  SAD ;
wire  SAE ;
wire  SAF ;
wire  SAG ;
wire  SAH ;
wire  SAI ;
wire  SAJ ;
wire  SAK ;
wire  SAL ;
wire  SAM ;
wire  SAN ;
wire  SAO ;
wire  SAP ;
wire  SAQ ;
wire  SAR ;
wire  SAS ;
wire  SAT ;
wire  SAU ;
wire  SAV ;
wire  SAW ;
wire  SAX ;
wire  SBA ;
wire  SBB ;
wire  SBC ;
wire  SBD ;
wire  SBE ;
wire  SBF ;
wire  SBG ;
wire  SBH ;
wire  SBI ;
wire  SBJ ;
wire  SBK ;
wire  SBL ;
wire  SBM ;
wire  SBN ;
wire  SBO ;
wire  SBP ;
wire  SBQ ;
wire  SBR ;
wire  SBS ;
wire  SBT ;
wire  SBU ;
wire  SBV ;
wire  SBW ;
wire  SBX ;
wire  SCA ;
wire  SCB ;
wire  SCC ;
wire  SCD ;
wire  SCE ;
wire  SCF ;
wire  SCG ;
wire  SCH ;
wire  SCI ;
wire  SCJ ;
wire  SCK ;
wire  SCL ;
wire  SCM ;
wire  SCN ;
wire  SCO ;
wire  SCP ;
wire  SCQ ;
wire  SCR ;
wire  SCS ;
wire  SCT ;
wire  SCU ;
wire  SCV ;
wire  SCW ;
wire  SCX ;
wire  SDA ;
wire  SDB ;
wire  SDC ;
wire  SDD ;
wire  SDE ;
wire  SDF ;
wire  SDG ;
wire  SDH ;
wire  SDI ;
wire  SDJ ;
wire  SDK ;
wire  SDL ;
wire  SDM ;
wire  SDN ;
wire  SDO ;
wire  SDP ;
wire  SDQ ;
wire  SDR ;
wire  SDS ;
wire  SDT ;
wire  SDU ;
wire  SDV ;
wire  SDW ;
wire  SDX ;
wire  SEA ;
wire  SEB ;
wire  SEC ;
wire  SED ;
wire  SEE ;
wire  SEF ;
wire  SEG ;
wire  SEH ;
wire  SEI ;
wire  SEJ ;
wire  SEK ;
wire  SEL ;
wire  SEM ;
wire  SEN ;
wire  SEO ;
wire  SEP ;
wire  SEQ ;
wire  SER ;
wire  SES ;
wire  SET ;
wire  SEU ;
wire  SEV ;
wire  SEW ;
wire  SEX ;
wire  SFA ;
wire  SFB ;
wire  SFC ;
wire  SFD ;
wire  SFE ;
wire  SFF ;
wire  SFG ;
wire  SFH ;
wire  SFI ;
wire  SFJ ;
wire  SFK ;
wire  SFL ;
wire  SFM ;
wire  SFN ;
wire  SFO ;
wire  SFP ;
wire  SFQ ;
wire  SFR ;
wire  SFS ;
wire  SFT ;
wire  SFU ;
wire  SFV ;
wire  SFW ;
wire  SFX ;
wire  SGA ;
wire  SGB ;
wire  SGC ;
wire  SGD ;
wire  SGE ;
wire  SGF ;
wire  SGG ;
wire  SGH ;
wire  SGI ;
wire  SGJ ;
wire  SGK ;
wire  SGL ;
wire  SGM ;
wire  SGN ;
wire  SGO ;
wire  SGP ;
wire  SGQ ;
wire  SGR ;
wire  SGS ;
wire  SGT ;
wire  SGU ;
wire  SGV ;
wire  SGW ;
wire  SGX ;
wire  SHA ;
wire  SHB ;
wire  SHC ;
wire  SHD ;
wire  SHE ;
wire  SHF ;
wire  SHG ;
wire  SHH ;
wire  SHI ;
wire  SHJ ;
wire  SHK ;
wire  SHL ;
wire  SHM ;
wire  SHN ;
wire  SHO ;
wire  SHP ;
wire  SHQ ;
wire  SHR ;
wire  SHS ;
wire  SHT ;
wire  SHU ;
wire  SHV ;
wire  SHW ;
wire  SHX ;
wire  SIA ;
wire  SIB ;
wire  SIC ;
wire  SID ;
wire  SIE ;
wire  SIF ;
wire  SIG ;
wire  SIH ;
wire  SII ;
wire  SIJ ;
wire  SIK ;
wire  SIL ;
wire  SIM ;
wire  SIN ;
wire  SIO ;
wire  SIP ;
wire  SIQ ;
wire  SIR ;
wire  SIS ;
wire  SIT ;
wire  SIU ;
wire  SIV ;
wire  SIW ;
wire  SIX ;
wire  SJA ;
wire  SJB ;
wire  SJC ;
wire  SJD ;
wire  SJE ;
wire  SJF ;
wire  SJG ;
wire  SJH ;
wire  SJI ;
wire  SJJ ;
wire  SJK ;
wire  SJL ;
wire  SJM ;
wire  SJN ;
wire  SJO ;
wire  SJP ;
wire  SJQ ;
wire  SJR ;
wire  SJS ;
wire  SJT ;
wire  SJU ;
wire  SJV ;
wire  SJW ;
wire  SJX ;
wire  taa ;
wire  tab ;
wire  tac ;
wire  tad ;
wire  tae ;
wire  taf ;
wire  tag ;
wire  tba ;
wire  tbb ;
wire  tbc ;
wire  tbd ;
wire  tbe ;
wire  tbf ;
wire  tca ;
wire  tcb ;
wire  tcc ;
wire  tcd ;
wire  tce ;
wire  tcf ;
wire  tcg ;
wire  tda ;
wire  tdb ;
wire  tdc ;
wire  tdd ;
wire  tde ;
wire  tdf ;
wire  tea ;
wire  teb ;
wire  tfa ;
wire  tfb ;
wire  tga ;
wire  tgb ;
wire  THA ;
wire  THB ;
wire  THC ;
wire  THD ;
wire  tia ;
wire  TIA ;
wire  tib ;
wire  TIB ;
wire  tic ;
wire  tid ;
wire  tie ;
wire  TIE ;
wire  tif ;
wire  TIF ;
wire  tja ;
wire  TJA ;
wire  tjb ;
wire  TJB ;
wire  tjc ;
wire  tjd ;
wire  tje ;
wire  TJE ;
wire  tjf ;
wire  TJF ;
wire  tka ;
wire  TKA ;
wire  tkb ;
wire  TKB ;
wire  tkc ;
wire  tkd ;
wire  tke ;
wire  TKE ;
wire  tkf ;
wire  TKF ;
wire  tla ;
wire  TLA ;
wire  tlb ;
wire  TLB ;
wire  tlc ;
wire  tld ;
wire  tle ;
wire  TLE ;
wire  tlf ;
wire  TLF ;
wire  tma ;
wire  tmb ;
wire  tmc ;
wire  tmd ;
wire  tna ;
wire  tnb ;
wire  tnc ;
wire  tnd ;
wire  waa ;
wire  wab ;
wire  wac ;
wire  wad ;
wire  wae ;
wire  waf ;
wire  wag ;
wire  wah ;
wire  wai ;
wire  waj ;
wire  wak ;
wire  wal ;
wire  wam ;
wire  wan ;
wire  wba ;
wire  wbb ;
wire  wbc ;
wire  wbd ;
wire  wbe ;
wire  wbf ;
wire  wbg ;
wire  wbh ;
wire  wbi ;
wire  wbj ;
wire  wbk ;
wire  wbl ;
wire  wbm ;
wire  wbn ;
wire  wca ;
wire  wcb ;
wire  wcc ;
wire  wcd ;
wire  wce ;
wire  wcf ;
wire  wcg ;
wire  wch ;
wire  wci ;
wire  wcj ;
wire  wck ;
wire  wcl ;
wire  wcm ;
wire  wcn ;
wire  wda ;
wire  wdb ;
wire  wdc ;
wire  wdd ;
wire  wde ;
wire  wdf ;
wire  wdg ;
wire  wdh ;
wire  wdi ;
wire  wdj ;
wire  wdk ;
wire  wdl ;
wire  wdm ;
wire  wdn ;
wire  xaa ;
wire  XAA ;
wire  xab ;
wire  XAB ;
wire  ZZI ;
wire  ZZO ;
assign ZZI = 1'b1;
assign ZZO = 1'b0;
assign PAA = ~paa;  //complement 
assign PBA = ~pba;  //complement 
assign PCA = ~pca;  //complement 
assign PDA = ~pda;  //complement 
assign PEA = ~pea;  //complement 
assign PFA = ~pfa;  //complement 
assign PGA = ~pga;  //complement 
assign PHA = ~pha;  //complement 
assign PIA = ~pia;  //complement 
assign PJA = ~pja;  //complement 
assign LCA =  CEA & CEB  |  CEA & CGB  |  CEB & CGB  ; 
assign lca = ~LCA; //complement 
assign PAB = ~pab;  //complement 
assign PBB = ~pbb;  //complement 
assign PCB = ~pcb;  //complement 
assign PDB = ~pdb;  //complement 
assign PEB = ~peb;  //complement 
assign PFB = ~pfb;  //complement 
assign PGB = ~pgb;  //complement 
assign PHB = ~phb;  //complement 
assign PIB = ~pib;  //complement 
assign PJB = ~pjb;  //complement 
assign DAB = ~dab;  //complement 
assign PAC = ~pac;  //complement 
assign PBC = ~pbc;  //complement 
assign PCC = ~pcc;  //complement 
assign PDC = ~pdc;  //complement 
assign PEC = ~pec;  //complement 
assign PFC = ~pfc;  //complement 
assign PGC = ~pgc;  //complement 
assign PHC = ~phc;  //complement 
assign PIC = ~pic;  //complement 
assign PJC = ~pjc;  //complement 
assign DAC = ~dac;  //complement 
assign DAD = ~dad;  //complement 
assign PAD = ~pad;  //complement 
assign PBD = ~pbd;  //complement 
assign PCD = ~pcd;  //complement 
assign PDD = ~pdd;  //complement 
assign PED = ~ped;  //complement 
assign PFD = ~pfd;  //complement 
assign PGD = ~pgd;  //complement 
assign PHD = ~phd;  //complement 
assign PID = ~pid;  //complement 
assign PJD = ~pjd;  //complement 
assign LCB =  CEC & CGC & CED  |  CEC & CGC & CGD  |  CED & CGD  ; 
assign lcb = ~LCB; //complement 
assign PAE = ~pae;  //complement 
assign PBE = ~pbe;  //complement 
assign PCE = ~pce;  //complement 
assign PDE = ~pde;  //complement 
assign PEE = ~pee;  //complement 
assign PFE = ~pfe;  //complement 
assign PGE = ~pge;  //complement 
assign PHE = ~phe;  //complement 
assign PIE = ~pie;  //complement 
assign PJE = ~pje;  //complement 
assign lbb =  cac & ccc  |  cad & ccd  ; 
assign LBB = ~lbb;  //complement 
assign ldb =  cec & cgc  |  ced & cgd  ; 
assign LDB = ~ldb;  //complement 
assign PAF = ~paf;  //complement 
assign PBF = ~pbf;  //complement 
assign PCF = ~pcf;  //complement 
assign PDF = ~pdf;  //complement 
assign PEF = ~pef;  //complement 
assign PFF = ~pff;  //complement 
assign PGF = ~pgf;  //complement 
assign PHF = ~phf;  //complement 
assign PIF = ~pif;  //complement 
assign PJF = ~pjf;  //complement 
assign PAR = ~par;  //complement 
assign PBR = ~pbr;  //complement 
assign PCR = ~pcr;  //complement 
assign PDR = ~pdr;  //complement 
assign PAM = ~pam;  //complement 
assign PBM = ~pbm;  //complement 
assign PCM = ~pcm;  //complement 
assign PDM = ~pdm;  //complement 
assign PEM = ~pem;  //complement 
assign PFM = ~pfm;  //complement 
assign PGM = ~pgm;  //complement 
assign PHM = ~phm;  //complement 
assign PJM = ~pjm;  //complement 
assign PIM = ~pim;  //complement 
assign PER = ~per;  //complement 
assign PFR = ~pfr;  //complement 
assign PGR = ~pgr;  //complement 
assign PHR = ~phr;  //complement 
assign PAN = ~pan;  //complement 
assign PBN = ~pbn;  //complement 
assign PCN = ~pcn;  //complement 
assign PDN = ~pdn;  //complement 
assign PEN = ~pen;  //complement 
assign PFN = ~pfn;  //complement 
assign PGN = ~pgn;  //complement 
assign PHN = ~phn;  //complement 
assign PIN = ~pin;  //complement 
assign PJN = ~pjn;  //complement 
assign PIR = ~pir;  //complement 
assign PJR = ~pjr;  //complement 
assign QAA = ~qaa;  //complement 
assign QAB = ~qab;  //complement 
assign cea = ~CEA;  //complement 
assign CGB = ~cgb;  //complement 
assign caa = ~CAA;  //complement 
assign CCB = ~ccb;  //complement 
assign eab = ~EAB;  //complement 
assign ebb = ~EBB;  //complement 
assign cab = ~CAB;  //complement 
assign CCC = ~ccc;  //complement 
assign eac = ~EAC;  //complement 
assign ebc = ~EBC;  //complement 
assign cec = ~CEC;  //complement 
assign CGD = ~cgd;  //complement 
assign cac = ~CAC;  //complement 
assign CCD = ~ccd;  //complement 
assign ead = ~EAD;  //complement 
assign ebd = ~EBD;  //complement 
assign bee =  AAD & acd & aed  |  aad & ACD & aed  |  aad & acd & AED  |  aad & acd & aed  ; 
assign BEE = ~bee;  //complement 
assign ced = ~CED;  //complement 
assign CGE = ~cge;  //complement 
assign cad = ~CAD;  //complement 
assign CCE = ~cce;  //complement 
assign tna = ~TNA;  //complement 
assign tnb = ~TNB;  //complement 
assign tnc = ~TNC;  //complement 
assign tnd = ~TND;  //complement 
assign LAB =  CAC & CCC & CAD  |  CAC & CCC & CCD  |  CAD & CCD  ; 
assign lab = ~LAB; //complement 
assign LAA =  CAA & CAB  |  CAA & CCB  |  CAB & CCB  ; 
assign laa = ~LAA; //complement 
assign THA = ~tha;  //complement 
assign THB = ~thb;  //complement 
assign THC = ~thc;  //complement 
assign THD = ~thd;  //complement 
assign jac =  dab  ; 
assign JAC = ~jac;  //complement 
assign jad =  dac & dab  |  dac & eac  ; 
assign JAD = ~jad;  //complement 
assign faa = ~FAA;  //complement 
assign fab = ~FAB;  //complement 
assign jae =  dab & dac & dad  |  eac & dac & dad  |  ead & dad  ; 
assign JAE = ~jae; //complement 
assign fac = ~FAC;  //complement 
assign fad = ~FAD;  //complement 
assign KAB =  fac & fad & fae & faf  ; 
assign kab = ~KAB;  //complement  
assign ceb = ~CEB;  //complement 
assign CGC = ~cgc;  //complement 
assign fae = ~FAE;  //complement 
assign faf = ~FAF;  //complement 
assign BAA =  AAA & aca & aea  |  aaa & ACA & aea  |  aaa & aca & AEA  |  AAA & ACA & AEA  ; 
assign baa = ~BAA; //complement 
assign bcb =  AAA & aca & aea  |  aaa & ACA & aea  |  aaa & aca & AEA  |  aaa & aca & aea  ; 
assign BCB = ~bcb;  //complement 
assign aaa = ~AAA;  //complement 
assign aab = ~AAB;  //complement 
assign aga = ~AGA;  //complement 
assign agb = ~AGB;  //complement 
assign AIA = ~aia;  //complement 
assign AIB = ~aib;  //complement 
assign BAB =  AAB & acb & aeb  |  aab & ACB & aeb  |  aab & acb & AEB  |  AAB & ACB & AEB  ; 
assign bab = ~BAB; //complement 
assign bcc =  AAB & acb & aeb  |  aab & ACB & aeb  |  aab & acb & AEB  |  aab & acb & aeb  ; 
assign BCC = ~bcc;  //complement 
assign aca = ~ACA;  //complement 
assign acb = ~ACB;  //complement 
assign aea = ~AEA;  //complement 
assign aeb = ~AEB;  //complement 
assign AKA = ~aka;  //complement 
assign AKB = ~akb;  //complement 
assign BAC =  AAC & acc & aec  |  aac & ACC & aec  |  aac & acc & AEC  |  AAC & ACC & AEC  ; 
assign bac = ~BAC; //complement 
assign bcd =  AAC & acc & aec  |  aac & ACC & aec  |  aac & acc & AEC  |  aac & acc & aec  ; 
assign BCD = ~bcd;  //complement 
assign aac = ~AAC;  //complement 
assign aad = ~AAD;  //complement 
assign agc = ~AGC;  //complement 
assign agd = ~AGD;  //complement 
assign AIC = ~aic;  //complement 
assign AID = ~aid;  //complement 
assign BAD =  AAD & acd & aed  |  aad & ACD & aed  |  aad & acd & AED  |  AAD & ACD & AED  ; 
assign bad = ~BAD; //complement 
assign bce =  AAD & acd & aed  |  aad & ACD & aed  |  aad & acd & AED  |  aad & acd & aed  ; 
assign BCE = ~bce;  //complement 
assign acc = ~ACC;  //complement 
assign acd = ~ACD;  //complement 
assign aec = ~AEC;  //complement 
assign aed = ~AED;  //complement 
assign AKC = ~akc;  //complement 
assign AKD = ~akd;  //complement 
assign tma = ~TMA;  //complement 
assign tmb = ~TMB;  //complement 
assign tmc = ~TMC;  //complement 
assign tmd = ~TMD;  //complement 
assign qac = ~QAC;  //complement 
assign tga = ~TGA;  //complement 
assign tgb = ~TGB;  //complement 
assign ohe = ~OHE;  //complement 
assign oam = ~OAM;  //complement 
assign wam = ~WAM;  //complement 
assign qma = ~QMA;  //complement 
assign qme = ~QME;  //complement 
assign TIA =  QBA & qma & qde & wak & wal  ; 
assign tia = ~TIA;  //complement  
assign oaa = ~OAA;  //complement 
assign waa = ~WAA;  //complement 
assign oab = ~OAB;  //complement 
assign wab = ~WAB;  //complement 
assign qba = ~QBA;  //complement 
assign qbe = ~QBE;  //complement 
assign KBA =  QBA & qma & QDA  ; 
assign kba = ~KBA;  //complement 
assign TIE =  QTA & qde  ; 
assign tie = ~TIE;  //complement 
assign oac = ~OAC;  //complement 
assign wac = ~WAC;  //complement 
assign oad = ~OAD;  //complement 
assign wad = ~WAD;  //complement 
assign qga = ~QGA;  //complement 
assign tic = ~TIC;  //complement 
assign tid = ~TID;  //complement 
assign QTA = ~qta;  //complement 
assign OHA = ~oha;  //complement 
assign oae = ~OAE;  //complement 
assign wae = ~WAE;  //complement 
assign oaf = ~OAF;  //complement 
assign waf = ~WAF;  //complement 
assign PAG = ~pag;  //complement 
assign PBG = ~pbg;  //complement 
assign PCG = ~pcg;  //complement 
assign PDG = ~pdg;  //complement 
assign PEG = ~peg;  //complement 
assign PFG = ~pfg;  //complement 
assign PGG = ~pgg;  //complement 
assign PHG = ~phg;  //complement 
assign PIG = ~pig;  //complement 
assign PIH = ~pih;  //complement 
assign PJG = ~pjg;  //complement 
assign LCC =  CEE & CGE & CEF  |  CEE & CGE & CGF  |  CEF & CGF  ; 
assign lcc = ~LCC; //complement 
assign PAH = ~pah;  //complement 
assign PBH = ~pbh;  //complement 
assign PCH = ~pch;  //complement 
assign PDH = ~pdh;  //complement 
assign PEH = ~peh;  //complement 
assign PFH = ~pfh;  //complement 
assign PGH = ~pgh;  //complement 
assign PHH = ~phh;  //complement 
assign ldc =  cee & cge  |  cef & cgf  ; 
assign LDC = ~ldc;  //complement 
assign ldd =  ceg & cgg  |  ceh & cgh  ; 
assign LDD = ~ldd;  //complement 
assign DAE = ~dae;  //complement 
assign DAF = ~daf;  //complement 
assign PAI = ~pai;  //complement 
assign PBI = ~pbi;  //complement 
assign PCI = ~pci;  //complement 
assign PDI = ~pdi;  //complement 
assign PEI = ~pei;  //complement 
assign PFI = ~pfi;  //complement 
assign PGI = ~pgi;  //complement 
assign PHI = ~phi;  //complement 
assign PII = ~pii;  //complement 
assign PJI = ~pji;  //complement 
assign PJH = ~pjh;  //complement 
assign DAG = ~dag;  //complement 
assign DAH = ~dah;  //complement 
assign PAJ = ~paj;  //complement 
assign PBJ = ~pbj;  //complement 
assign PCJ = ~pcj;  //complement 
assign PDJ = ~pdj;  //complement 
assign PEJ = ~pej;  //complement 
assign PFJ = ~pfj;  //complement 
assign PGJ = ~pgj;  //complement 
assign PHJ = ~phj;  //complement 
assign LCD =  CEG & CGG & CEH  |  CEG & CGG & CGH  |  CEH & CGH  ; 
assign lcd = ~LCD; //complement 
assign JAG =  DAB & EAC & EAD & EAE & EAF  |  DAC & EAD & EAE & EAF  |  DAD & EAE & EAF  |  DAE & EAF  |  DAF  ; 
assign jag = ~JAG;  //complement 
assign PAK = ~pak;  //complement 
assign PBK = ~pbk;  //complement 
assign PCK = ~pck;  //complement 
assign PDK = ~pdk;  //complement 
assign PEK = ~pek;  //complement 
assign PFK = ~pfk;  //complement 
assign PGK = ~pgk;  //complement 
assign PHK = ~phk;  //complement 
assign PIK = ~pik;  //complement 
assign PJK = ~pjk;  //complement 
assign PIJ = ~pij;  //complement 
assign PJJ = ~pjj;  //complement 
assign fem = ~FEM;  //complement 
assign fen = ~FEN;  //complement 
assign PAQ = ~paq;  //complement 
assign PBQ = ~pbq;  //complement 
assign PCQ = ~pcq;  //complement 
assign PDQ = ~pdq;  //complement 
assign PEQ = ~peq;  //complement 
assign PFQ = ~pfq;  //complement 
assign PGQ = ~pgq;  //complement 
assign PHQ = ~phq;  //complement 
assign qnb = ~QNB;  //complement 
assign qnc = ~QNC;  //complement 
assign qnd = ~QND;  //complement 
assign qne = ~QNE;  //complement 
assign qnf = ~QNF;  //complement 
assign qng = ~QNG;  //complement 
assign qnh = ~QNH;  //complement 
assign qni = ~QNI;  //complement 
assign PAO = ~pao;  //complement 
assign PBO = ~pbo;  //complement 
assign PCO = ~pco;  //complement 
assign PDO = ~pdo;  //complement 
assign PEO = ~peo;  //complement 
assign PFO = ~pfo;  //complement 
assign PGO = ~pgo;  //complement 
assign PHO = ~pho;  //complement 
assign PJO = ~pjo;  //complement 
assign PIO = ~pio;  //complement 
assign mba = ~MBA;  //complement 
assign PAP = ~pap;  //complement 
assign PBP = ~pbp;  //complement 
assign PCP = ~pcp;  //complement 
assign PDP = ~pdp;  //complement 
assign PEP = ~pep;  //complement 
assign PFP = ~pfp;  //complement 
assign PGP = ~pgp;  //complement 
assign PHP = ~php;  //complement 
assign PIP = ~pip;  //complement 
assign PJP = ~pjp;  //complement 
assign qnj = ~QNJ;  //complement 
assign eae = ~EAE;  //complement 
assign ebe = ~EBE;  //complement 
assign cee = ~CEE;  //complement 
assign CGF = ~cgf;  //complement 
assign cae = ~CAE;  //complement 
assign CCF = ~ccf;  //complement 
assign eaf = ~EAF;  //complement 
assign ebf = ~EBF;  //complement 
assign cef = ~CEF;  //complement 
assign CGG = ~cgg;  //complement 
assign caf = ~CAF;  //complement 
assign CCG = ~ccg;  //complement 
assign eag = ~EAG;  //complement 
assign ebg = ~EBG;  //complement 
assign ceg = ~CEG;  //complement 
assign CGH = ~cgh;  //complement 
assign cag = ~CAG;  //complement 
assign CCH = ~cch;  //complement 
assign eah = ~EAH;  //complement 
assign ebh = ~EBH;  //complement 
assign bei =  AAH & ach & aeh  |  aah & ACH & aeh  |  aah & ach & AEH  |  aah & ach & aeh  ; 
assign BEI = ~bei;  //complement 
assign ceh = ~CEH;  //complement 
assign CGI = ~cgi;  //complement 
assign cah = ~CAH;  //complement 
assign CCI = ~cci;  //complement 
assign JFA =  FAM  |  fca & fen & TNA  |  fda & FEN & TNB  ; 
assign jfa = ~JFA; //complement 
assign lbc =  cae & cce  |  caf & ccf  ; 
assign LBC = ~lbc;  //complement 
assign lbd =  cag & ccg  |  cah & cch  ; 
assign LBD = ~lbd;  //complement 
assign LAD =  CAG & CCG & CAH  |  CAG & CCG & CCH  |  CAH & CCH  ; 
assign lad = ~LAD; //complement 
assign LAC =  CAE & CCE & CAF  |  CAE & CCE & CCF  |  CAF & CCF  ; 
assign lac = ~LAC; //complement 
assign JAF =  DAB & EAC & EAD & EAE  |  DAC & EAD & EAE  |  DAD & EAE  |  DAE  ; 
assign jaf = ~JAF;  //complement 
assign fag = ~FAG;  //complement 
assign fah = ~FAH;  //complement 
assign qna = ~QNA;  //complement 
assign fai = ~FAI;  //complement 
assign faj = ~FAJ;  //complement 
assign fea = ~FEA;  //complement 
assign fei = ~FEI;  //complement 
assign fak = ~FAK;  //complement 
assign fal = ~FAL;  //complement 
assign KAA =  QNA & QMA  |  QNJ & QMA  |  QEB  ; 
assign kaa = ~KAA;  //complement 
assign BAE =  AAE & ace & aee  |  aae & ACE & aee  |  aae & ace & AEE  |  AAE & ACE & AEE  ; 
assign bae = ~BAE; //complement 
assign bcf =  AAE & ace & aee  |  aae & ACE & aee  |  aae & ace & AEE  |  aae & ace & aee  ; 
assign BCF = ~bcf;  //complement 
assign aae = ~AAE;  //complement 
assign aaf = ~AAF;  //complement 
assign age = ~AGE;  //complement 
assign agf = ~AGF;  //complement 
assign AIE = ~aie;  //complement 
assign AIF = ~aif;  //complement 
assign BAF =  AAF & acf & aef  |  aaf & ACF & aef  |  aaf & acf & AEF  |  AAF & ACF & AEF  ; 
assign baf = ~BAF; //complement 
assign bcg =  AAF & acf & aef  |  aaf & ACF & aef  |  aaf & acf & AEF  |  aaf & acf & aef  ; 
assign BCG = ~bcg;  //complement 
assign ace = ~ACE;  //complement 
assign acf = ~ACF;  //complement 
assign aee = ~AEE;  //complement 
assign aef = ~AEF;  //complement 
assign AKE = ~ake;  //complement 
assign AKF = ~akf;  //complement 
assign BAG =  AAG & acg & aeg  |  aag & ACG & aeg  |  aag & acg & AEG  |  AAG & ACG & AEG  ; 
assign bag = ~BAG; //complement 
assign bch =  AAG & acg & aeg  |  aag & ACG & aeg  |  aag & acg & AEG  |  aag & acg & aeg  ; 
assign BCH = ~bch;  //complement 
assign aag = ~AAG;  //complement 
assign aah = ~AAH;  //complement 
assign agg = ~AGG;  //complement 
assign agh = ~AGH;  //complement 
assign AIG = ~aig;  //complement 
assign AIH = ~aih;  //complement 
assign BAH =  AAH & ach & aeh  |  aah & ACH & aeh  |  aah & ach & AEH  |  AAH & ACH & AEH  ; 
assign bah = ~BAH; //complement 
assign bci =  AAH & ach & aeh  |  aah & ACH & aeh  |  aah & ach & AEH  |  aah & ach & aeh  ; 
assign BCI = ~bci;  //complement 
assign acg = ~ACG;  //complement 
assign ach = ~ACH;  //complement 
assign aeg = ~AEG;  //complement 
assign aeh = ~AEH;  //complement 
assign AKG = ~akg;  //complement 
assign AKH = ~akh;  //complement 
assign tac = ~TAC;  //complement 
assign tad = ~TAD;  //complement 
assign tag = ~TAG;  //complement 
assign taa = ~TAA;  //complement 
assign tab = ~TAB;  //complement 
assign oia = ~OIA;  //complement 
assign tae = ~TAE;  //complement 
assign taf = ~TAF;  //complement 
assign oan = ~OAN;  //complement 
assign wan = ~WAN;  //complement 
assign oie = ~OIE;  //complement 
assign ola = ~OLA;  //complement 
assign qca = ~QCA;  //complement 
assign TIB =  QBE & qme & qda & wak & wal  ; 
assign tib = ~TIB;  //complement  
assign KCA =  QBE & qme & qda  ; 
assign kca = ~KCA;  //complement 
assign oag = ~OAG;  //complement 
assign wag = ~WAG;  //complement 
assign oah = ~OAH;  //complement 
assign wah = ~WAH;  //complement 
assign QDA = ~qda;  //complement 
assign QDE = ~qde;  //complement 
assign KBE =  QBE & qme  ; 
assign kbe = ~KBE;  //complement 
assign TIF =  QTA & qda  ; 
assign tif = ~TIF;  //complement 
assign oai = ~OAI;  //complement 
assign wai = ~WAI;  //complement 
assign oaj = ~OAJ;  //complement 
assign waj = ~WAJ;  //complement 
assign qeb = ~QEB;  //complement 
assign OFA = ~ofa;  //complement 
assign qfa = ~QFA;  //complement 
assign oak = ~OAK;  //complement 
assign wak = ~WAK;  //complement 
assign oal = ~OAL;  //complement 
assign wal = ~WAL;  //complement 
assign LCE =  CEI & CGI & CEJ  |  CEI & CGI & CGJ  |  CEJ & CGJ  ; 
assign lce = ~LCE; //complement 
assign JDB =  DAH  ; 
assign jdb = ~JDB;  //complement 
assign JDC =  EAI & DAH  |  DAI  ; 
assign jdc = ~JDC;  //complement 
assign DAI = ~dai;  //complement 
assign DAJ = ~daj;  //complement 
assign lde =  cei & cgi  |  cej & cgj  ; 
assign LDE = ~lde;  //complement 
assign ldf =  cek & cgk  |  cel & cgl  ; 
assign LDF = ~ldf;  //complement 
assign JDD =  DAH & EAI & EAJ  |  DAI & EAJ  |  DAJ  ; 
assign jdd = ~JDD; //complement 
assign DAK = ~dak;  //complement 
assign DAL = ~dal;  //complement 
assign PIQ = ~piq;  //complement 
assign PJQ = ~pjq;  //complement 
assign LCF =  CEK & CGK & CEL  |  CEK & CGK & CGL  |  CEL & CGL  ; 
assign lcf = ~LCF; //complement 
assign jeb =  dah & eah & eah  ; 
assign JEB = ~jeb;  //complement 
assign jec =  dai & dah & eah  |  dai & eai  ; 
assign JEC = ~jec;  //complement 
assign jed =  eah & dah & dai & daj  |  eai & dai & daj  |  eaj & daj  ; 
assign JED = ~jed;  //complement 
assign SAA = ~saa;  //complement 
assign SBA = ~sba;  //complement 
assign SCA = ~sca;  //complement 
assign SDA = ~sda;  //complement 
assign SEA = ~sea;  //complement 
assign SFA = ~sfa;  //complement 
assign SGA = ~sga;  //complement 
assign SHA = ~sha;  //complement 
assign SIA = ~sia;  //complement 
assign SJA = ~sja;  //complement 
assign fca = ~FCA;  //complement 
assign fda = ~FDA;  //complement 
assign SAB = ~sab;  //complement 
assign SBB = ~sbb;  //complement 
assign SCB = ~scb;  //complement 
assign SDB = ~sdb;  //complement 
assign SEB = ~seb;  //complement 
assign SFB = ~sfb;  //complement 
assign SGB = ~sgb;  //complement 
assign SHB = ~shb;  //complement 
assign SIB = ~sib;  //complement 
assign SJB = ~sjb;  //complement 
assign fcb = ~FCB;  //complement 
assign fdb = ~FDB;  //complement 
assign SAC = ~sac;  //complement 
assign SBC = ~sbc;  //complement 
assign SCC = ~scc;  //complement 
assign SDC = ~sdc;  //complement 
assign SEC = ~sec;  //complement 
assign SFC = ~sfc;  //complement 
assign SGC = ~sgc;  //complement 
assign SHC = ~shc;  //complement 
assign fcc = ~FCC;  //complement 
assign fdc = ~FDC;  //complement 
assign SAD = ~sad;  //complement 
assign SBD = ~sbd;  //complement 
assign SCD = ~scd;  //complement 
assign SDD = ~sdd;  //complement 
assign SED = ~sed;  //complement 
assign SFD = ~sfd;  //complement 
assign SGD = ~sgd;  //complement 
assign SHD = ~shd;  //complement 
assign SID = ~sid;  //complement 
assign SJD = ~sjd;  //complement 
assign SIC = ~sic;  //complement 
assign SJC = ~sjc;  //complement 
assign fcd = ~FCD;  //complement 
assign fdd = ~FDD;  //complement 
assign eai = ~EAI;  //complement 
assign cei = ~CEI;  //complement 
assign CGJ = ~cgj;  //complement 
assign cai = ~CAI;  //complement 
assign CCJ = ~ccj;  //complement 
assign eaj = ~EAJ;  //complement 
assign cej = ~CEJ;  //complement 
assign CGK = ~cgk;  //complement 
assign caj = ~CAJ;  //complement 
assign CCK = ~cck;  //complement 
assign eak = ~EAK;  //complement 
assign cek = ~CEK;  //complement 
assign CGL = ~cgl;  //complement 
assign cak = ~CAK;  //complement 
assign CCL = ~ccl;  //complement 
assign eal = ~EAL;  //complement 
assign bem =  AAL & acl & ael  |  aal & ACL & ael  |  aal & acl & AEL  |  aal & acl & ael  ; 
assign BEM = ~bem;  //complement 
assign cel = ~CEL;  //complement 
assign CGM = ~cgm;  //complement 
assign cal = ~CAL;  //complement 
assign CCM = ~ccm;  //complement 
assign JFB =  FAN  |  FCA & fem & TNC  |  FDA & FEM & TND  ; 
assign jfb = ~JFB; //complement 
assign LAF =  CAK & CCK & CAL  |  CAK & CCK & CCL  |  CAL & CCL  ; 
assign laf = ~LAF; //complement 
assign LAE =  CAI & CCI & CAJ  |  CAI & CCI & CCJ  |  CAJ & CCJ  ; 
assign lae = ~LAE; //complement 
assign haa = ~HAA;  //complement 
assign oea = ~OEA;  //complement 
assign fam = ~FAM;  //complement 
assign fan = ~FAN;  //complement 
assign hac = ~HAC;  //complement 
assign oec = ~OEC;  //complement 
assign lbe =  cai & cci  |  caj & ccj  ; 
assign LBE = ~lbe;  //complement 
assign lbf =  cak & cck  |  cal & ccl  ; 
assign LBF = ~lbf;  //complement 
assign hab = ~HAB;  //complement 
assign oeb = ~OEB;  //complement 
assign FFB = ~ffb;  //complement 
assign FFJ = ~ffj;  //complement 
assign maa = ~MAA;  //complement 
assign feb = ~FEB;  //complement 
assign fej = ~FEJ;  //complement 
assign gaa =  fea  ; 
assign GAA = ~gaa;  //complement 
assign had = ~HAD;  //complement 
assign oed = ~OED;  //complement 
assign BAI =  AAI & aci & aei  |  aai & ACI & aei  |  aai & aci & AEI  |  AAI & ACI & AEI  ; 
assign bai = ~BAI; //complement 
assign bcj =  AAI & aci & aei  |  aai & ACI & aei  |  aai & aci & AEI  |  aai & aci & aei  ; 
assign BCJ = ~bcj;  //complement 
assign aai = ~AAI;  //complement 
assign aaj = ~AAJ;  //complement 
assign agi = ~AGI;  //complement 
assign agj = ~AGJ;  //complement 
assign AII = ~aii;  //complement 
assign AIJ = ~aij;  //complement 
assign BAJ =  AAJ & acj & aej  |  aaj & ACJ & aej  |  aaj & acj & AEJ  |  AAJ & ACJ & AEJ  ; 
assign baj = ~BAJ; //complement 
assign bck =  AAJ & acj & aej  |  aaj & ACJ & aej  |  aaj & acj & AEJ  |  aaj & acj & aej  ; 
assign BCK = ~bck;  //complement 
assign aci = ~ACI;  //complement 
assign acj = ~ACJ;  //complement 
assign aei = ~AEI;  //complement 
assign aej = ~AEJ;  //complement 
assign AKI = ~aki;  //complement 
assign AKJ = ~akj;  //complement 
assign BAK =  AAK & ack & aek  |  aak & ACK & aek  |  aak & ack & AEK  |  AAK & ACK & AEK  ; 
assign bak = ~BAK; //complement 
assign bcl =  AAK & ack & aek  |  aak & ACK & aek  |  aak & ack & AEK  |  aak & ack & aek  ; 
assign BCL = ~bcl;  //complement 
assign aak = ~AAK;  //complement 
assign aal = ~AAL;  //complement 
assign agk = ~AGK;  //complement 
assign agl = ~AGL;  //complement 
assign AIK = ~aik;  //complement 
assign AIL = ~ail;  //complement 
assign BAL =  AAL & acl & ael  |  aal & ACL & ael  |  aal & acl & AEL  |  AAL & ACL & AEL  ; 
assign bal = ~BAL; //complement 
assign bcm =  AAL & acl & ael  |  aal & ACL & ael  |  aal & acl & AEL  |  aal & acl & ael  ; 
assign BCM = ~bcm;  //complement 
assign ack = ~ACK;  //complement 
assign acl = ~ACL;  //complement 
assign aek = ~AEK;  //complement 
assign ael = ~AEL;  //complement 
assign AKK = ~akk;  //complement 
assign AKL = ~akl;  //complement 
assign tba = ~TBA;  //complement 
assign tbb = ~TBB;  //complement 
assign tbc = ~TBC;  //complement 
assign tbd = ~TBD;  //complement 
assign tbe = ~TBE;  //complement 
assign tbf = ~TBF;  //complement 
assign obm = ~OBM;  //complement 
assign wbm = ~WBM;  //complement 
assign qmb = ~QMB;  //complement 
assign qmf = ~QMF;  //complement 
assign TJA =  QBB & qmb & qdf & wbk & wbl  ; 
assign tja = ~TJA;  //complement  
assign oba = ~OBA;  //complement 
assign wba = ~WBA;  //complement 
assign obb = ~OBB;  //complement 
assign wbb = ~WBB;  //complement 
assign qbb = ~QBB;  //complement 
assign qbf = ~QBF;  //complement 
assign KBB =  QBB & qmb & QDB  ; 
assign kbb = ~KBB;  //complement 
assign TJE =  QTB & qdf  ; 
assign tje = ~TJE;  //complement 
assign obc = ~OBC;  //complement 
assign wbc = ~WBC;  //complement 
assign obd = ~OBD;  //complement 
assign wbd = ~WBD;  //complement 
assign qgb = ~QGB;  //complement 
assign tjc = ~TJC;  //complement 
assign tjd = ~TJD;  //complement 
assign QTB = ~qtb;  //complement 
assign OHB = ~ohb;  //complement 
assign obe = ~OBE;  //complement 
assign wbe = ~WBE;  //complement 
assign obf = ~OBF;  //complement 
assign wbf = ~WBF;  //complement 
assign LCG =  CEM & CGM & CEN  |  CEM & CGM & CGN  |  CEN & CGN  ; 
assign lcg = ~LCG; //complement 
assign JDF =  DAL  ; 
assign jdf = ~JDF;  //complement 
assign JDG =  EAM & DAL  |  DAM  ; 
assign jdg = ~JDG;  //complement 
assign DAM = ~dam;  //complement 
assign DAN = ~dan;  //complement 
assign ldg =  cem & cgm  |  cen & cgn  ; 
assign LDG = ~ldg;  //complement 
assign ldh =  ceo & cgo  |  cep & cgp  ; 
assign LDH = ~ldh;  //complement 
assign JDH =  DAL & EAM & EAN  |  DAM & EAN  |  DAN  ; 
assign jdh = ~JDH;  //complement 
assign DAO = ~dao;  //complement 
assign DAP = ~dap;  //complement 
assign LCH =  CEO & CGO & CEP  |  CEO & CGO & CGP  |  CEP & CGP  ; 
assign lch = ~LCH; //complement 
assign jef =  dal & eal & eal  ; 
assign JEF = ~jef;  //complement 
assign jeg =  dam & dal & eal  |  dam & eam  ; 
assign JEG = ~jeg;  //complement 
assign jeh =  eal & dal & dam & dan  |  eam & dam & dan  |  ean & dan  ; 
assign JEH = ~jeh;  //complement 
assign SAE = ~sae;  //complement 
assign SBE = ~sbe;  //complement 
assign SCE = ~sce;  //complement 
assign SDE = ~sde;  //complement 
assign SEE = ~see;  //complement 
assign SFE = ~sfe;  //complement 
assign SGE = ~sge;  //complement 
assign SHE = ~she;  //complement 
assign SIE = ~sie;  //complement 
assign SJE = ~sje;  //complement 
assign fce = ~FCE;  //complement 
assign fde = ~FDE;  //complement 
assign SAF = ~saf;  //complement 
assign SBF = ~sbf;  //complement 
assign SCF = ~scf;  //complement 
assign SDF = ~sdf;  //complement 
assign SEF = ~sef;  //complement 
assign SFF = ~sff;  //complement 
assign SGF = ~sgf;  //complement 
assign SHF = ~shf;  //complement 
assign SIF = ~sif;  //complement 
assign SIG = ~sig;  //complement 
assign fcf = ~FCF;  //complement 
assign fdf = ~FDF;  //complement 
assign SAG = ~sag;  //complement 
assign SBG = ~sbg;  //complement 
assign SCG = ~scg;  //complement 
assign SDG = ~sdg;  //complement 
assign SEG = ~seg;  //complement 
assign SFG = ~sfg;  //complement 
assign SGG = ~sgg;  //complement 
assign SHG = ~shg;  //complement 
assign SJG = ~sjg;  //complement 
assign fcg = ~FCG;  //complement 
assign fdg = ~FDG;  //complement 
assign SAH = ~sah;  //complement 
assign SBH = ~sbh;  //complement 
assign SCH = ~sch;  //complement 
assign SDH = ~sdh;  //complement 
assign SEH = ~seh;  //complement 
assign SFH = ~sfh;  //complement 
assign SGH = ~sgh;  //complement 
assign SHH = ~shh;  //complement 
assign SIH = ~sih;  //complement 
assign SJH = ~sjh;  //complement 
assign SJF = ~sjf;  //complement 
assign fch = ~FCH;  //complement 
assign fdh = ~FDH;  //complement 
assign eam = ~EAM;  //complement 
assign cem = ~CEM;  //complement 
assign CGN = ~cgn;  //complement 
assign cam = ~CAM;  //complement 
assign CCN = ~ccn;  //complement 
assign ean = ~EAN;  //complement 
assign cen = ~CEN;  //complement 
assign CGO = ~cgo;  //complement 
assign can = ~CAN;  //complement 
assign CCO = ~cco;  //complement 
assign eao = ~EAO;  //complement 
assign ceo = ~CEO;  //complement 
assign CGP = ~cgp;  //complement 
assign eap = ~EAP;  //complement 
assign bfa =  AAP & acp & aep  |  aap & ACP & aep  |  aap & acp & AEP  |  aap & acp & aep  ; 
assign BFA = ~bfa;  //complement 
assign cep = ~CEP;  //complement 
assign CHA = ~cha;  //complement 
assign cap = ~CAP;  //complement 
assign CDA = ~cda;  //complement 
assign lbg =  cam & ccm  |  can & ccn  ; 
assign LBG = ~lbg;  //complement 
assign lbh =  cao & cco  |  cap & ccp  ; 
assign LBH = ~lbh;  //complement 
assign LAH =  CAO & CCO & CAP  |  CAO & CCO & CCP  |  CAP & CCP  ; 
assign lah = ~LAH; //complement 
assign LAG =  CAM & CCM & CAN  |  CAM & CCM & CCN  |  CAN & CCN  ; 
assign lag = ~LAG; //complement 
assign hae = ~HAE;  //complement 
assign oee = ~OEE;  //complement 
assign mbb = ~MBB;  //complement 
assign mab = ~MAB;  //complement 
assign haf = ~HAF;  //complement 
assign oef = ~OEF;  //complement 
assign FFC = ~ffc;  //complement 
assign FFK = ~ffk;  //complement 
assign NAB = ~nab;  //complement 
assign hag = ~HAG;  //complement 
assign oeg = ~OEG;  //complement 
assign fec = ~FEC;  //complement 
assign fek = ~FEK;  //complement 
assign gab =  feb & fea  |  feb & ffb  ; 
assign GAB = ~gab; //complement 
assign hah = ~HAH;  //complement 
assign oeh = ~OEH;  //complement 
assign BAM =  AAM & acm & aem  |  aam & ACM & aem  |  aam & acm & AEM  |  AAM & ACM & AEM  ; 
assign bam = ~BAM; //complement 
assign bcn =  AAM & acm & aem  |  aam & ACM & aem  |  aam & acm & AEM  |  aam & acm & aem  ; 
assign BCN = ~bcn;  //complement 
assign aam = ~AAM;  //complement 
assign aan = ~AAN;  //complement 
assign agm = ~AGM;  //complement 
assign agn = ~AGN;  //complement 
assign AIM = ~aim;  //complement 
assign AIN = ~ain;  //complement 
assign BAN =  AAN & acn & aen  |  aan & ACN & aen  |  aan & acn & AEN  |  AAN & ACN & AEN  ; 
assign ban = ~BAN; //complement 
assign bco =  AAN & acn & aen  |  aan & ACN & aen  |  aan & acn & AEN  |  aan & acn & aen  ; 
assign BCO = ~bco;  //complement 
assign acm = ~ACM;  //complement 
assign acn = ~ACN;  //complement 
assign aem = ~AEM;  //complement 
assign aen = ~AEN;  //complement 
assign AKM = ~akm;  //complement 
assign AKN = ~akn;  //complement 
assign BAO =  AAO & aco & aeo  |  aao & ACO & aeo  |  aao & aco & AEO  |  AAO & ACO & AEO  ; 
assign bao = ~BAO; //complement 
assign bcp =  AAO & aco & aeo  |  aao & ACO & aeo  |  aao & aco & AEO  |  aao & aco & aeo  ; 
assign BCP = ~bcp;  //complement 
assign aao = ~AAO;  //complement 
assign aap = ~AAP;  //complement 
assign ago = ~AGO;  //complement 
assign agp = ~AGP;  //complement 
assign AIO = ~aio;  //complement 
assign AIP = ~aip;  //complement 
assign BAP =  AAP & acp & aep  |  aap & ACP & aep  |  aap & acp & AEP  |  AAP & ACP & AEP  ; 
assign bap = ~BAP; //complement 
assign bda =  AAP & acp & aep  |  aap & ACP & aep  |  aap & acp & AEP  |  aap & acp & aep  ; 
assign BDA = ~bda;  //complement 
assign aco = ~ACO;  //complement 
assign acp = ~ACP;  //complement 
assign aeo = ~AEO;  //complement 
assign aep = ~AEP;  //complement 
assign AKO = ~ako;  //complement 
assign AKP = ~akp;  //complement 
assign qrb = ~QRB;  //complement 
assign oib = ~OIB;  //complement 
assign qra = ~QRA;  //complement 
assign obn = ~OBN;  //complement 
assign wbn = ~WBN;  //complement 
assign oif = ~OIF;  //complement 
assign olb = ~OLB;  //complement 
assign qcb = ~QCB;  //complement 
assign TJB =  QBF & qmf & qdb & wbk & wbl  ; 
assign tjb = ~TJB;  //complement  
assign KCB =  QBF & qmf & qdb  ; 
assign kcb = ~KCB;  //complement 
assign obg = ~OBG;  //complement 
assign wbg = ~WBG;  //complement 
assign obh = ~OBH;  //complement 
assign wbh = ~WBH;  //complement 
assign QDB = ~qdb;  //complement 
assign QDF = ~qdf;  //complement 
assign KBF =  QBF & qmf  ; 
assign kbf = ~KBF;  //complement 
assign TJF =  QTB & qdb  ; 
assign tjf = ~TJF;  //complement 
assign obi = ~OBI;  //complement 
assign wbi = ~WBI;  //complement 
assign obj = ~OBJ;  //complement 
assign wbj = ~WBJ;  //complement 
assign OFB = ~ofb;  //complement 
assign qfb = ~QFB;  //complement 
assign obk = ~OBK;  //complement 
assign wbk = ~WBK;  //complement 
assign obl = ~OBL;  //complement 
assign wbl = ~WBL;  //complement 
assign ldi =  cfa & cha  |  cfb & chb  ; 
assign LDI = ~ldi;  //complement 
assign ldj =  cfc & chc  |  cfd & chd  ; 
assign LDJ = ~ldj;  //complement 
assign SAK = ~sak;  //complement 
assign SBK = ~sbk;  //complement 
assign SCK = ~sck;  //complement 
assign SDK = ~sdk;  //complement 
assign LCI =  CFA & CHA & CFB  |  CFA & CHA & CHB  |  CFB & CHB  ; 
assign lci = ~LCI; //complement 
assign fcl = ~FCL;  //complement 
assign fdl = ~FDL;  //complement 
assign JDJ =  DAP  ; 
assign jdj = ~JDJ;  //complement 
assign JDK =  EDA & DAP  |  DBA  ; 
assign jdk = ~JDK;  //complement 
assign DBA = ~dba;  //complement 
assign DBB = ~dbb;  //complement 
assign SIK = ~sik;  //complement 
assign SIL = ~sil;  //complement 
assign SJL = ~sjl;  //complement 
assign JDL =  DAP & EDA & EDB  |  DBA & EDB  |  DBB  ; 
assign jdl = ~JDL;  //complement 
assign DBC = ~dbc;  //complement 
assign DBD = ~dbd;  //complement 
assign LCJ =  CFC & CHC & CFD  |  CFC & CHC & CHD  |  CFD & CHD  ; 
assign lcj = ~LCJ; //complement 
assign jej =  dap & eap & eap  ; 
assign JEJ = ~jej;  //complement 
assign jek =  dba & dap & eap  |  dba & eda  ; 
assign JEK = ~jek;  //complement 
assign jel =  eap & dap & dba & dbb  |  eda & dba & dbb  |  edb & dbb  ; 
assign JEL = ~jel;  //complement 
assign SAI = ~sai;  //complement 
assign SBI = ~sbi;  //complement 
assign SCI = ~sci;  //complement 
assign SDI = ~sdi;  //complement 
assign SEI = ~sei;  //complement 
assign SFI = ~sfi;  //complement 
assign SGI = ~sgi;  //complement 
assign SHI = ~shi;  //complement 
assign SII = ~sii;  //complement 
assign SJI = ~sji;  //complement 
assign fci = ~FCI;  //complement 
assign fdi = ~FDI;  //complement 
assign SAJ = ~saj;  //complement 
assign SBJ = ~sbj;  //complement 
assign SCJ = ~scj;  //complement 
assign SDJ = ~sdj;  //complement 
assign SEJ = ~sej;  //complement 
assign SFJ = ~sfj;  //complement 
assign SGJ = ~sgj;  //complement 
assign SHJ = ~shj;  //complement 
assign SIJ = ~sij;  //complement 
assign SJJ = ~sjj;  //complement 
assign fcj = ~FCJ;  //complement 
assign fdj = ~FDJ;  //complement 
assign FFD = ~ffd;  //complement 
assign FFL = ~ffl;  //complement 
assign SEK = ~sek;  //complement 
assign SFK = ~sfk;  //complement 
assign SGK = ~sgk;  //complement 
assign SHK = ~shk;  //complement 
assign SJK = ~sjk;  //complement 
assign fck = ~FCK;  //complement 
assign fdk = ~FDK;  //complement 
assign SAL = ~sal;  //complement 
assign SBL = ~sbl;  //complement 
assign SCL = ~scl;  //complement 
assign SDL = ~sdl;  //complement 
assign SEL = ~sel;  //complement 
assign SFL = ~sfl;  //complement 
assign SGL = ~sgl;  //complement 
assign SHL = ~shl;  //complement 
assign GAC =  FEA & FFB & FFC  |  FEB & FFC  |  FEC  ; 
assign gac = ~GAC;  //complement 
assign oel = ~OEL;  //complement 
assign eda = ~EDA;  //complement 
assign cfa = ~CFA;  //complement 
assign CHB = ~chb;  //complement 
assign cba = ~CBA;  //complement 
assign CDB = ~cdb;  //complement 
assign edb = ~EDB;  //complement 
assign cfb = ~CFB;  //complement 
assign CHC = ~chc;  //complement 
assign cbb = ~CBB;  //complement 
assign CDC = ~cdc;  //complement 
assign edc = ~EDC;  //complement 
assign cfc = ~CFC;  //complement 
assign CHD = ~chd;  //complement 
assign cbc = ~CBC;  //complement 
assign CDD = ~cdd;  //complement 
assign edd = ~EDD;  //complement 
assign bfe =  ABD & add & afd  |  abd & ADD & afd  |  abd & add & AFD  |  abd & add & afd  ; 
assign BFE = ~bfe;  //complement 
assign cfd = ~CFD;  //complement 
assign CHE = ~che;  //complement 
assign cbd = ~CBD;  //complement 
assign CDE = ~cde;  //complement 
assign lbi =  cba & cda  |  cbb & cdb  ; 
assign LBI = ~lbi;  //complement 
assign lbj =  cbc & cdc  |  cbd & cdd  ; 
assign LBJ = ~lbj;  //complement 
assign LAJ =  CBC & CDC & CBD  |  CBC & CDC & CDD  |  CBD & CDD  ; 
assign laj = ~LAJ; //complement 
assign LAI =  CBA & CDA & CBB  |  CBA & CDA & CDB  |  CBB & CDB  ; 
assign lai = ~LAI; //complement 
assign hai = ~HAI;  //complement 
assign oei = ~OEI;  //complement 
assign mbc = ~MBC;  //complement 
assign mac = ~MAC;  //complement 
assign haj = ~HAJ;  //complement 
assign oej = ~OEJ;  //complement 
assign hak = ~HAK;  //complement 
assign oek = ~OEK;  //complement 
assign fed = ~FED;  //complement 
assign fel = ~FEL;  //complement 
assign hal = ~HAL;  //complement 
assign BBA =  ABA & ada & afa  |  aba & ADA & afa  |  aba & ada & AFA  |  ABA & ADA & AFA  ; 
assign bba = ~BBA; //complement 
assign bdb =  ABA & ada & afa  |  aba & ADA & afa  |  aba & ada & AFA  |  aba & ada & afa  ; 
assign BDB = ~bdb;  //complement 
assign aba = ~ABA;  //complement 
assign abb = ~ABB;  //complement 
assign aha = ~AHA;  //complement 
assign ahb = ~AHB;  //complement 
assign AJA = ~aja;  //complement 
assign AJB = ~ajb;  //complement 
assign BBB =  ABB & adb & afb  |  abb & ADB & afb  |  abb & adb & AFB  |  ABB & ADB & AFB  ; 
assign bbb = ~BBB; //complement 
assign bdc =  ABB & adb & afb  |  abb & ADB & afb  |  abb & adb & AFB  |  abb & adb & afb  ; 
assign BDC = ~bdc;  //complement 
assign ada = ~ADA;  //complement 
assign adb = ~ADB;  //complement 
assign afa = ~AFA;  //complement 
assign afb = ~AFB;  //complement 
assign ALA = ~ala;  //complement 
assign ALB = ~alb;  //complement 
assign BBC =  ABC & adc & afc  |  abc & ADC & afc  |  abc & adc & AFC  |  ABC & ADC & AFC  ; 
assign bbc = ~BBC; //complement 
assign bdd =  ABC & adc & afc  |  abc & ADC & afc  |  abc & adc & AFC  |  abc & adc & afc  ; 
assign BDD = ~bdd;  //complement 
assign abc = ~ABC;  //complement 
assign abd = ~ABD;  //complement 
assign ahc = ~AHC;  //complement 
assign ahd = ~AHD;  //complement 
assign AJC = ~ajc;  //complement 
assign AJD = ~ajd;  //complement 
assign BBD =  ABD & add & afd  |  abd & ADD & afd  |  abd & add & AFD  |  ABD & ADD & AFD  ; 
assign bbd = ~BBD; //complement 
assign bde =  ABD & add & afd  |  abd & ADD & afd  |  abd & add & AFD  |  abd & add & afd  ; 
assign BDE = ~bde;  //complement 
assign adc = ~ADC;  //complement 
assign add = ~ADD;  //complement 
assign afc = ~AFC;  //complement 
assign afd = ~AFD;  //complement 
assign ALC = ~alc;  //complement 
assign ALD = ~ald;  //complement 
assign tda = ~TDA;  //complement 
assign tdb = ~TDB;  //complement 
assign tdc = ~TDC;  //complement 
assign tdd = ~TDD;  //complement 
assign tde = ~TDE;  //complement 
assign tdf = ~TDF;  //complement 
assign ocm = ~OCM;  //complement 
assign wcm = ~WCM;  //complement 
assign qmc = ~QMC;  //complement 
assign qmg = ~QMG;  //complement 
assign TKA =  QBC & qmc & qdg & wck & wcl  ; 
assign tka = ~TKA;  //complement  
assign oca = ~OCA;  //complement 
assign wca = ~WCA;  //complement 
assign ocb = ~OCB;  //complement 
assign wcb = ~WCB;  //complement 
assign qbc = ~QBC;  //complement 
assign qbg = ~QBG;  //complement 
assign KBC =  QBC & qmc & QDC  ; 
assign kbc = ~KBC;  //complement 
assign TKE =  QTC & qdg  ; 
assign tke = ~TKE;  //complement 
assign occ = ~OCC;  //complement 
assign wcc = ~WCC;  //complement 
assign ocd = ~OCD;  //complement 
assign wcd = ~WCD;  //complement 
assign qgc = ~QGC;  //complement 
assign tkc = ~TKC;  //complement 
assign tkd = ~TKD;  //complement 
assign QTC = ~qtc;  //complement 
assign OHC = ~ohc;  //complement 
assign oce = ~OCE;  //complement 
assign wce = ~WCE;  //complement 
assign ocf = ~OCF;  //complement 
assign wcf = ~WCF;  //complement 
assign LCK =  CFE & CHE & CFF  |  CFE & CHE & CHF  |  CFF & CHF  ; 
assign lck = ~LCK; //complement 
assign JDN =  DBD  ; 
assign jdn = ~JDN;  //complement 
assign JDO =  EDE & DBD  |  DBE  ; 
assign jdo = ~JDO;  //complement 
assign DBE = ~dbe;  //complement 
assign DBF = ~dbf;  //complement 
assign ldk =  cfe & che  |  cff & chf  ; 
assign LDK = ~ldk;  //complement 
assign ldl =  cfg & chg  |  cfh & chh  ; 
assign LDL = ~ldl;  //complement 
assign JDP =  DBD & EDE & EDF  |  DBE & EDF  |  DBF  ; 
assign jdp = ~JDP;  //complement 
assign DBG = ~dbg;  //complement 
assign DBH = ~dbh;  //complement 
assign LCL =  CFG & CHG & CFH  |  CFG & CHG & CHH  |  CFH & CHH  ; 
assign lcl = ~LCL; //complement 
assign jen =  dbd & edd & edd  ; 
assign JEN = ~jen;  //complement 
assign jeo =  dbe & dbd & edd  |  dbe & ede  ; 
assign JEO = ~jeo;  //complement 
assign jep =  edd & dbd & dbe & dbf  |  ede & dbe & dbf  |  edf & dbf  ; 
assign JEP = ~jep;  //complement 
assign SAM = ~sam;  //complement 
assign SBM = ~sbm;  //complement 
assign SCM = ~scm;  //complement 
assign SDM = ~sdm;  //complement 
assign SEM = ~sem;  //complement 
assign SFM = ~sfm;  //complement 
assign SGM = ~sgm;  //complement 
assign SHM = ~shm;  //complement 
assign SIM = ~sim;  //complement 
assign SJM = ~sjm;  //complement 
assign fcm = ~FCM;  //complement 
assign fdm = ~FDM;  //complement 
assign SAN = ~san;  //complement 
assign SBN = ~sbn;  //complement 
assign SCN = ~scn;  //complement 
assign SDN = ~sdn;  //complement 
assign SEN = ~sen;  //complement 
assign SFN = ~sfn;  //complement 
assign SGN = ~sgn;  //complement 
assign SHN = ~shn;  //complement 
assign SIN = ~sin;  //complement 
assign SJN = ~sjn;  //complement 
assign fcn = ~FCN;  //complement 
assign fdn = ~FDN;  //complement 
assign SAO = ~sao;  //complement 
assign SBO = ~sbo;  //complement 
assign SCO = ~sco;  //complement 
assign SDO = ~sdo;  //complement 
assign SEO = ~seo;  //complement 
assign SFO = ~sfo;  //complement 
assign SGO = ~sgo;  //complement 
assign SHO = ~sho;  //complement 
assign SJO = ~sjo;  //complement 
assign SIO = ~sio;  //complement 
assign fco = ~FCO;  //complement 
assign fdo = ~FDO;  //complement 
assign SAP = ~sap;  //complement 
assign SBP = ~sbp;  //complement 
assign SCP = ~scp;  //complement 
assign SDP = ~sdp;  //complement 
assign SEP = ~sep;  //complement 
assign SFP = ~sfp;  //complement 
assign SGP = ~sgp;  //complement 
assign SHP = ~shp;  //complement 
assign SIP = ~sip;  //complement 
assign SJP = ~sjp;  //complement 
assign fcp = ~FCP;  //complement 
assign fdp = ~FDP;  //complement 
assign ede = ~EDE;  //complement 
assign cfe = ~CFE;  //complement 
assign CHF = ~chf;  //complement 
assign cbe = ~CBE;  //complement 
assign CDF = ~cdf;  //complement 
assign edf = ~EDF;  //complement 
assign cff = ~CFF;  //complement 
assign CHG = ~chg;  //complement 
assign cbf = ~CBF;  //complement 
assign CDG = ~cdg;  //complement 
assign edg = ~EDG;  //complement 
assign cfg = ~CFG;  //complement 
assign CHH = ~chh;  //complement 
assign cbg = ~CBG;  //complement 
assign CDH = ~cdh;  //complement 
assign edh = ~EDH;  //complement 
assign bfi =  ABH & adh & afh  |  abh & ADH & afh  |  abh & adh & AFH  |  abh & adh & afh  ; 
assign BFI = ~bfi;  //complement 
assign cfh = ~CFH;  //complement 
assign CHI = ~chi;  //complement 
assign cbh = ~CBH;  //complement 
assign CDI = ~cdi;  //complement 
assign lbk =  cbe & cde  |  cbf & cdf  ; 
assign LBK = ~lbk;  //complement 
assign lbl =  cbg & cdg  |  cbh & cdh  ; 
assign LBL = ~lbl;  //complement 
assign LAL =  CBG & CDG & CBH  |  CBG & CDG & CDH  |  CBH & CDH  ; 
assign lal = ~LAL; //complement 
assign LAK =  CBE & CDE & CBF  |  CBE & CDE & CDF  |  CBF & CDF  ; 
assign lak = ~LAK; //complement 
assign ham = ~HAM;  //complement 
assign oem = ~OEM;  //complement 
assign NBB = ~nbb;  //complement 
assign NAC = ~nac;  //complement 
assign han = ~HAN;  //complement 
assign oen = ~OEN;  //complement 
assign FFE = ~ffe;  //complement 
assign FFM = ~ffm;  //complement 
assign hao = ~HAO;  //complement 
assign oeo = ~OEO;  //complement 
assign fee = ~FEE;  //complement 
assign GAD =  FEA & FFB & FFC & FFD  |  FEB & FFC & FFD  |  FEC & FFD  |  FED  ; 
assign gad = ~GAD;  //complement 
assign hap = ~HAP;  //complement 
assign oep = ~OEP;  //complement 
assign BBE =  ABE & ade & afe  |  abe & ADE & afe  |  abe & ade & AFE  |  ABE & ADE & AFE  ; 
assign bbe = ~BBE; //complement 
assign bdf =  ABE & ade & afe  |  abe & ADE & afe  |  abe & ade & AFE  |  abe & ade & afe  ; 
assign BDF = ~bdf;  //complement 
assign abe = ~ABE;  //complement 
assign abf = ~ABF;  //complement 
assign ahe = ~AHE;  //complement 
assign ahf = ~AHF;  //complement 
assign AJE = ~aje;  //complement 
assign AJF = ~ajf;  //complement 
assign BBF =  ABF & adf & aff  |  abf & ADF & aff  |  abf & adf & AFF  |  ABF & ADF & AFF  ; 
assign bbf = ~BBF; //complement 
assign bdg =  ABF & adf & aff  |  abf & ADF & aff  |  abf & adf & AFF  |  abf & adf & aff  ; 
assign BDG = ~bdg;  //complement 
assign ade = ~ADE;  //complement 
assign adf = ~ADF;  //complement 
assign afe = ~AFE;  //complement 
assign aff = ~AFF;  //complement 
assign ALE = ~ale;  //complement 
assign ALF = ~alf;  //complement 
assign BBG =  ABG & adg & afg  |  abg & ADG & afg  |  abg & adg & AFG  |  ABG & ADG & AFG  ; 
assign bbg = ~BBG; //complement 
assign bdh =  ABG & adg & afg  |  abg & ADG & afg  |  abg & adg & AFG  |  abg & adg & afg  ; 
assign BDH = ~bdh;  //complement 
assign abg = ~ABG;  //complement 
assign abh = ~ABH;  //complement 
assign ahg = ~AHG;  //complement 
assign ahh = ~AHH;  //complement 
assign AJG = ~ajg;  //complement 
assign AJH = ~ajh;  //complement 
assign BBH =  ABH & adh & afh  |  abh & ADH & afh  |  abh & adh & AFH  |  ABH & ADH & AFH  ; 
assign bbh = ~BBH; //complement 
assign bdi =  ABH & adh & afh  |  abh & ADH & afh  |  abh & adh & AFH  |  abh & adh & afh  ; 
assign BDI = ~bdi;  //complement 
assign adg = ~ADG;  //complement 
assign adh = ~ADH;  //complement 
assign afg = ~AFG;  //complement 
assign afh = ~AFH;  //complement 
assign ALG = ~alg;  //complement 
assign ALH = ~alh;  //complement 
assign tca = ~TCA;  //complement 
assign tcb = ~TCB;  //complement 
assign tcg = ~TCG;  //complement 
assign tcc = ~TCC;  //complement 
assign tcd = ~TCD;  //complement 
assign oic = ~OIC;  //complement 
assign tce = ~TCE;  //complement 
assign tcf = ~TCF;  //complement 
assign ocn = ~OCN;  //complement 
assign wcn = ~WCN;  //complement 
assign oig = ~OIG;  //complement 
assign olc = ~OLC;  //complement 
assign qcc = ~QCC;  //complement 
assign TKB =  QBG & qmg & qdc & wck & wcl  ; 
assign tkb = ~TKB;  //complement  
assign KCC =  QBG & qmg & qdc  ; 
assign kcc = ~KCC;  //complement 
assign ocg = ~OCG;  //complement 
assign wcg = ~WCG;  //complement 
assign och = ~OCH;  //complement 
assign wch = ~WCH;  //complement 
assign QDC = ~qdc;  //complement 
assign QDG = ~qdg;  //complement 
assign KBG =  QBG & qmg  ; 
assign kbg = ~KBG;  //complement 
assign TKF =  QTC & qdc  ; 
assign tkf = ~TKF;  //complement 
assign oci = ~OCI;  //complement 
assign wci = ~WCI;  //complement 
assign ocj = ~OCJ;  //complement 
assign wcj = ~WCJ;  //complement 
assign OFC = ~ofc;  //complement 
assign qfc = ~QFC;  //complement 
assign ock = ~OCK;  //complement 
assign wck = ~WCK;  //complement 
assign ocl = ~OCL;  //complement 
assign wcl = ~WCL;  //complement 
assign LCM =  CFI & CHI & CFJ  |  CFI & CHI & CHJ  |  CFJ & CHJ  ; 
assign lcm = ~LCM; //complement 
assign JDR =  DBH  ; 
assign jdr = ~JDR;  //complement 
assign JDS =  EDI & DBH  |  DBI  ; 
assign jds = ~JDS;  //complement 
assign DBI = ~dbi;  //complement 
assign DBJ = ~dbj;  //complement 
assign ldm =  cfi & chi  |  cfj & chj  ; 
assign LDM = ~ldm;  //complement 
assign ldn =  cfk & chk  |  cfl & chl  ; 
assign LDN = ~ldn;  //complement 
assign JDT =  DBH & EDI & EDJ  |  DBI & EDJ  |  DBJ  ; 
assign jdt = ~JDT;  //complement 
assign DBK = ~dbk;  //complement 
assign DBL = ~dbl;  //complement 
assign LCN =  CFK & CHK & CFL  |  CFK & CHK & CHL  |  CFL & CHL  ; 
assign lcn = ~LCN; //complement 
assign jer =  dbh & edh & edh  ; 
assign JER = ~jer;  //complement 
assign jes =  dbi & dbh & edh  |  dbi & edi  ; 
assign JES = ~jes;  //complement 
assign jet =  edh & dbh & dbi & dbj  |  edi & dbi & dbj  |  edj & dbj  ; 
assign JET = ~jet;  //complement 
assign SAQ = ~saq;  //complement 
assign SBQ = ~sbq;  //complement 
assign SCQ = ~scq;  //complement 
assign SDQ = ~sdq;  //complement 
assign SEQ = ~seq;  //complement 
assign SFQ = ~sfq;  //complement 
assign SGQ = ~sgq;  //complement 
assign SHQ = ~shq;  //complement 
assign SIQ = ~siq;  //complement 
assign SJQ = ~sjq;  //complement 
assign fcq = ~FCQ;  //complement 
assign fdq = ~FDQ;  //complement 
assign SAR = ~sar;  //complement 
assign SBR = ~sbr;  //complement 
assign SCR = ~scr;  //complement 
assign SDR = ~sdr;  //complement 
assign SER = ~ser;  //complement 
assign SFR = ~sfr;  //complement 
assign SGR = ~sgr;  //complement 
assign SHR = ~shr;  //complement 
assign SIR = ~sir;  //complement 
assign SJR = ~sjr;  //complement 
assign fcr = ~FCR;  //complement 
assign fdr = ~FDR;  //complement 
assign SAS = ~sas;  //complement 
assign SBS = ~sbs;  //complement 
assign SCS = ~scs;  //complement 
assign SDS = ~sds;  //complement 
assign SES = ~ses;  //complement 
assign SFS = ~sfs;  //complement 
assign SGS = ~sgs;  //complement 
assign SHS = ~shs;  //complement 
assign SIS = ~sis;  //complement 
assign SJS = ~sjs;  //complement 
assign fcs = ~FCS;  //complement 
assign fds = ~FDS;  //complement 
assign SAT = ~sat;  //complement 
assign SBT = ~sbt;  //complement 
assign SCT = ~sct;  //complement 
assign SDT = ~sdt;  //complement 
assign SET = ~set;  //complement 
assign SFT = ~sft;  //complement 
assign SGT = ~sgt;  //complement 
assign SHT = ~sht;  //complement 
assign SIT = ~sit;  //complement 
assign SJT = ~sjt;  //complement 
assign fct = ~FCT;  //complement 
assign fdt = ~FDT;  //complement 
assign edi = ~EDI;  //complement 
assign cfi = ~CFI;  //complement 
assign CHJ = ~chj;  //complement 
assign cbi = ~CBI;  //complement 
assign CDJ = ~cdj;  //complement 
assign edj = ~EDJ;  //complement 
assign cfj = ~CFJ;  //complement 
assign CHK = ~chk;  //complement 
assign cbj = ~CBJ;  //complement 
assign CDK = ~cdk;  //complement 
assign edk = ~EDK;  //complement 
assign cfk = ~CFK;  //complement 
assign CHL = ~chl;  //complement 
assign cbk = ~CBK;  //complement 
assign CDL = ~cdl;  //complement 
assign edl = ~EDL;  //complement 
assign bfm =  ABL & adl & afl  |  abl & ADL & afl  |  abl & adl & AFL  |  abl & adl & afl  ; 
assign BFM = ~bfm;  //complement 
assign cfl = ~CFL;  //complement 
assign CHM = ~chm;  //complement 
assign cbl = ~CBL;  //complement 
assign CDM = ~cdm;  //complement 
assign lbm =  cbi & cdi  |  cbj & cdj  ; 
assign LBM = ~lbm;  //complement 
assign lbn =  cbk & cdk  |  cbl & cdl  ; 
assign LBN = ~lbn;  //complement 
assign LAN =  CBK & CDK & CBL  |  CBK & CDK & CDL  |  CBL & CDL  ; 
assign lan = ~LAN; //complement 
assign LAM =  CBI & CDI & CBJ  |  CBI & CDI & CDJ  |  CBJ & CDJ  ; 
assign lam = ~LAM; //complement 
assign haq = ~HAQ;  //complement 
assign oeq = ~OEQ;  //complement 
assign NBC = ~nbc;  //complement 
assign mad = ~MAD;  //complement 
assign har = ~HAR;  //complement 
assign oer = ~OER;  //complement 
assign FFF = ~fff;  //complement 
assign NAD = ~nad;  //complement 
assign has = ~HAS;  //complement 
assign oes = ~OES;  //complement 
assign fef = ~FEF;  //complement 
assign GAE =  FEI & FFJ & FFK & FFL & FFM  |  FEJ & FFK & FFL & FFM  |  FEK & FFL & FFM  |  FEL & FFM  |  FEE  ; 
assign gae = ~GAE;  //complement 
assign hat = ~HAT;  //complement 
assign oet = ~OET;  //complement 
assign BBI =  ABI & adi & afi  |  abi & ADI & afi  |  abi & adi & AFI  |  ABI & ADI & AFI  ; 
assign bbi = ~BBI; //complement 
assign bdj =  ABI & adi & afi  |  abi & ADI & afi  |  abi & adi & AFI  |  abi & adi & afi  ; 
assign BDJ = ~bdj;  //complement 
assign abi = ~ABI;  //complement 
assign abj = ~ABJ;  //complement 
assign ahi = ~AHI;  //complement 
assign ahj = ~AHJ;  //complement 
assign AJI = ~aji;  //complement 
assign AJJ = ~ajj;  //complement 
assign BBJ =  ABJ & adj & afj  |  abj & ADJ & afj  |  abj & adj & AFJ  |  ABJ & ADJ & AFJ  ; 
assign bbj = ~BBJ; //complement 
assign bdk =  ABJ & adj & afj  |  abj & ADJ & afj  |  abj & adj & AFJ  |  abj & adj & afj  ; 
assign BDK = ~bdk;  //complement 
assign adi = ~ADI;  //complement 
assign adj = ~ADJ;  //complement 
assign afi = ~AFI;  //complement 
assign afj = ~AFJ;  //complement 
assign ALI = ~ali;  //complement 
assign ALJ = ~alj;  //complement 
assign BBK =  ABK & adk & afk  |  abk & ADK & afk  |  abk & adk & AFK  |  ABK & ADK & AFK  ; 
assign bbk = ~BBK; //complement 
assign bdl =  ABK & adk & afk  |  abk & ADK & afk  |  abk & adk & AFK  |  abk & adk & afk  ; 
assign BDL = ~bdl;  //complement 
assign abk = ~ABK;  //complement 
assign abl = ~ABL;  //complement 
assign ahk = ~AHK;  //complement 
assign ahl = ~AHL;  //complement 
assign AJK = ~ajk;  //complement 
assign AJL = ~ajl;  //complement 
assign adk = ~ADK;  //complement 
assign adl = ~ADL;  //complement 
assign BBL =  ABL & adl & afl  |  abl & ADL & afl  |  abl & adl & AFL  |  ABL & ADL & AFL  ; 
assign bbl = ~BBL; //complement 
assign bdm =  ABL & adl & afl  |  abl & ADL & afl  |  abl & adl & AFL  |  abl & adl & afl  ; 
assign BDM = ~bdm;  //complement 
assign afk = ~AFK;  //complement 
assign afl = ~AFL;  //complement 
assign ALK = ~alk;  //complement 
assign ALL = ~all;  //complement 
assign tea = ~TEA;  //complement 
assign teb = ~TEB;  //complement 
assign tfa = ~TFA;  //complement 
assign tfb = ~TFB;  //complement 
assign odm = ~ODM;  //complement 
assign wdm = ~WDM;  //complement 
assign qmd = ~QMD;  //complement 
assign qmh = ~QMH;  //complement 
assign TLA =  QBD & qmd & qdh & wdk & wdl  ; 
assign tla = ~TLA;  //complement  
assign oda = ~ODA;  //complement 
assign wda = ~WDA;  //complement 
assign odb = ~ODB;  //complement 
assign wdb = ~WDB;  //complement 
assign qbd = ~QBD;  //complement 
assign qbh = ~QBH;  //complement 
assign KBD =  QBD & qmd & QDD  ; 
assign kbd = ~KBD;  //complement 
assign TLE =  QTD & qdh  ; 
assign tle = ~TLE;  //complement 
assign odc = ~ODC;  //complement 
assign wdc = ~WDC;  //complement 
assign odd = ~ODD;  //complement 
assign wdd = ~WDD;  //complement 
assign qgd = ~QGD;  //complement 
assign tlc = ~TLC;  //complement 
assign tld = ~TLD;  //complement 
assign QTD = ~qtd;  //complement 
assign OHD = ~ohd;  //complement 
assign ode = ~ODE;  //complement 
assign wde = ~WDE;  //complement 
assign odf = ~ODF;  //complement 
assign wdf = ~WDF;  //complement 
assign LCO =  CFM & CHM & CFN  |  CFM & CHM & CHN  |  CFN & CHN  ; 
assign lco = ~LCO; //complement 
assign DBM = ~dbm;  //complement 
assign DBN = ~dbn;  //complement 
assign SIW = ~siw;  //complement 
assign ldo =  cfm & chm  |  cfn & chn  ; 
assign LDO = ~ldo;  //complement 
assign ldp =  cfo & cho  |  cfp & chp  ; 
assign LDP = ~ldp;  //complement 
assign DBO = ~dbo;  //complement 
assign DBP = ~dbp;  //complement 
assign LCP =  CFO & CHO & CFP  |  CFO & CHO & CHP  |  CFP & CHP  ; 
assign lcp = ~LCP; //complement 
assign JDV =  DBL  ; 
assign jdv = ~JDV;  //complement 
assign jev =  dbl & edl  ; 
assign JEV = ~jev;  //complement 
assign SAU = ~sau;  //complement 
assign SBU = ~sbu;  //complement 
assign SCU = ~scu;  //complement 
assign SDU = ~sdu;  //complement 
assign SEU = ~seu;  //complement 
assign SFU = ~sfu;  //complement 
assign SGU = ~sgu;  //complement 
assign SHU = ~shu;  //complement 
assign SIU = ~siu;  //complement 
assign SJU = ~sju;  //complement 
assign fcu = ~FCU;  //complement 
assign fdu = ~FDU;  //complement 
assign SAV = ~sav;  //complement 
assign SBV = ~sbv;  //complement 
assign SCV = ~scv;  //complement 
assign SDV = ~sdv;  //complement 
assign SEV = ~sev;  //complement 
assign SFV = ~sfv;  //complement 
assign SGV = ~sgv;  //complement 
assign SHV = ~shv;  //complement 
assign SIV = ~siv;  //complement 
assign SJV = ~sjv;  //complement 
assign fcv = ~FCV;  //complement 
assign fdv = ~FDV;  //complement 
assign SBW = ~sbw;  //complement 
assign SCW = ~scw;  //complement 
assign SDW = ~sdw;  //complement 
assign SAW = ~saw;  //complement 
assign SEW = ~sew;  //complement 
assign SFW = ~sfw;  //complement 
assign SGW = ~sgw;  //complement 
assign SHW = ~shw;  //complement 
assign SJW = ~sjw;  //complement 
assign SAX = ~sax;  //complement 
assign SBX = ~sbx;  //complement 
assign SCX = ~scx;  //complement 
assign SDX = ~sdx;  //complement 
assign SEX = ~sex;  //complement 
assign SFX = ~sfx;  //complement 
assign SGX = ~sgx;  //complement 
assign SHX = ~shx;  //complement 
assign SIX = ~six;  //complement 
assign SJX = ~sjx;  //complement 
assign edm = ~EDM;  //complement 
assign cfm = ~CFM;  //complement 
assign CHN = ~chn;  //complement 
assign cbm = ~CBM;  //complement 
assign CDN = ~cdn;  //complement 
assign edn = ~EDN;  //complement 
assign cfn = ~CFN;  //complement 
assign CHO = ~cho;  //complement 
assign cbn = ~CBN;  //complement 
assign CDO = ~cdo;  //complement 
assign edo = ~EDO;  //complement 
assign cfo = ~CFO;  //complement 
assign CHP = ~chp;  //complement 
assign cbo = ~CBO;  //complement 
assign CDP = ~cdp;  //complement 
assign edp = ~EDP;  //complement 
assign cfp = ~CFP;  //complement 
assign cbp = ~CBP;  //complement 
assign lbo =  cbm & cdm  |  cbn & cdn  ; 
assign LBO = ~lbo;  //complement 
assign lbp =  cbo & cdo  |  cbp & cdp  ; 
assign LBP = ~lbp;  //complement 
assign LAP =  CBO & CDO & CBP  |  CBO & CDO & CDP  |  CBP & CDP  ; 
assign lap = ~LAP; //complement 
assign LAO =  CBM & CDM & CBN  |  CBM & CDM & CDN  |  CBN & CDN  ; 
assign lao = ~LAO; //complement 
assign hau = ~HAU;  //complement 
assign oeu = ~OEU;  //complement 
assign mbd = ~MBD;  //complement 
assign XAA =  MAA & NAB & NAC & NAD & QEA  |  MAB & NAC & NAD & QEA  |  MAC & NAD & QEA  |  MAD & QEA  ; 
assign xaa = ~XAA;  //complement 
assign hav = ~HAV;  //complement 
assign oev = ~OEV;  //complement 
assign NBD = ~nbd;  //complement 
assign XAB =  MBA & NBB & NBC & NBD & QEA  |  MBB & NBC & NBD & QEA  |  MBC & NBD & QEA  |  MBD & QEA  ; 
assign xab = ~XAB;  //complement 
assign haw = ~HAW;  //complement 
assign OEX = ~oex;  //complement 
assign hax = ~HAX;  //complement 
assign GAF =  FEI & FFJ & FFK & FFL & FFM & FFF  |  FEJ & FFK & FFL & FFM & FFF  |  FEK & FFL & FFM & FFF  |  FEL & FFM & FFF  |  FFE & FFF  |  FEF  ; 
assign gaf = ~GAF;  //complement 
assign OEW = ~oew;  //complement 
assign BBM =  ABM & adm & afm  |  abm & ADM & afm  |  abm & adm & AFM  |  ABM & ADM & AFM  ; 
assign bbm = ~BBM; //complement 
assign bdn =  ABM & adm & afm  |  abm & ADM & afm  |  abm & adm & AFM  |  abm & adm & afm  ; 
assign BDN = ~bdn;  //complement 
assign abm = ~ABM;  //complement 
assign abn = ~ABN;  //complement 
assign ahm = ~AHM;  //complement 
assign ahn = ~AHN;  //complement 
assign AJM = ~ajm;  //complement 
assign AJN = ~ajn;  //complement 
assign BBN =  ABN & adn & afn  |  abn & ADN & afn  |  abn & adn & AFN  |  ABN & ADN & AFN  ; 
assign bbn = ~BBN; //complement 
assign bdo =  ABN & adn & afn  |  abn & ADN & afn  |  abn & adn & AFN  |  abn & adn & afn  ; 
assign BDO = ~bdo;  //complement 
assign adm = ~ADM;  //complement 
assign adn = ~ADN;  //complement 
assign afm = ~AFM;  //complement 
assign afn = ~AFN;  //complement 
assign ALM = ~alm;  //complement 
assign ALN = ~aln;  //complement 
assign BBO =  ABO & ado & afo  |  abo & ADO & afo  |  abo & ado & AFO  |  ABO & ADO & AFO  ; 
assign bbo = ~BBO; //complement 
assign bdp =  ABO & ado & afo  |  abo & ADO & afo  |  abo & ado & AFO  |  abo & ado & afo  ; 
assign BDP = ~bdp;  //complement 
assign abo = ~ABO;  //complement 
assign abp = ~ABP;  //complement 
assign aho = ~AHO;  //complement 
assign ahp = ~AHP;  //complement 
assign cao = ~CAO;  //complement 
assign CCP = ~ccp;  //complement 
assign BBP =  ABP & adp & afp  |  abp & ADP & afp  |  abp & adp & AFP  |  ABP & ADP & AFP  ; 
assign bbp = ~BBP; //complement 
assign ado = ~ADO;  //complement 
assign adp = ~ADP;  //complement 
assign afo = ~AFO;  //complement 
assign afp = ~AFP;  //complement 
assign ALO = ~alo;  //complement 
assign ALP = ~alp;  //complement 
assign oid = ~OID;  //complement 
assign qea = ~QEA;  //complement 
assign qec = ~QEC;  //complement 
assign OFD = ~ofd;  //complement 
assign oka = ~OKA;  //complement 
assign odn = ~ODN;  //complement 
assign wdn = ~WDN;  //complement 
assign oih = ~OIH;  //complement 
assign old = ~OLD;  //complement 
assign qcd = ~QCD;  //complement 
assign TLB =  QBH & qmh & qdd & wdk & wdl  ; 
assign tlb = ~TLB;  //complement  
assign KCD =  QBH & qmh & qdd  ; 
assign kcd = ~KCD;  //complement 
assign odg = ~ODG;  //complement 
assign wdg = ~WDG;  //complement 
assign odh = ~ODH;  //complement 
assign wdh = ~WDH;  //complement 
assign QDD = ~qdd;  //complement 
assign QDH = ~qdh;  //complement 
assign KBH =  QBH & qmh  ; 
assign kbh = ~KBH;  //complement 
assign TLF =  QTD & qdd  ; 
assign tlf = ~TLF;  //complement 
assign odi = ~ODI;  //complement 
assign wdi = ~WDI;  //complement 
assign odj = ~ODJ;  //complement 
assign wdj = ~WDJ;  //complement 
assign AJO = ~ajo;  //complement 
assign AJP = ~ajp;  //complement 
assign qfd = ~QFD;  //complement 
assign odk = ~ODK;  //complement 
assign wdk = ~WDK;  //complement 
assign odl = ~ODL;  //complement 
assign wdl = ~WDL;  //complement 
assign iaa = ~IAA; //complement 
assign iab = ~IAB; //complement 
assign iac = ~IAC; //complement 
assign iad = ~IAD; //complement 
assign iae = ~IAE; //complement 
assign iaf = ~IAF; //complement 
assign iag = ~IAG; //complement 
assign iah = ~IAH; //complement 
assign iai = ~IAI; //complement 
assign iaj = ~IAJ; //complement 
assign iak = ~IAK; //complement 
assign ial = ~IAL; //complement 
assign iam = ~IAM; //complement 
assign ian = ~IAN; //complement 
assign iao = ~IAO; //complement 
assign iap = ~IAP; //complement 
assign iba = ~IBA; //complement 
assign ibb = ~IBB; //complement 
assign ibc = ~IBC; //complement 
assign ibd = ~IBD; //complement 
assign ibe = ~IBE; //complement 
assign ibf = ~IBF; //complement 
assign ibg = ~IBG; //complement 
assign ibh = ~IBH; //complement 
assign ibi = ~IBI; //complement 
assign ibj = ~IBJ; //complement 
assign ibk = ~IBK; //complement 
assign ibl = ~IBL; //complement 
assign ibm = ~IBM; //complement 
assign ibn = ~IBN; //complement 
assign ibo = ~IBO; //complement 
assign ibp = ~IBP; //complement 
assign ica = ~ICA; //complement 
assign icb = ~ICB; //complement 
assign icc = ~ICC; //complement 
assign icd = ~ICD; //complement 
assign ice = ~ICE; //complement 
assign icf = ~ICF; //complement 
assign icg = ~ICG; //complement 
assign ich = ~ICH; //complement 
assign ici = ~ICI; //complement 
assign icj = ~ICJ; //complement 
assign ick = ~ICK; //complement 
assign icl = ~ICL; //complement 
assign icm = ~ICM; //complement 
assign icn = ~ICN; //complement 
assign ico = ~ICO; //complement 
assign icp = ~ICP; //complement 
assign ida = ~IDA; //complement 
assign idb = ~IDB; //complement 
assign idc = ~IDC; //complement 
assign idd = ~IDD; //complement 
assign ide = ~IDE; //complement 
assign idf = ~IDF; //complement 
assign idg = ~IDG; //complement 
assign idh = ~IDH; //complement 
assign idi = ~IDI; //complement 
assign idj = ~IDJ; //complement 
assign idk = ~IDK; //complement 
assign idl = ~IDL; //complement 
assign idm = ~IDM; //complement 
assign idn = ~IDN; //complement 
assign ido = ~IDO; //complement 
assign idp = ~IDP; //complement 
assign iea = ~IEA; //complement 
assign ieb = ~IEB; //complement 
assign iec = ~IEC; //complement 
assign ied = ~IED; //complement 
assign iee = ~IEE; //complement 
assign ief = ~IEF; //complement 
assign ieg = ~IEG; //complement 
assign ieh = ~IEH; //complement 
assign iei = ~IEI; //complement 
assign iej = ~IEJ; //complement 
assign iek = ~IEK; //complement 
assign iel = ~IEL; //complement 
assign iem = ~IEM; //complement 
assign ien = ~IEN; //complement 
assign ieo = ~IEO; //complement 
assign iep = ~IEP; //complement 
assign ifa = ~IFA; //complement 
assign ifb = ~IFB; //complement 
assign ifc = ~IFC; //complement 
assign ifd = ~IFD; //complement 
assign ife = ~IFE; //complement 
assign ifff  = ~IFFF ; //complement 
assign ifg = ~IFG; //complement 
assign ifh = ~IFH; //complement 
assign ifi = ~IFI; //complement 
assign ifj = ~IFJ; //complement 
assign ifk = ~IFK; //complement 
assign ifl = ~IFL; //complement 
assign ifm = ~IFM; //complement 
assign ifn = ~IFN; //complement 
assign ifo = ~IFO; //complement 
assign ifp = ~IFP; //complement 
assign iga = ~IGA; //complement 
assign igb = ~IGB; //complement 
assign igc = ~IGC; //complement 
assign igd = ~IGD; //complement 
assign ige = ~IGE; //complement 
assign igf = ~IGF; //complement 
assign igg = ~IGG; //complement 
assign igh = ~IGH; //complement 
assign igi = ~IGI; //complement 
assign igj = ~IGJ; //complement 
assign igk = ~IGK; //complement 
assign igl = ~IGL; //complement 
assign igm = ~IGM; //complement 
assign ign = ~IGN; //complement 
assign igo = ~IGO; //complement 
assign igp = ~IGP; //complement 
assign iha = ~IHA; //complement 
assign ihb = ~IHB; //complement 
assign ihc = ~IHC; //complement 
assign ihd = ~IHD; //complement 
assign ihe = ~IHE; //complement 
assign ihf = ~IHF; //complement 
assign ihg = ~IHG; //complement 
assign ihh = ~IHH; //complement 
assign ihi = ~IHI; //complement 
assign ihj = ~IHJ; //complement 
assign ihk = ~IHK; //complement 
assign ihl = ~IHL; //complement 
assign ihm = ~IHM; //complement 
assign ihn = ~IHN; //complement 
assign iho = ~IHO; //complement 
assign ihp = ~IHP; //complement 
assign iia = ~IIA; //complement 
assign iib = ~IIB; //complement 
assign iic = ~IIC; //complement 
assign iid = ~IID; //complement 
assign iie = ~IIE; //complement 
assign iif = ~IIF; //complement 
assign ija = ~IJA; //complement 
assign ijb = ~IJB; //complement 
assign ijc = ~IJC; //complement 
assign ijd = ~IJD; //complement 
assign ije = ~IJE; //complement 
assign ijf = ~IJF; //complement 
assign ijg = ~IJG; //complement 
assign ijh = ~IJH; //complement 
assign ika = ~IKA; //complement 
assign ikb = ~IKB; //complement 
assign ikc = ~IKC; //complement 
assign ikd = ~IKD; //complement 
assign ike = ~IKE; //complement 
assign ikf = ~IKF; //complement 
assign ikg = ~IKG; //complement 
assign ikh = ~IKH; //complement 
assign iki = ~IKI; //complement 
assign ikj = ~IKJ; //complement 
assign ikk = ~IKK; //complement 
assign ikm = ~IKM; //complement 
assign ikn = ~IKN; //complement 
assign iko = ~IKO; //complement 
assign ikp = ~IKP; //complement 
assign ikq = ~IKQ; //complement 
assign ikr = ~IKR; //complement 
assign iks = ~IKS; //complement 
assign ikt = ~IKT; //complement 
assign iku = ~IKU; //complement 
assign ila = ~ILA; //complement 
always@(posedge IZZ )
   begin 
 paa <= faa ; 
 pba <= paa ; 
 pca <= pba ; 
 pda <= pca ; 
 pea <= pda ; 
 pfa <= pea ; 
 pga <= pfa ; 
 pha <= pga ; 
 pia <= pha ; 
 pja <= pia ; 
 pab <= fab ; 
 pbb <= pab ; 
 pcb <= pbb ; 
 pdb <= pcb ; 
 peb <= pdb ; 
 pfb <= peb ; 
 pgb <= pfb ; 
 phb <= pgb ; 
 pib <= phb ; 
 pjb <= pib ; 
 dab <=  bab  |  bcb  |  TGA  ; 
 pac <= fac ; 
 pbc <= pac ; 
 pcc <= pbc ; 
 pdc <= pcc ; 
 pec <= pdc ; 
 pfc <= pec ; 
 pgc <= pfc ; 
 phc <= pgc ; 
 pic <= phc ; 
 pjc <= pic ; 
 dac <=  bac  |  bcc  |  TGB  ; 
 dad <=  bad  |  bcd  |  TGB  ; 
 pad <= fad ; 
 pbd <= pad ; 
 pcd <= pbd ; 
 pdd <= pcd ; 
 ped <= pdd ; 
 pfd <= ped ; 
 pgd <= pfd ; 
 phd <= pgd ; 
 pid <= phd ; 
 pjd <= pid ; 
 pae <= fae ; 
 pbe <= pae ; 
 pce <= pbe ; 
 pde <= pce ; 
 pee <= pde ; 
 pfe <= pee ; 
 pge <= pfe ; 
 phe <= pge ; 
 pie <= phe ; 
 pje <= pie ; 
 paf <= faf ; 
 pbf <= paf ; 
 pcf <= pbf ; 
 pdf <= pcf ; 
 pef <= pdf ; 
 pff <= pef ; 
 pgf <= pff ; 
 phf <= pgf ; 
 pif <= phf ; 
 pjf <= pif ; 
 par <= jfb ; 
 pbr <= par ; 
 pcr <= pbr ; 
 pdr <= pcr ; 
 pam <= qba ; 
 pbm <= pam ; 
 pcm <= pbm ; 
 pdm <= pcm ; 
 pem <= pdm ; 
 pfm <= pem ; 
 pgm <= pfm ; 
 phm <= pgm ; 
 pjm <= pim ; 
 pim <= phm ; 
 per <= pdr ; 
 pfr <= per ; 
 pgr <= pfr ; 
 phr <= pgr ; 
 pan <= qbb ; 
 pbn <= pan ; 
 pcn <= pbn ; 
 pdn <= pcn ; 
 pen <= pdn ; 
 pfn <= pen ; 
 pgn <= pfn ; 
 phn <= pgn ; 
 pin <= phn ; 
 pjn <= pin ; 
 pir <= phr ; 
 pjr <= pir ; 
 qaa <=  BAA  |  ika  ; 
 qab <=  baa  |  ika  ; 
 CEA <=  BAA & AIA  |  baa & aia  |  baa & AIA  |  BAA & aia  ;
 cgb <=  BAA & AIA  |  baa & aia  |  baa & AIA  |  baa & AIA  ;
 CAA <=  BAA & AKA  |  baa & aka  |  baa & AKA  |  BAA & aka  ;
 ccb <=  BAA & AKA  |  baa & aka  |  baa & AKA  |  baa & AKA  ;
 EAB <=  BAB & bcb  |  bab & BCB  ; 
 EBB <=  BAB & bcb  |  bab & BCB  ; 
 CAB <=  BAB & bcb & AKB  |  bab & BCB & AKB  |  bab & bcb & akb  |  BAB & BCB & akb  ;
 ccc <=  BAB & bcb & AKB  |  bab & BCB & AKB  |  bab & bcb & akb  |  bab & bcb & AKB  ;
 EAC <=  BAC & bcc  |  bac & BCC  ; 
 EBC <=  BAC & bcc  |  bac & BCC  ; 
 CEC <=  BAC & bcc & AIC  |  bac & BCC & AIC  |  bac & bcc & aic  |  BAC & BCC & aic  ;
 cgd <=  BAC & bcc & AIC  |  bac & BCC & AIC  |  bac & bcc & aic  |  bac & bcc & AIC  ;
 CAC <=  BAC & bcc & AKC  |  bac & BCC & AKC  |  bac & bcc & akc  |  BAC & BCC & akc  ;
 ccd <=  BAC & bcc & AKC  |  bac & BCC & AKC  |  bac & bcc & akc  |  bac & bcc & AKC  ;
 EAD <=  BAD & bcd  |  bad & BCD  ; 
 EBD <=  BAD & bcd  |  bad & BCD  ; 
 CED <=  BAD & bcd & AID  |  bad & BCD & AID  |  bad & bcd & aid  |  BAD & BCD & aid  ;
 cge <=  BAD & bcd & AID  |  bad & BCD & AID  |  bad & bcd & aid  |  bad & bcd & AID  ;
 CAD <=  BAD & bcd & AKD  |  bad & BCD & AKD  |  bad & bcd & akd  |  BAD & BCD & akd  ;
 cce <=  BAD & bcd & AKD  |  bad & BCD & AKD  |  bad & bcd & akd  |  bad & bcd & AKD  ;
 TNA <= qra & thd ; 
 TNB <= qra & thd ; 
 TNC <= qra & thd ; 
 TND <= qra & thd ; 
 tha <= tga ; 
 thb <= tga ; 
 thc <= tga ; 
 thd <= tga ; 
 FAA <=  IIA & tha  |  PJA & THA  ; 
 FAB <=  IIB & tha  |  PJB & THA  ; 
 FAC <=  IIC & tha  |  PJC & THA  ; 
 FAD <=  IID & tha  |  PJD & THA  ; 
 CEB <=  BAB & bcb & AIB  |  bab & BCB & AIB  |  bab & bcb & aib  |  BAB & BCB & aib  ;
 cgc <=  BAB & bcb & AIB  |  bab & BCB & AIB  |  bab & bcb & aib  |  bab & bcb & AIB  ;
 FAE <=  IIE & tha  |  PJE & THA  ; 
 FAF <=  IIF & tha  |  PJF & THA  ; 
 AAA <=  IAA & TAA  |  QAC & TAC  |  AAA & TAE  ; 
 AAB <=  IAB & TAA  |  BCB & TAC  |  AAB & TAE  ; 
 AGA <=  IAA & TDA  |  IEA & TDC  |  AGA & TDE  ; 
 AGB <=  IAB & TDA  |  IEB & TDC  |  AGB & TDE  ; 
 aia <=  iea & TEA  |  aia & tea  ; 
 aib <=  ieb & TEA  |  aib & tea  ; 
 ACA <=  IGA & TBA  |  BAA & TBC  |  ACA & TBE  ; 
 ACB <=  IGB & TBA  |  BAB & TBC  |  ACB & TBE  ; 
 AEA <=  ICA & TCA  |  AGA & TCC  |  AIA & TCE  ; 
 AEB <=  ICB & TCA  |  AGB & TCC  |  AIB & TCE  ; 
 aka <=  iea & TFA  |  aka & tfa  ; 
 akb <=  ieb & TFA  |  akb & tfa  ; 
 AAC <=  IAC & TAB  |  BCC & TAD  |  AAC & TAF  ; 
 AAD <=  IAD & TAB  |  BCD & TAD  |  AAD & TAF  ; 
 AGC <=  IAC & TDB  |  IEC & TDD  |  AGC & TDF  ; 
 AGD <=  IAD & TDB  |  IED & TDD  |  AGD & TDF  ; 
 aic <=  iec & TEB  |  aic & teb  ; 
 aid <=  ied & TEB  |  aid & teb  ; 
 ACC <=  IGC & TBB  |  BAC & TBD  |  ACC & TBF  ; 
 ACD <=  IGD & TBB  |  BAD & TBD  |  ACD & TBF  ; 
 AEC <=  ICC & TCB  |  AGC & TCD  |  AIC & TCF  ; 
 AED <=  ICD & TCB  |  AGD & TCD  |  AID & TCF  ; 
 akc <=  iec & TFB  |  akc & tfb  ; 
 akd <=  ied & TFB  |  akd & tfb  ; 
 TMA <= THA ; 
 TMB <= THA ; 
 TMC <= THA ; 
 TMD <= THA ; 
 QAC <= IKF ; 
 TGA <= IKB ; 
 TGB <= IKB ; 
 OHE <= QME ; 
 OAM <=  WAM & tid & tif  |  PCQ & TIC  |  JFA & TIA  ; 
 WAM <=  WAM & tid & tif  |  PCQ & TIC  |  JFA & TIA  ; 
 QMA <=  KBA  |  KBB  |  KBC  |  KBD  |  KAA  ; 
 QME <=  KBA  |  KBB  |  KBC  |  KBD  |  KAA  ; 
 OAA <=  WAA & tic & tie  |  PCA & TIC  |  FAA & TIA  ; 
 WAA <=  WAA & tic & tie  |  PCA & TIC  |  FAA & TIA  ; 
 OAB <=  WAB & tic & tie  |  PCB & TIC  |  FAB & TIA  ; 
 WAB <=  WAB & tic & tie  |  PCB & TIC  |  FAB & TIA  ; 
 QBA <=  QAA & eab & thc  |  PJM & THC  ; 
 QBE <=  QAA & eab & thc  |  PJM & THC  ; 
 OAC <=  WAC & tic & tie  |  PCC & TIC  |  FAC & TIA  ; 
 WAC <=  WAC & tic & tie  |  PCC & TIC  |  FAC & TIA  ; 
 OAD <=  WAD & tic & tie  |  PCD & TIC  |  FAD & TIA  ; 
 WAD <=  WAD & tic & tie  |  PCD & TIC  |  FAD & TIA  ; 
 QGA <= QFA ; 
 TIC <= QGA ; 
 TID <= QGA ; 
 qta <= ike ; 
 oha <=  kbd & kba & kbb & kbc  ; 
 OAE <=  WAE & tic & tie  |  PCE & TIC  |  FAE & TIA  ; 
 WAE <=  WAE & tic & tie  |  PCE & TIC  |  FAE & TIA  ; 
 OAF <=  WAF & tic & tie  |  PCF & TIC  |  FAF & TIA  ; 
 WAF <=  WAF & tic & tie  |  PCF & TIC  |  FAF & TIA  ; 
 pag <= fag ; 
 pbg <= pag ; 
 pcg <= pbg ; 
 pdg <= pcg ; 
 peg <= pdg ; 
 pfg <= peg ; 
 pgg <= pfg ; 
 phg <= pgg ; 
 pig <= phg ; 
 pih <= phh ; 
 pjg <= pig ; 
 pah <= fah ; 
 pbh <= pah ; 
 pch <= pbh ; 
 pdh <= pch ; 
 peh <= pdh ; 
 pfh <= peh ; 
 pgh <= pfh ; 
 phh <= pgh ; 
 dae <=  bae  |  bce  |  TGA  ; 
 daf <=  baf  |  bcf  |  TGA  ; 
 pai <= fai ; 
 pbi <= pai ; 
 pci <= pbi ; 
 pdi <= pci ; 
 pei <= pdi ; 
 pfi <= pei ; 
 pgi <= pfi ; 
 phi <= pgi ; 
 pii <= phi ; 
 pji <= pii ; 
 pjh <= pih ; 
 dag <=  bag  |  bcg  |  TGB  ; 
 dah <=  bah  |  bch  |  TGB  ; 
 paj <= faj ; 
 pbj <= paj ; 
 pcj <= pbj ; 
 pdj <= pcj ; 
 pej <= pdj ; 
 pfj <= pej ; 
 pgj <= pfj ; 
 phj <= pgj ; 
 pak <= fak ; 
 pbk <= pak ; 
 pck <= pbk ; 
 pdk <= pck ; 
 pek <= pdk ; 
 pfk <= pek ; 
 pgk <= pfk ; 
 phk <= pgk ; 
 pik <= phk ; 
 pjk <= pik ; 
 pij <= phj ; 
 pjj <= pij ; 
 FEM <=  JAG & EAG  |  DAG  ; 
 FEN <=  JAG & EAG  |  DAG  ; 
 paq <= jfa ; 
 pbq <= paq ; 
 pcq <= pbq ; 
 pdq <= pcq ; 
 peq <= pdq ; 
 pfq <= peq ; 
 pgq <= pfq ; 
 phq <= pgq ; 
 QNB <= QMA ; 
 QNC <= QNB ; 
 QND <= QNC ; 
 QNE <= QND ; 
 QNF <= QNE ; 
 QNG <= QNF ; 
 QNH <= QNG ; 
 QNI <= QNH ; 
 pao <= qbc ; 
 pbo <= pao ; 
 pco <= pbo ; 
 pdo <= pco ; 
 peo <= pdo ; 
 pfo <= peo ; 
 pgo <= pfo ; 
 pho <= pgo ; 
 pjo <= pio ; 
 pio <= pho ; 
 MBA <=  LCA & LDB & LDC & LDD  |  LCB & LDC & LDD  |  LCC & LDD  |  LCD  ; 
 pap <= qbd ; 
 pbp <= pap ; 
 pcp <= pbp ; 
 pdp <= pcp ; 
 pep <= pdp ; 
 pfp <= pep ; 
 pgp <= pfp ; 
 php <= pgp ; 
 pip <= php ; 
 pjp <= pip ; 
 QNJ <=  qnf  |  qng  |  qnh  |  qni  ; 
 EAE <=  BAE & bee  |  bae & BEE  ; 
 EBE <=  BAE & bee  |  bae & BEE  ; 
 CEE <=  BAE & bce & AIE  |  bae & BCE & AIE  |  bae & bce & aie  |  BAE & BCE & aie  ;
 cgf <=  BAE & bce & AIE  |  bae & BCE & AIE  |  bae & bce & aie  |  bae & bce & AIE  ;
 CAE <=  BAE & bce & AKE  |  bae & BCE & AKE  |  bae & bce & ake  |  BAE & BCE & ake  ;
 ccf <=  BAE & bce & AKE  |  bae & BCE & AKE  |  bae & bce & ake  |  bae & bce & AKE  ;
 EAF <=  BAF & bcf  |  baf & BCF  ; 
 EBF <=  BAF & bcf  |  baf & BCF  ; 
 CEF <=  BAF & bcf & AIF  |  baf & BCF & AIF  |  baf & bcf & aif  |  BAF & BCF & aif  ;
 cgg <=  BAF & bcf & AIF  |  baf & BCF & AIF  |  baf & bcf & aif  |  baf & bcf & AIF  ;
 CAF <=  BAF & bcf & AKF  |  baf & BCF & AKF  |  baf & bcf & akf  |  BAF & BCF & akf  ;
 ccg <=  BAF & bcf & AKF  |  baf & BCF & AKF  |  baf & bcf & akf  |  baf & bcf & AKF  ;
 EAG <=  BAG & bcg  |  bag & BCG  ; 
 EBG <=  BAG & bcg  |  bag & BCG  ; 
 CEG <=  BAG & bcg & AIG  |  bag & BCG & AIG  |  bag & bcg & aig  |  BAG & BCG & aig  ;
 cgh <=  BAG & bcg & AIG  |  bag & BCG & AIG  |  bag & bcg & aig  |  bag & bcg & AIG  ;
 CAG <=  BAG & bcg & AKG  |  bag & BCG & AKG  |  bag & bcg & akg  |  BAG & BCG & akg  ;
 cch <=  BAG & bcg & AKG  |  bag & BCG & AKG  |  bag & bcg & akg  |  bag & bcg & AKG  ;
 EAH <=  BAH & bch  |  bah & BCH  ; 
 EBH <=  BAH & bch  |  bah & BCH  ; 
 CEH <=  BAH & bch & AIH  |  bah & BCH & AIH  |  bah & bch & aih  |  BAH & BCH & aih  ;
 cgi <=  BAH & bch & AIH  |  bah & BCH & AIH  |  bah & bch & aih  |  bah & bch & AIH  ;
 CAH <=  BAH & bch & AKH  |  bah & BCH & AKH  |  bah & bch & akh  |  BAH & BCH & akh  ;
 cci <=  BAH & bch & AKH  |  bah & BCH & AKH  |  bah & bch & akh  |  bah & bch & AKH  ;
 FAG <=  EBC & jac & thb  |  PJG & THB  |  ebc & JAC  ; 
 FAH <=  EBD & jad & thb  |  PJH & THB  |  ebd & JAD  ; 
 QNA <=  qma  |  qnb  |  qnc  |  qnd  |  qne  ; 
 FAI <=  EBE & jae & thb  |  PJI & THB  |  ebe & JAE  ; 
 FAJ <=  EBF & jaf & thb  |  PJJ & THB  |  ebf & JAF  ; 
 FEA <=  JAG & EAG  |  DAG  ; 
 FEI <=  JAG & EAG  |  DAG  ; 
 FAK <=  EBG & jag & thb  |  PJK & THB  |  ebg & JAG  ; 
 FAL <=  EBG & jag & thb  |  PJK & THB  |  ebg & JAG  ; 
 AAE <=  IAE & TAA  |  BCE & TAC  |  AAE & TAE  ; 
 AAF <=  IAF & TAA  |  BCF & TAC  |  AAF & TAE  ; 
 AGE <=  IAE & TDA  |  IEE & TDC  |  AGE & TDE  ; 
 AGF <=  IAF & TDA  |  IEF & TDC  |  AGF & TDE  ; 
 aie <=  iee & TEA  |  aie & tea  ; 
 aif <=  ief & TEA  |  aif & tea  ; 
 ACE <=  IGE & TBA  |  BAE & TBC  |  ACE & TBE  ; 
 ACF <=  IGF & TBA  |  BAF & TBC  |  ACF & TBE  ; 
 AEE <=  ICE & TCA  |  AGE & TCC  |  AIE & TCE  ; 
 AEF <=  ICF & TCA  |  AGF & TCC  |  AIF & TCE  ; 
 ake <=  iee & TFA  |  ake & tfa  ; 
 akf <=  ief & TFA  |  akf & tfa  ; 
 AAG <=  IAG & TAB  |  BCG & TAD  |  AAG & TAF  ; 
 AAH <=  IAH & TAB  |  BCH & TAD  |  AAH & TAF  ; 
 AGG <=  IAG & TDB  |  IEG & TDD  |  AGG & TDF  ; 
 AGH <=  IAH & TDB  |  IEH & TDD  |  AGH & TDF  ; 
 aig <=  ieg & TEB  |  aig & teb  ; 
 aih <=  ieh & TEB  |  aih & teb  ; 
 ACG <=  IGG & TBB  |  BAG & TBD  |  ACG & TBF  ; 
 ACH <=  IGH & TBB  |  BAH & TBD  |  ACH & TBF  ; 
 AEG <=  ICG & TCB  |  AGG & TCD  |  AIG & TCF  ; 
 AEH <=  ICH & TCB  |  AGH & TCD  |  AIH & TCF  ; 
 akg <=  ieg & TFB  |  akg & tfb  ; 
 akh <=  ieh & TFB  |  akh & tfb  ; 
 TAC <=  IKH  ; 
 TAD <=  IKH  ; 
 TAG <=  IKH  ; 
 TAA <= IKG ; 
 TAB <= IKG ; 
 OIA <= QDE ; 
 TAE <= IKI ; 
 TAF <= IKI ; 
 OAN <=  WAN & tid & tif  |  PCR & TID  |  JFB & TIB  ; 
 WAN <=  WAN & tid & tif  |  PCR & TID  |  JFB & TIB  ; 
 OIE <=  QCA & ija & ijb  |  QDA  |  KBE  ; 
 OLA <=  QCA & ija & ijb  |  QDA  |  KBE  ; 
 QCA <=  QCA & ija & ijb  |  QDA  |  KBE  ; 
 OAG <=  WAG & tid & tif  |  PCG & TID  |  FAG & TIB  ; 
 WAG <=  WAG & tid & tif  |  PCG & TID  |  FAG & TIB  ; 
 OAH <=  WAH & tid & tif  |  PCH & TID  |  FAH & TIB  ; 
 WAH <=  WAH & tid & tif  |  PCH & TID  |  FAH & TIB  ; 
 qda <=  qda & kbe  |  qda & qca  |  IJA  |  IJB  ; 
 qde <=  qda & kbe  |  qda & qca  |  IJA  |  IJB  ; 
 OAI <=  WAI & tid & tif  |  PCI & TID  |  FAI & TIB  ; 
 WAI <=  WAI & tid & tif  |  PCI & TID  |  FAI & TIB  ; 
 OAJ <=  WAJ & tid & tif  |  PCJ & TID  |  FAJ & TIB  ; 
 WAJ <=  WAJ & tid & tif  |  PCJ & TID  |  FAJ & TIB  ; 
 QEB <= IKD ; 
 ofa <= kbe ; 
 QFA <=  KCA & WAK  |  KCA & WAL  ; 
 OAK <=  WAK & tid & tif  |  pck & TID  |  fal & TIB  ; 
 WAK <=  WAK & tid & tif  |  pck & TID  |  fal & TIB  ; 
 OAL <=  WAL & tid & tif  |  PCK & TID  |  FAL & TIB  ; 
 WAL <=  WAL & tid & tif  |  PCK & TID  |  FAL & TIB  ; 
 dai <=  bai  |  bci  |  TGA  ; 
 daj <=  baj  |  bcj  |  TGA  ; 
 dak <=  bak  |  bck  |  TGB  ; 
 dal <=  bal  |  bcl  |  TGB  ; 
 piq <= phq ; 
 pjq <= piq ; 
 saa <= haa ; 
 sba <= saa ; 
 sca <= sba ; 
 sda <= sca ; 
 sea <= sda ; 
 sfa <= sea ; 
 sga <= sfa ; 
 sha <= sga ; 
 sia <= sha ; 
 sja <= sia ; 
 FCA <=  EAH  ; 
 FDA <=  eah  ; 
 sab <= hab ; 
 sbb <= sab ; 
 scb <= sbb ; 
 sdb <= scb ; 
 seb <= sdb ; 
 sfb <= seb ; 
 sgb <= sfb ; 
 shb <= sgb ; 
 sib <= shb ; 
 sjb <= sib ; 
 FCB <=  JDB & eai  |  jdb & EAI  ; 
 FDB <=  JEB & eai  |  jeb & EAI  ; 
 sac <= hac ; 
 sbc <= sac ; 
 scc <= sbc ; 
 sdc <= scc ; 
 sec <= sdc ; 
 sfc <= sec ; 
 sgc <= sfc ; 
 shc <= sgc ; 
 FCC <=  JDC & eaj  |  jdc & EAJ  ; 
 FDC <=  JEC & eaj  |  jec & EAJ  ; 
 sad <= had ; 
 sbd <= sad ; 
 scd <= sbd ; 
 sdd <= scd ; 
 sed <= sdd ; 
 sfd <= sed ; 
 sgd <= sfd ; 
 shd <= sgd ; 
 sid <= shd ; 
 sjd <= sid ; 
 sic <= shc ; 
 sjc <= sic ; 
 FCD <=  JDD & eak  |  jdd & EAK  ; 
 FDD <=  JED & eak  |  jed & EAK  ; 
 EAI <=  BAI & bei  |  bai & BEI  ; 
 CEI <=  BAI & bci & AII  |  bai & BCI & AII  |  bai & bci & aii  |  BAI & BCI & aii  ;
 cgj <=  BAI & bci & AII  |  bai & BCI & AII  |  bai & bci & aii  |  bai & bci & AII  ;
 CAI <=  BAI & bci & AKI  |  bai & BCI & AKI  |  bai & bci & aki  |  BAI & BCI & aki  ;
 ccj <=  BAI & bci & AKI  |  bai & BCI & AKI  |  bai & bci & aki  |  bai & bci & AKI  ;
 EAJ <=  BAJ & bcj  |  baj & BCJ  ; 
 CEJ <=  BAJ & bcj & AIJ  |  baj & BCJ & AIJ  |  baj & bcj & aij  |  BAJ & BCJ & aij  ;
 cgk <=  BAJ & bcj & AIJ  |  baj & BCJ & AIJ  |  baj & bcj & aij  |  baj & bcj & AIJ  ;
 CAJ <=  BAJ & bcj & AKJ  |  baj & BCJ & AKJ  |  baj & bcj & akj  |  BAJ & BCJ & akj  ;
 cck <=  BAJ & bcj & AKJ  |  baj & BCJ & AKJ  |  baj & bcj & akj  |  baj & bcj & AKJ  ;
 EAK <=  BAK & bck  |  bak & BCK  ; 
 CEK <=  BAK & bck & AIK  |  bak & BCK & AIK  |  bak & bck & aik  |  BAK & BCK & aik  ;
 cgl <=  BAK & bck & AIK  |  bak & BCK & AIK  |  bak & bck & aik  |  bak & bck & AIK  ;
 CAK <=  BAK & bck & AKK  |  bak & BCK & AKK  |  bak & bck & akk  |  BAK & BCK & akk  ;
 ccl <=  BAK & bck & AKK  |  bak & BCK & AKK  |  bak & bck & akk  |  bak & bck & AKK  ;
 EAL <=  BAL & bcl  |  bal & BCL  ; 
 CEL <=  BAL & bcl & AIL  |  bal & BCL & AIL  |  bal & bcl & ail  |  BAL & BCL & ail  ;
 cgm <=  BAL & bcl & AIL  |  bal & BCL & AIL  |  bal & bcl & ail  |  bal & bcl & AIL  ;
 CAL <=  BAL & bcl & AKL  |  bal & BCL & AKL  |  bal & bcl & akl  |  BAL & BCL & akl  ;
 ccm <=  BAL & bcl & AKL  |  bal & BCL & AKL  |  bal & bcl & akl  |  bal & bcl & AKL  ;
 HAA <=  FCA & gaa & tma  |  SJA & TMA  |  FDA & GAA  ; 
 OEA <=  FCA & gaa & tma  |  SJA & TMA  |  FDA & GAA  ; 
 FAM <= THD & PJQ ; 
 FAN <= THD & PJR ; 
 HAC <=  FCC & gaa & tmc  |  SJC & TMC  |  FDC & GAA  ; 
 OEC <=  FCC & gaa & tmc  |  SJC & TMC  |  FDC & GAA  ; 
 HAB <=  FCB & gaa & tmb  |  SJB & TMB  |  FDB & GAA  ; 
 OEB <=  FCB & gaa & tmb  |  SJB & TMB  |  FDB & GAA  ; 
 ffb <=  eah  |  eai  |  eaj  |  eak  ; 
 ffj <=  eah  |  eai  |  eaj  |  eak  ; 
 MAA <=  LAA & LBB & LBC & LBD  |  LAB & LBC & LBD  |  LAC & LBD  |  LAD  ; 
 FEB <=  JDD & EAK  |  DAK  ; 
 FEJ <=  JDD & EAK  |  DAK  ; 
 HAD <=  FCD & gaa & tmd  |  SJD & TMD  |  FDD & GAA  ; 
 OED <=  FCD & gaa & tmd  |  SJD & TMD  |  FDD & GAA  ; 
 AAI <=  IAI & TAA  |  BCI & TAC  |  AAI & TAE  ; 
 AAJ <=  IAJ & TAA  |  BCJ & TAC  |  AAJ & TAE  ; 
 AGI <=  IAI & TDA  |  IEI & TDC  |  AGI & TDE  ; 
 AGJ <=  IAJ & TDA  |  IEJ & TDC  |  AGJ & TDE  ; 
 aii <=  iei & TEA  |  aii & tea  ; 
 aij <=  iej & TEA  |  aij & tea  ; 
 ACI <=  IGI & TBA  |  BAI & TBC  |  ACI & TBE  ; 
 ACJ <=  IGJ & TBA  |  BAJ & TBC  |  ACJ & TBE  ; 
 AEI <=  ICI & TCA  |  AGI & TCC  |  AII & TCE  ; 
 AEJ <=  ICJ & TCA  |  AGJ & TCC  |  AIJ & TCE  ; 
 aki <=  iei & TFA  |  aki & tfa  ; 
 akj <=  iej & TFA  |  akj & tfa  ; 
 AAK <=  IAK & TAB  |  BCK & TAD  |  AAK & TAF  ; 
 AAL <=  IAL & TAB  |  BCL & TAD  |  AAL & TAF  ; 
 AGK <=  IAK & TDB  |  IEK & TDD  |  AGK & TDF  ; 
 AGL <=  IAL & TDB  |  IEL & TDD  |  AGL & TDF  ; 
 aik <=  iek & TEB  |  aik & teb  ; 
 ail <=  iel & TEB  |  ail & teb  ; 
 ACK <=  IGK & TBB  |  BAK & TBD  |  ACK & TBF  ; 
 ACL <=  IGL & TBB  |  BAL & TBD  |  ACL & TBF  ; 
 AEK <=  ICK & TCB  |  AGK & TCD  |  AIK & TCF  ; 
 AEL <=  ICL & TCB  |  AGL & TCD  |  AIL & TCF  ; 
 akk <=  iek & TFB  |  akk & tfb  ; 
 akl <=  iel & TFB  |  akl & tfb  ; 
 TBA <= IKJ ; 
 TBB <= IKJ ; 
 TBC <= IKK ; 
 TBD <= IKK ; 
 TBE <= IKM ; 
 TBF <= IKM ; 
 OBM <=  WBM & tjc & tje  |  PCQ & TJC  |  JFA & TJA  ; 
 WBM <=  WBM & tjc & tje  |  PCQ & TJC  |  JFA & TJA  ; 
 QMB <=  KBA  |  KBB  |  KBC  |  KBD  |  KAA  ; 
 QMF <=  KBA  |  KBB  |  KBC  |  KBD  |  KAA  ; 
 OBA <=  WBA & tjc & tje  |  PCA & TJC  |  FAA & TJA  ; 
 WBA <=  WBA & tjc & tje  |  PCA & TJC  |  FAA & TJA  ; 
 OBB <=  WBB & tjc & tje  |  PCB & TJC  |  FAB & TJA  ; 
 WBB <=  WBB & tjc & tje  |  PCB & TJC  |  FAB & TJA  ; 
 QBB <=  QAB & eab & thc  |  PJN & THC  ; 
 QBF <=  QAB & eab & thc  |  PJN & THC  ; 
 OBC <=  WBC & tjc & tje  |  PCC & TJC  |  FAC & TJA  ; 
 WBC <=  WBC & tjc & tje  |  PCC & TJC  |  FAC & TJA  ; 
 OBD <=  WBD & tjc & tje  |  PCD & TJC  |  FAD & TJA  ; 
 WBD <=  WBD & tjc & tje  |  PCD & TJC  |  FAD & TJA  ; 
 QGB <= QFB ; 
 TJC <= QGB ; 
 TJD <= QGB ; 
 qtb <= qta ; 
 ohb <=  kbd & kba & kbb & kbc  ; 
 OBE <=  WBE & tjc & tje  |  PCE & TJC  |  FAE & TJA  ; 
 WBE <=  WBE & tjc & tje  |  PCE & TJC  |  FAE & TJA  ; 
 OBF <=  WBF & tjc & tje  |  PCF & TJC  |  FAF & TJA  ; 
 WBF <=  WBF & tjc & tje  |  PCF & TJC  |  FAF & TJA  ; 
 dam <=  bam  |  bcm  |  TGA  ; 
 dan <=  ban  |  bcn  |  TGA  ; 
 dao <=  bao  |  bco  |  TGB  ; 
 dap <=  bap  |  bcp  |  TGB  ; 
 sae <= hae ; 
 sbe <= sae ; 
 sce <= sbe ; 
 sde <= sce ; 
 see <= sde ; 
 sfe <= see ; 
 sge <= sfe ; 
 she <= sge ; 
 sie <= she ; 
 sje <= sie ; 
 FCE <=  EAL  ; 
 FDE <=  eal  ; 
 saf <= haf ; 
 sbf <= saf ; 
 scf <= sbf ; 
 sdf <= scf ; 
 sef <= sdf ; 
 sff <= sef ; 
 sgf <= sff ; 
 shf <= sgf ; 
 sif <= shf ; 
 sig <= shg ; 
 FCF <=  JDF & eam  |  jdf & EAM  ; 
 FDF <=  JEF & eam  |  jef & EAM  ; 
 sag <= hag ; 
 sbg <= sag ; 
 scg <= sbg ; 
 sdg <= scg ; 
 seg <= sdg ; 
 sfg <= seg ; 
 sgg <= sfg ; 
 shg <= sgg ; 
 sjg <= sig ; 
 FCG <=  JDG & ean  |  jdg & EAN  ; 
 FDG <=  JEG & ean  |  jeg & EAN  ; 
 sah <= hah ; 
 sbh <= sah ; 
 sch <= sbh ; 
 sdh <= sch ; 
 seh <= sdh ; 
 sfh <= seh ; 
 sgh <= sfh ; 
 shh <= sgh ; 
 sih <= shh ; 
 sjh <= sih ; 
 sjf <= sif ; 
 FCH <=  JDH & eao  |  jdh & EAO  ; 
 FDH <=  JEH & eao  |  jeh & EAO  ; 
 EAM <=  BAM & bem  |  bam & BEM  ; 
 CEM <=  BAM & bcm & AIM  |  bam & BCM & AIM  |  bam & bcm & aim  |  BAM & BCM & aim  ;
 cgn <=  BAM & bcm & AIM  |  bam & BCM & AIM  |  bam & bcm & aim  |  bam & bcm & AIM  ;
 CAM <=  BAM & bcm & AKM  |  bam & BCM & AKM  |  bam & bcm & akm  |  BAM & BCM & akm  ;
 ccn <=  BAM & bcm & AKM  |  bam & BCM & AKM  |  bam & bcm & akm  |  bam & bcm & AKM  ;
 EAN <=  BAM & bcn  |  ban & BCN  ; 
 CEN <=  BAN & bcn & AIN  |  ban & BCN & AIN  |  ban & bcn & ain  |  BAN & BCN & ain  ;
 cgo <=  BAN & bcn & AIN  |  ban & BCN & AIN  |  ban & bcn & ain  |  ban & bcn & AIN  ;
 CAN <=  BAN & bcn & AKN  |  ban & BCN & AKN  |  ban & bcn & akn  |  BAN & BCN & akn  ;
 cco <=  BAN & bcn & AKN  |  ban & BCN & AKN  |  ban & bcn & akn  |  ban & bcn & AKN  ;
 EAO <=  BAO & bco  |  bao & BCO  ; 
 CEO <=  BAO & bco & AIO  |  bao & BCO & AIO  |  bao & bco & aio  |  BAO & BCO & aio  ;
 cgp <=  BAO & bco & AIO  |  bao & BCO & AIO  |  bao & bco & aio  |  bao & bco & AIO  ;
 EAP <=  BAP & bcp  |  bap & BCP  ; 
 CEP <=  BAP & bcp & AIP  |  bap & BCP & AIP  |  bap & bcp & aip  |  BAP & BCP & aip  ;
 cha <=  BAP & bcp & AIP  |  bap & BCP & AIP  |  bap & bcp & aip  |  bap & bcp & AIP  ;
 CAP <=  BAP & bcp & AKP  |  bap & BCP & AKP  |  bap & bcp & akp  |  BAP & BCP & akp  ;
 cda <=  BAP & bcp & AKP  |  bap & BCP & AKP  |  bap & bcp & akp  |  bap & bcp & AKP  ;
 HAE <=  FCE & gab & tma  |  SJE & TMA  |  FDE & GAB  ; 
 OEE <=  FCE & gab & tma  |  SJE & TMA  |  FDE & GAB  ; 
 MBB <=  LCE & LDF & LDG & LDH  |  LCF & LDG & LDH  |  LCG & LDH  |  LCH  ; 
 MAB <=  LAE & LBF & LBG & LBH  |  LAF & LBG & LBH  |  LAG & LBH  |  LAH  ; 
 HAF <=  FCF & gab & tmb  |  SJF & TMB  |  FDF & GAB  ; 
 OEF <=  FCF & gab & tmb  |  SJF & TMB  |  FDF & GAB  ; 
 ffc <=  eal  |  eam  |  ean  |  eao  ; 
 ffk <=  eal  |  eam  |  ean  |  eao  ; 
 nab <=  lbe  |  lbf  |  lbg  |  lbh  ; 
 HAG <=  FCG & gab & tmc  |  SJG & TMC  |  FDG & GAB  ; 
 OEG <=  FCG & gab & tmc  |  SJG & TMC  |  FDG & GAB  ; 
 FEC <=  JDH & EAO  |  DAO  ; 
 FEK <=  JDH & EAO  |  DAO  ; 
 HAH <=  FCH & gab & tmd  |  SJH & TMD  |  FDH & GAB  ; 
 OEH <=  FCH & gab & tmd  |  SJH & TMD  |  FDH & GAB  ; 
 AAM <=  IAM & TAA  |  BCM & TAC  |  AAM & TAE  ; 
 AAN <=  IAN & TAA  |  BCN & TAC  |  AAN & TAE  ; 
 AGM <=  IAM & TDA  |  IEM & TDC  |  AGM & TDE  ; 
 AGN <=  IAN & TDA  |  IEN & TDC  |  AGN & TDE  ; 
 aim <=  iem & TEA  |  aim & tea  ; 
 ain <=  ien & TEA  |  ain & tea  ; 
 ACM <=  IGM & TBA  |  BAM & TBC  |  ACM & TBE  ; 
 ACN <=  IGN & TBA  |  BAN & TBC  |  ACN & TBE  ; 
 AEM <=  ICM & TCA  |  AGM & TCC  |  AIM & TCE  ; 
 AEN <=  ICN & TCA  |  AGN & TCC  |  AIN & TCE  ; 
 akm <=  iem & TFA  |  akm & tfa  ; 
 akn <=  ien & TFA  |  akn & tfa  ; 
 AAO <=  IAO & TAB  |  BCO & TAD  |  AAO & TAF  ; 
 AAP <=  IAP & TAB  |  BCP & TAD  |  AAP & TAF  ; 
 AGO <=  IAO & TDB  |  IEO & TDD  |  AGO & TDF  ; 
 AGP <=  IAP & TDB  |  IEP & TDD  |  AGP & TDF  ; 
 aio <=  ieo & TEB  |  aio & teb  ; 
 aip <=  iep & TEB  |  aip & teb  ; 
 ACO <=  IGO & TBB  |  BAO & TBD  |  ACO & TBF  ; 
 ACP <=  IGP & TBB  |  BAP & TBD  |  ACP & TBF  ; 
 AEO <=  ICO & TCB  |  AGO & TCD  |  AIO & TCF  ; 
 AEP <=  ICP & TCB  |  AGP & TCD  |  AIP & TCF  ; 
 ako <=  ieo & TFB  |  ako & tfb  ; 
 akp <=  iep & TFB  |  akp & tfb  ; 
 QRB <= QRA ; 
 OIB <= QDF ; 
 QRA <=  ILA & TCG  |  QRA & TAG  ; 
 OBN <=  WBN & tjd & tjf  |  PCR & TJD  |  JFB & TJB  ; 
 WBN <=  WBN & tjd & tjf  |  PCR & TJD  |  JFB & TJB  ; 
 OIF <=  QCB & ijc & ijd  |  QDB  |  KBF  ; 
 OLB <=  QCB & ijc & ijd  |  QDB  |  KBF  ; 
 QCB <=  QCB & ijc & ijd  |  QDB  |  KBF  ; 
 OBG <=  WBG & tjd & tjf  |  PCG & TJD  |  FAG & TJB  ; 
 WBG <=  WBG & tjd & tjf  |  PCG & TJD  |  FAG & TJB  ; 
 OBH <=  WBH & tjd & tjf  |  PCH & TJD  |  FAH & TJB  ; 
 WBH <=  WBH & tjd & tjf  |  PCH & TJD  |  FAH & TJB  ; 
 qdb <=  qdb & kbf  |  qdb & qcb  |  IJC  |  IJD  ; 
 qdf <=  qdb & kbf  |  qdb & qcb  |  IJC  |  IJD  ; 
 OBI <=  WBI & tjd & tjf  |  PCI & TJD  |  FAI & TJB  ; 
 WBI <=  WBI & tjd & tjf  |  PCI & TJD  |  FAI & TJB  ; 
 OBJ <=  WBJ & tjd & tjf  |  PCJ & TJD  |  FAJ & TJB  ; 
 WBJ <=  WBJ & tjd & tjf  |  PCJ & TJD  |  FAJ & TJB  ; 
 ofb <= kbf ; 
 QFB <=  KCB & WBK  |  KCB & WBL  ; 
 OBK <=  WBK & tjd & tjf  |  pck & TJD  |  fal & TJB  ; 
 WBK <=  WBK & tjd & tjf  |  pck & TJD  |  fal & TJB  ; 
 OBL <=  WBL & tjd & tjf  |  PCK & TJD  |  FAL & TJB  ; 
 WBL <=  WBL & tjd & tjf  |  PCK & TJD  |  FAL & TJB  ; 
 sak <= hak ; 
 sbk <= sak ; 
 sck <= sbk ; 
 sdk <= sck ; 
 FCL <=  JDL & edc  |  jdl & EDC  ; 
 FDL <=  JEL & edc  |  jel & EDC  ; 
 dba <=  bba  |  bda  |  TGA  ; 
 dbb <=  bbb  |  bdb  |  TGA  ; 
 sik <= shk ; 
 sil <= shl ; 
 sjl <= sil ; 
 dbc <=  bbc  |  bdc  |  TGB  ; 
 dbd <=  bbd  |  bdd  |  TGB  ; 
 sai <= hai ; 
 sbi <= sai ; 
 sci <= sbi ; 
 sdi <= sci ; 
 sei <= sdi ; 
 sfi <= sei ; 
 sgi <= sfi ; 
 shi <= sgi ; 
 sii <= shi ; 
 sji <= sii ; 
 FCI <=  EAP  ; 
 FDI <=  eae  ; 
 saj <= haj ; 
 sbj <= saj ; 
 scj <= sbj ; 
 sdj <= scj ; 
 sej <= sdj ; 
 sfj <= sej ; 
 sgj <= sfj ; 
 shj <= sgj ; 
 sij <= shj ; 
 sjj <= sij ; 
 FCJ <=  JDJ & eda  |  jdj & EDA  ; 
 FDJ <=  JEJ & eda  |  jej & EDA  ; 
 ffd <=  eap  |  eda  |  edb  |  edc  ; 
 ffl <=  eap  |  eda  |  edb  |  edc  ; 
 sek <= sdk ; 
 sfk <= sek ; 
 sgk <= sfk ; 
 shk <= sgk ; 
 sjk <= sik ; 
 FCK <=  JDK & edb  |  jdk & EDB  ; 
 FDK <=  JEK & edb  |  jek & EDB  ; 
 sal <= hal ; 
 sbl <= sal ; 
 scl <= sbl ; 
 sdl <= scl ; 
 sel <= sdl ; 
 sfl <= sel ; 
 sgl <= sfl ; 
 shl <= sgl ; 
 OEL <=  FCL & gac & tmd  |  SJL & TMD  |  FDL & GAC  ; 
 EDA <=  BBA & bfa  |  bba & BFA  ; 
 CFA <=  BBA & bda & AJA  |  bba & BDA & AJA  |  bba & bda & aja  |  BBA & BDA & aja  ;
 chb <=  BBA & bda & AJA  |  bba & BDA & AJA  |  bba & bda & aja  |  bba & bda & AJA  ;
 CBA <=  BBA & bda & ALA  |  bba & BDA & ALA  |  bba & bda & ala  |  BBA & BDA & ala  ;
 cdb <=  BBA & bda & ALA  |  bba & BDA & ALA  |  bba & bda & ala  |  bba & bda & ALA  ;
 EDB <=  BBB & bdb & BDB  |  bbb & BDB  ; 
 CFB <=  BBB & bdb & AJB  |  bbb & BDB & AJB  |  bbb & bdb & ajb  |  BBB & BDB & ajb  ;
 chc <=  BBB & bdb & AJB  |  bbb & BDB & AJB  |  bbb & bdb & ajb  |  bbb & bdb & AJB  ;
 CBB <=  BBB & bdb & ALB  |  bbb & BDB & ALB  |  bbb & bdb & alb  |  BBB & BDB & alb  ;
 cdc <=  BBB & bdb & ALB  |  bbb & BDB & ALB  |  bbb & bdb & alb  |  bbb & bdb & ALB  ;
 EDC <=  BBC & bdc  |  bbc & BDC  ; 
 CFC <=  BBC & bdc & AJC  |  bbc & BDC & AJC  |  bbc & bdc & ajc  |  BBC & BDC & ajc  ;
 chd <=  BBC & bdc & AJC  |  bbc & BDC & AJC  |  bbc & bdc & ajc  |  bbc & bdc & AJC  ;
 CBC <=  BBC & bdc & ALC  |  bbc & BDC & ALC  |  bbc & bdc & alc  |  BBC & BDC & alc  ;
 cdd <=  BBC & bdc & ALC  |  bbc & BDC & ALC  |  bbc & bdc & alc  |  bbc & bdc & ALC  ;
 EDD <=  BBD & bdd  |  bbd & BDD  ; 
 CFD <=  BBD & bdd & AJD  |  bbd & BDD & AJD  |  bbd & bdd & ajd  |  BBD & BDD & ajd  ;
 che <=  BBD & bdd & AJD  |  bbd & BDD & AJD  |  bbd & bdd & ajd  |  bbd & bdd & AJD  ;
 CBD <=  BBD & bdd & ALD  |  bbd & BDD & ALD  |  bbd & bdd & ald  |  BBD & BDD & ald  ;
 cde <=  BBD & bdd & ALD  |  bbd & BDD & ALD  |  bbd & bdd & ald  |  bbd & bdd & ALD  ;
 HAI <=  FCI & gac & tma  |  SJI & TMA  |  FDI & GAC  ; 
 OEI <=  FCI & gac & tma  |  SJI & TMA  |  FDI & GAC  ; 
 MBC <=  LCI & LDJ & LDK & LDL  |  LCJ & LDK & LDL  |  LCK & LDL  |  LCL  ; 
 MAC <=  LAI & LBJ & LBK & LBL  |  LAJ & LBK & LBL  |  LAK & LBL  |  LAL  ; 
 HAJ <=  FCJ & gac & tmb  |  SJJ & TMB  |  FDJ & GAC  ; 
 OEJ <=  FCJ & gac & tmb  |  SJJ & TMB  |  FDJ & GAC  ; 
 HAK <=  FCK & gac & tmc  |  SJK & TMC  |  FDK & GAC  ; 
 OEK <=  FCK & gac & tmc  |  SJK & TMC  |  FDK & GAC  ; 
 FED <=  JDL & EDC  |  DBC  ; 
 FEL <=  JDL & EDC  |  DBC  ; 
 HAL <=  FCL & gac & tmd  |  SJL & TMD  |  FDL & GAC  ; 
 ABA <=  IBA & TAA  |  BDA & TAC  |  ABA & TAE  ; 
 ABB <=  IBB & TAA  |  BDB & TAC  |  ABB & TAE  ; 
 AHA <=  IBA & TDA  |  IFA & TDC  |  AHA & TDE  ; 
 AHB <=  IBB & TDA  |  IFB & TDC  |  AHB & TDE  ; 
 aja <=  ifa & TEA  |  aja & tea  ; 
 ajb <=  ifb & TEA  |  ajb & tea  ; 
 ADA <=  IHA & TBA  |  BBA & TBC  |  ADA & TBE  ; 
 ADB <=  IHB & TBA  |  BBB & TBC  |  ADB & TBE  ; 
 AFA <=  IDA & TCA  |  AHA & TCC  |  AJA & TCE  ; 
 AFB <=  IDB & TCA  |  AHB & TCC  |  AJB & TCE  ; 
 ala <=  ifa & TFA  |  ala & tfa  ; 
 alb <=  ifb & TFA  |  alb & tfa  ; 
 ABC <=  IBC & TAB  |  BDC & TAD  |  ABC & TAF  ; 
 ABD <=  IBD & TAB  |  BDD & TAD  |  ABD & TAF  ; 
 AHC <=  IBC & TDB  |  IFC & TDD  |  AHC & TDF  ; 
 AHD <=  IBD & TDB  |  IFD & TDD  |  AHD & TDF  ; 
 ajc <=  ifc & TEB  |  ajc & teb  ; 
 ajd <=  ifd & TEB  |  ajd & teb  ; 
 ADC <=  IHC & TBB  |  BBC & TBD  |  ADC & TBF  ; 
 ADD <=  IHD & TBB  |  BBD & TBD  |  ADD & TBF  ; 
 AFC <=  IDC & TCB  |  AHC & TCD  |  AJC & TCF  ; 
 AFD <=  IDD & TCB  |  AHD & TCD  |  AJD & TCF  ; 
 alc <=  ifc & TFB  |  alc & tfb  ; 
 ald <=  ifd & TFB  |  ald & tfb  ; 
 TDA <= IKQ ; 
 TDB <= IKQ ; 
 TDC <= IKR ; 
 TDD <= IKR ; 
 TDE <= IKS ; 
 TDF <= IKS ; 
 OCM <=  WCM & tkc & tke  |  PCQ & TKC  |  JFA & TKA  ; 
 WCM <=  WCM & tkc & tke  |  PCQ & TKC  |  JFA & TKA  ; 
 QMC <=  KBA  |  KBB  |  KBC  |  KBD  |  KAA  ; 
 QMG <=  KBA  |  KBB  |  KBC  |  KBD  |  KAA  ; 
 OCA <=  WCA & tkc & tke  |  PCA & TKC  |  FAA & TKA  ; 
 WCA <=  WCA & tkc & tke  |  PCA & TKC  |  FAA & TKA  ; 
 OCB <=  WCB & tkc & tke  |  PCB & TKC  |  FAB & TKA  ; 
 WCB <=  WCB & tkc & tke  |  PCB & TKC  |  FAB & TKA  ; 
 QBC <=  QAA & EAB & thc  |  PJO & THC  ; 
 QBG <=  QAA & EAB & thc  |  PJO & THC  ; 
 OCC <=  WCC & tkc & tke  |  PCC & TKC  |  FAC & TKA  ; 
 WCC <=  WCC & tkc & tke  |  PCC & TKC  |  FAC & TKA  ; 
 OCD <=  WCD & tkc & tke  |  PCD & TKC  |  FAD & TKA  ; 
 WCD <=  WCD & tkc & tke  |  PCD & TKC  |  FAD & TKA  ; 
 QGC <= QFC ; 
 TKC <= QGC ; 
 TKD <= QGC ; 
 qtc <= qtb ; 
 ohc <=  kbd & kba & kbb & kbc  ; 
 OCE <=  WCE & tkc & tke  |  PCE & TKC  |  FAE & TKA  ; 
 WCE <=  WCE & tkc & tke  |  PCE & TKC  |  FAE & TKA  ; 
 OCF <=  WCF & tkc & tke  |  PCF & TKC  |  FAF & TKA  ; 
 WCF <=  WCF & tkc & tke  |  PCF & TKC  |  FAF & TKA  ; 
 dbe <=  bbe  |  bde  |  TGA  ; 
 dbf <=  bbf  |  bdf  |  TGA  ; 
 dbg <=  bbg  |  bdg  |  TGB  ; 
 dbh <=  bbh  |  bdh  |  TGB  ; 
 sam <= ham ; 
 sbm <= sam ; 
 scm <= sbm ; 
 sdm <= scm ; 
 sem <= sdm ; 
 sfm <= sem ; 
 sgm <= sfm ; 
 shm <= sgm ; 
 sim <= shm ; 
 sjm <= sim ; 
 FCM <=  EDD  ; 
 FDM <=  edd  ; 
 san <= han ; 
 sbn <= san ; 
 scn <= sbn ; 
 sdn <= scn ; 
 sen <= sdn ; 
 sfn <= sen ; 
 sgn <= sfn ; 
 shn <= sgn ; 
 sin <= shn ; 
 sjn <= sin ; 
 FCN <=  JDN & ede  |  jdn & EDE  ; 
 FDN <=  JEN & ede  |  jen & EDE  ; 
 sao <= hao ; 
 sbo <= sao ; 
 sco <= sbo ; 
 sdo <= sco ; 
 seo <= sdo ; 
 sfo <= seo ; 
 sgo <= sfo ; 
 sho <= sgo ; 
 sjo <= sio ; 
 sio <= sho ; 
 FCO <=  JDO & edf  |  jdo & EDF  ; 
 FDO <=  JEO & edf  |  jeo & EDF  ; 
 sap <= hap ; 
 sbp <= sap ; 
 scp <= sbp ; 
 sdp <= scp ; 
 sep <= sdp ; 
 sfp <= sep ; 
 sgp <= sfp ; 
 shp <= sgp ; 
 sip <= shp ; 
 sjp <= sip ; 
 FCP <=  JDP & edg  |  jdp & EDG  ; 
 FDP <=  JEP & edg  |  jep & EDG  ; 
 EDE <=  BBE & bfe  |  bbe & BFE  ; 
 CFE <=  BBE & bde & AJE  |  bbe & BDE & AJE  |  bbe & bde & aje  |  BBE & BDE & aje  ;
 chf <=  BBE & bde & AJE  |  bbe & BDE & AJE  |  bbe & bde & aje  |  bbe & bde & AJE  ;
 CBE <=  BBE & bde & ALE  |  bbe & BDE & ALE  |  bbe & bde & ale  |  BBE & BDE & ale  ;
 cdf <=  BBE & bde & ALE  |  bbe & BDE & ALE  |  bbe & bde & ale  |  bbe & bde & ALE  ;
 EDF <=  BBF & bdf  |  bbf & BDF  ; 
 CFF <=  BBF & bdf & AJF  |  bbf & BDF & AJF  |  bbf & bdf & ajf  |  BBF & BDF & ajf  ;
 chg <=  BBF & bdf & AJF  |  bbf & BDF & AJF  |  bbf & bdf & ajf  |  bbf & bdf & AJF  ;
 CBF <=  BBF & bdf & ALF  |  bbf & BDF & ALF  |  bbf & bdf & alf  |  BBF & BDF & alf  ;
 cdg <=  BBF & bdf & ALF  |  bbf & BDF & ALF  |  bbf & bdf & alf  |  bbf & bdf & ALF  ;
 EDG <=  BBG & bdg  |  bbg & BDG  ; 
 CFG <=  BBG & bdg & AJG  |  bbg & BDG & AJG  |  bbg & bdg & ajg  |  BBG & BDG & ajg  ;
 chh <=  BBG & bdg & AJG  |  bbg & BDG & AJG  |  bbg & bdg & ajg  |  bbg & bdg & AJG  ;
 CBG <=  BBG & bdg & ALG  |  bbg & BDG & ALG  |  bbg & bdg & alg  |  BBG & BDG & alg  ;
 cdh <=  BBG & bdg & ALG  |  bbg & BDG & ALG  |  bbg & bdg & alg  |  bbg & bdg & ALG  ;
 EDH <=  BBH & bdh  |  bbh & BDH  ; 
 CFH <=  BBH & bdh & AJH  |  bbh & BDH & AJH  |  bbh & bdh & ajh  |  BBH & BDH & ajh  ;
 chi <=  BBH & bdh & AJH  |  bbh & BDH & AJH  |  bbh & bdh & ajh  |  bbh & bdh & AJH  ;
 CBH <=  BBH & bdh & ALH  |  bbh & BDH & ALH  |  bbh & bdh & alh  |  BBH & BDH & alh  ;
 cdi <=  BBH & bdh & ALH  |  bbh & BDH & ALH  |  bbh & bdh & alh  |  bbh & bdh & ALH  ;
 HAM <=  FCM & gad & tma  |  SJM & TMA  |  FDM & GAD  ; 
 OEM <=  FCM & gad & tma  |  SJM & TMA  |  FDM & GAD  ; 
 nbb <=  lde  |  ldf  |  ldg  |  ldh  ; 
 nac <=  lbi  |  lbj  |  lbk  |  lbl  ; 
 HAN <=  FCN & gad & tmb  |  SJN & TMB  |  FDN & GAD  ; 
 OEN <=  FCN & gad & tmb  |  SJN & TMB  |  FDN & GAD  ; 
 ffe <=  edd  |  ede  |  edf  |  edg  ; 
 ffm <=  edd  |  ede  |  edf  |  edg  ; 
 HAO <=  FCO & gad & tmc  |  SJO & TMC  |  FDO & GAD  ; 
 OEO <=  FCO & gad & tmc  |  SJO & TMC  |  FDO & GAD  ; 
 FEE <=  JDP & EDG  |  DBG  ; 
 HAP <=  FCP & gad & tmd  |  SJP & TMD  |  FDP & GAD  ; 
 OEP <=  FCP & gad & tmd  |  SJP & TMD  |  FDP & GAD  ; 
 ABE <=  IBE & TAA  |  BDE & TAC  |  ABE & TAE  ; 
 ABF <=  IBF & TAA  |  BDF & TAC  |  ABF & TAE  ; 
 AHE <=  IBE & TDA  |  IFE & TDC  |  AHE & TDE  ; 
 AHF <=  IBF & TDA  |  IFFF  & TDC  |  AHF & TDE  ; 
 aje <=  ife & TEA  |  aje & tea  ; 
 ajf <=  ifff  & TEA  |  ajf & tea  ; 
 ADE <=  IHE & TBA  |  BBE & TBC  |  ADE & TBE  ; 
 ADF <=  IHF & TBA  |  BBF & TBC  |  ADF & TBE  ; 
 AFE <=  IDE & TCA  |  AHE & TCC  |  AJE & TCE  ; 
 AFF <=  IDF & TCA  |  AHF & TCC  |  AJF & TCE  ; 
 ale <=  ife & TFA  |  ale & tfa  ; 
 alf <=  ifff  & TFA  |  alf & tfa  ; 
 ABG <=  IBG & TAB  |  BDG & TAD  |  ABG & TAF  ; 
 ABH <=  IBH & TAB  |  BDH & TAD  |  ABH & TAF  ; 
 AHG <=  IBG & TDB  |  IFG & TDD  |  AHG & TDF  ; 
 AHH <=  IBH & TDB  |  IFH & TDD  |  AHH & TDF  ; 
 ajg <=  ifg & TEB  |  ajg & teb  ; 
 ajh <=  ifh & TEB  |  ajh & teb  ; 
 ADG <=  IHG & TBB  |  BBG & TBD  |  ADG & TBF  ; 
 ADH <=  IHH & TBB  |  BBH & TBD  |  ADH & TBF  ; 
 AFG <=  IDG & TCB  |  AHG & TCD  |  AJG & TCF  ; 
 AFH <=  IDH & TCB  |  AHH & TCD  |  AJH & TCF  ; 
 alg <=  ifg & TFB  |  alg & tfb  ; 
 alh <=  ifh & TFB  |  alh & tfb  ; 
 TCA <=  IKN  ; 
 TCB <=  IKN  ; 
 TCG <=  IKN  ; 
 TCC <= IKO ; 
 TCD <= IKO ; 
 OIC <= QDG ; 
 TCE <= IKP ; 
 TCF <= IKP ; 
 OCN <=  WCN & tkd & tkf  |  PCR & TKD  |  JFB & TKB  ; 
 WCN <=  WCN & tkd & tkf  |  PCR & TKD  |  JFB & TKB  ; 
 OIG <=  QCC & ije & ijf  |  QDC  |  KBG  ; 
 OLC <=  QCC & ije & ijf  |  QDC  |  KBG  ; 
 QCC <=  QCC & ije & ijf  |  QDC  |  KBG  ; 
 OCG <=  WCG & tkd & tkf  |  PCG & TKD  |  FAG & TKB  ; 
 WCG <=  WCG & tkd & tkf  |  PCG & TKD  |  FAG & TKB  ; 
 OCH <=  WCH & tkd & tkf  |  PCH & TKD  |  FAH & TKB  ; 
 WCH <=  WCH & tkd & tkf  |  PCH & TKD  |  FAH & TKB  ; 
 qdc <=  qdc & kbg  |  qdc & qcc  |  IJE  |  IJF  ; 
 qdg <=  qdc & kbg  |  qdc & qcc  |  IJE  |  IJF  ; 
 OCI <=  WCI & tkd & tkf  |  PCI & TKD  |  FAI & TKB  ; 
 WCI <=  WCI & tkd & tkf  |  PCI & TKD  |  FAI & TKB  ; 
 OCJ <=  WCJ & tkd & tkf  |  PCJ & TKD  |  FAJ & TKB  ; 
 WCJ <=  WCJ & tkd & tkf  |  PCJ & TKD  |  FAJ & TKB  ; 
 ofc <= kbg ; 
 QFC <=  KCC & WCK  |  KCC & WCL  ; 
 OCK <=  WCK & tkd & tkf  |  pck & TKD  |  fal & TKB  ; 
 WCK <=  WCK & tkd & tkf  |  pck & TKD  |  fal & TKB  ; 
 OCL <=  WCL & tkd & tkf  |  PCK & TKD  |  FAL & TKB  ; 
 WCL <=  WCL & tkd & tkf  |  PCK & TKD  |  FAL & TKB  ; 
 dbi <=  bbi  |  bdi  |  TGA  ; 
 dbj <=  bbj  |  bdj  |  TGA  ; 
 dbk <=  bbk  |  bdk  |  TGB  ; 
 dbl <=  bbl  |  bdl  |  TGB  ; 
 saq <= haq ; 
 sbq <= saq ; 
 scq <= sbq ; 
 sdq <= scq ; 
 seq <= sdq ; 
 sfq <= seq ; 
 sgq <= sfq ; 
 shq <= sgq ; 
 siq <= shq ; 
 sjq <= siq ; 
 FCQ <=  EDH  ; 
 FDQ <=  edh  ; 
 sar <= har ; 
 sbr <= sar ; 
 scr <= sbr ; 
 sdr <= scr ; 
 ser <= sdr ; 
 sfr <= ser ; 
 sgr <= sfr ; 
 shr <= sgr ; 
 sir <= shr ; 
 sjr <= sir ; 
 FCR <=  JDR & edi  |  jdr & EDI  ; 
 FDR <=  JER & edi  |  jer & EDI  ; 
 sas <= has ; 
 sbs <= sas ; 
 scs <= sbs ; 
 sds <= scs ; 
 ses <= sds ; 
 sfs <= ses ; 
 sgs <= sfs ; 
 shs <= sgs ; 
 sis <= shs ; 
 sjs <= sis ; 
 FCS <=  JDS & edj  |  jds & EDJ  ; 
 FDS <=  JES & edj  |  jes & EDJ  ; 
 sat <= hat ; 
 sbt <= sat ; 
 sct <= sbt ; 
 sdt <= sct ; 
 set <= sdt ; 
 sft <= set ; 
 sgt <= sft ; 
 sht <= sgt ; 
 sit <= sht ; 
 sjt <= sit ; 
 FCT <=  JDT & edk  |  jdt & EDK  ; 
 FDT <=  JET & edk  |  jet & EDK  ; 
 EDI <=  BBI & bfi  |  bbi & BFI  ; 
 CFI <=  BBI & bdi & AJI  |  bbi & BDI & AJI  |  bbi & bdi & aji  |  BBI & BDI & aji  ;
 chj <=  BBI & bdi & AJI  |  bbi & BDI & AJI  |  bbi & bdi & aji  |  bbi & bdi & AJI  ;
 CBI <=  BBI & bdi & ALI  |  bbi & BDI & ALI  |  bbi & bdi & ali  |  BBI & BDI & ali  ;
 cdj <=  BBI & bdi & ALI  |  bbi & BDI & ALI  |  bbi & bdi & ali  |  bbi & bdi & ALI  ;
 EDJ <=  BBJ & bdj  |  bbj & BDJ  ; 
 CFJ <=  BBJ & bdj & AJJ  |  bbj & BDJ & AJJ  |  bbj & bdj & ajj  |  BBJ & BDJ & ajj  ;
 chk <=  BBJ & bdj & AJJ  |  bbj & BDJ & AJJ  |  bbj & bdj & ajj  |  bbj & bdj & AJJ  ;
 CBJ <=  BBJ & bdj & ALJ  |  bbj & BDJ & ALJ  |  bbj & bdj & alj  |  BBJ & BDJ & alj  ;
 cdk <=  BBJ & bdj & ALJ  |  bbj & BDJ & ALJ  |  bbj & bdj & alj  |  bbj & bdj & ALJ  ;
 EDK <=  BBK & bdk  |  bbk & BDK  ; 
 CFK <=  BBK & bdk & AJK  |  bbk & BDK & AJK  |  bbk & bdk & ajk  |  BBK & BDK & ajk  ;
 chl <=  BBK & bdk & AJK  |  bbk & BDK & AJK  |  bbk & bdk & ajk  |  bbk & bdk & AJK  ;
 CBK <=  BBK & bdk & ALK  |  bbk & BDK & ALK  |  bbk & bdk & alk  |  BBK & BDK & alk  ;
 cdl <=  BBK & bdk & ALK  |  bbk & BDK & ALK  |  bbk & bdk & alk  |  bbk & bdk & ALK  ;
 EDL <=  BBL & bdl  |  bbl & BDL  ; 
 CFL <=  BBL & bdl & AJL  |  bbl & BDL & AJL  |  bbl & bdl & ajl  |  BBL & BDL & ajl  ;
 chm <=  BBL & bdl & AJL  |  bbl & BDL & AJL  |  bbl & bdl & ajl  |  bbl & bdl & AJL  ;
 CBL <=  BBL & bdl & ALL  |  bbl & BDL & ALL  |  bbl & bdl & all  |  BBL & BDL & all  ;
 cdm <=  BBL & bdl & ALL  |  bbl & BDL & ALL  |  bbl & bdl & all  |  bbl & bdl & ALL  ;
 HAQ <=  FCQ & gae & tma  |  SJQ & TMA  |  FDQ & GAE  ; 
 OEQ <=  FCQ & gae & tma  |  SJQ & TMA  |  FDQ & GAE  ; 
 nbc <=  ldi  |  ldj  |  ldk  |  ldl  ; 
 MAD <=  LAM & LBN & LBO & LBP  |  LAN & LBO & LBP  |  LAO & LBP  |  LAP  ; 
 HAR <=  FCR & gae & tmb  |  SJR & TMB  |  FDR & GAE  ; 
 OER <=  FCR & gae & tmb  |  SJR & TMB  |  FDR & GAE  ; 
 fff <=  edh  |  edi  |  edj  |  edk  ; 
 nad <=  lbm  |  lbn  |  lbo  |  lbp  ; 
 HAS <=  FCS & gae & tmc  |  SJS & TMC  |  FDS & GAE  ; 
 OES <=  FCS & gae & tmc  |  SJS & TMC  |  FDS & GAE  ; 
 FEF <=  JDT & EDK  |  DBK  ; 
 HAT <=  FCT & gae & tmd  |  SJT & TMD  |  FDT & GAE  ; 
 OET <=  FCT & gae & tmd  |  SJT & TMD  |  FDT & GAE  ; 
 ABI <=  IBI & TAA  |  BDI & TAC  |  ABI & TAE  ; 
 ABJ <=  IBJ & TAA  |  BDJ & TAC  |  ABJ & TAE  ; 
 AHI <=  IBI & TDA  |  IFI & TDC  |  AHI & TDE  ; 
 AHJ <=  IBJ & TDA  |  IFJ & TDC  |  AHJ & TDE  ; 
 aji <=  ifi & TEA  |  aji & tea  ; 
 ajj <=  ifj & TEA  |  ajj & tea  ; 
 ADI <=  IHI & TBA  |  BBI & TBC  |  ADI & TBE  ; 
 ADJ <=  IHJ & TBA  |  BBJ & TBC  |  ADJ & TBE  ; 
 AFI <=  IDI & TCA  |  AHI & TCC  |  AJI & TCE  ; 
 AFJ <=  IDJ & TCA  |  AHJ & TCC  |  AJJ & TCE  ; 
 ali <=  ifi & TFA  |  ali & tfa  ; 
 alj <=  ifj & TFA  |  alj & tfa  ; 
 ABK <=  IBK & TAB  |  BDK & TAD  |  ABK & TAF  ; 
 ABL <=  IBL & TAB  |  BDL & TAD  |  ABL & TAF  ; 
 AHK <=  IBK & TDB  |  IFK & TDD  |  AHK & TDF  ; 
 AHL <=  IBL & TDB  |  IFL & TDD  |  AHL & TDF  ; 
 ajk <=  ifk & TEB  |  ajk & teb  ; 
 ajl <=  ifl & TEB  |  ajl & teb  ; 
 ADK <=  IHK & TBB  |  BBK & TBD  |  ADK & TBF  ; 
 ADL <=  IHL & TBB  |  BBL & TBD  |  ADL & TBF  ; 
 AFK <=  IDK & TCB  |  AHK & TCD  |  AJK & TCF  ; 
 AFL <=  IDL & TCB  |  AHL & TCD  |  AJL & TCF  ; 
 alk <=  ifk & TFB  |  alk & tfb  ; 
 all <=  ifl & TFB  |  all & tfb  ; 
 TEA <= IKT ; 
 TEB <= IKT ; 
 TFA <= IKU ; 
 TFB <= IKU ; 
 ODM <=  WDM & tlc & tle  |  PCQ & TLC  |  JFA & TLA  ; 
 WDM <=  WDM & tlc & tle  |  PCQ & TLC  |  JFA & TLA  ; 
 QMD <=  KBA  |  KBB  |  KBC  |  KBD  |  KAA  ; 
 QMH <=  KBA  |  KBB  |  KBC  |  KBD  |  KAA  ; 
 ODA <=  WDA & tlc & tle  |  PCA & TLC  |  FAA & TLA  ; 
 WDA <=  WDA & tlc & tle  |  PCA & TLC  |  FAA & TLA  ; 
 ODB <=  WDB & tlc & tle  |  PCB & TLC  |  FAB & TLA  ; 
 WDB <=  WDB & tlc & tle  |  PCB & TLC  |  FAB & TLA  ; 
 QBD <=  QAB & EAB & thc  |  PJP & THC  ; 
 QBH <=  QAB & EAB & thc  |  PJP & THC  ; 
 ODC <=  WDC & tlc & tle  |  PCC & TLC  |  FAC & TLA  ; 
 WDC <=  WDC & tlc & tle  |  PCC & TLC  |  FAC & TLA  ; 
 ODD <=  WDD & tlc & tle  |  PCD & TLC  |  FAD & TLA  ; 
 WDD <=  WDD & tlc & tle  |  PCD & TLC  |  FAD & TLA  ; 
 QGD <= QFD ; 
 TLC <= QGD ; 
 TLD <= QGD ; 
 qtd <= qtc ; 
 ohd <=  kbd & kba & kbb & kbc  ; 
 ODE <=  WDE & tlc & tle  |  PCE & TLC  |  FAE & TLA  ; 
 WDE <=  WDE & tlc & tle  |  PCE & TLC  |  FAE & TLA  ; 
 ODF <=  WDF & tlc & tle  |  PCF & TLC  |  FAF & TLA  ; 
 WDF <=  WDF & tlc & tle  |  PCF & TLC  |  FAF & TLA  ; 
 dbm <=  bbm  |  bfm  |  TGA  ; 
 dbn <=  bbn  |  bdn  |  TGA  ; 
 siw <= shw ; 
 dbo <=  bbo  |  bdo  |  TGB  ; 
 dbp <=  bbp  |  bdp  |  TGB  ; 
 sau <= hau ; 
 sbu <= sau ; 
 scu <= sbu ; 
 sdu <= scu ; 
 seu <= sdu ; 
 sfu <= seu ; 
 sgu <= sfu ; 
 shu <= sgu ; 
 siu <= shu ; 
 sju <= siu ; 
 FCU <=  EDL  ; 
 FDU <=  edl  ; 
 sav <= hav ; 
 sbv <= sav ; 
 scv <= sbv ; 
 sdv <= scv ; 
 sev <= sdv ; 
 sfv <= sev ; 
 sgv <= sfv ; 
 shv <= sgv ; 
 siv <= shv ; 
 sjv <= siv ; 
 FCV <=  JDV & edm  |  jdv & EDM  ; 
 FDV <=  JEV & edm  |  jev & EDM  ; 
 sbw <= saw ; 
 scw <= sbw ; 
 sdw <= scw ; 
 saw <= haw ; 
 sew <= sdw ; 
 sfw <= sew ; 
 sgw <= sfw ; 
 shw <= sgw ; 
 sjw <= siw ; 
 sax <= hax ; 
 sbx <= sax ; 
 scx <= sbx ; 
 sdx <= scx ; 
 sex <= sdx ; 
 sfx <= sex ; 
 sgx <= sfx ; 
 shx <= sgx ; 
 six <= shx ; 
 sjx <= six ; 
 EDM <=  BBM & bfm  |  bbm & BFM  ; 
 CFM <=  BBM & bdm & AJM  |  bbm & BDM & AJM  |  bbm & bdm & ajm  |  BBM & BDM & ajm  ;
 chn <=  BBM & bdm & AJM  |  bbm & BDM & AJM  |  bbm & bdm & ajm  |  bbm & bdm & AJM  ;
 CBM <=  BBM & bdm & ALM  |  bbm & BDM & ALM  |  bbm & bdm & alm  |  BBM & BDM & alm  ;
 cdn <=  BBM & bdm & ALM  |  bbm & BDM & ALM  |  bbm & bdm & alm  |  bbm & bdm & ALM  ;
 EDN <=  BBN & bdn  |  bbn & BDN  ; 
 CFN <=  BBN & bdn & AJN  |  bbn & BDN & AJN  |  bbn & bdn & ajn  |  BBN & BDN & ajn  ;
 cho <=  BBN & bdn & AJN  |  bbn & BDN & AJN  |  bbn & bdn & ajn  |  bbn & bdn & AJN  ;
 CBN <=  BBN & bdn & ALN  |  bbn & BDN & ALN  |  bbn & bdn & aln  |  BBN & BDN & aln  ;
 cdo <=  BBN & bdn & ALN  |  bbn & BDN & ALN  |  bbn & bdn & aln  |  bbn & bdn & ALN  ;
 EDO <=  BBO & bdo  |  bbo & BDO  ; 
 CFO <=  BBO & bdo & AJO  |  bbo & BDO & AJO  |  bbo & bdo & ajo  |  BBO & BDO & ajo  ;
 chp <=  BBO & bdo & AJO  |  bbo & BDO & AJO  |  bbo & bdo & ajo  |  bbo & bdo & AJO  ;
 CBO <=  BBO & bdo & ALO  |  bbo & BDO & ALO  |  bbo & bdo & alo  |  BBO & BDO & alo  ;
 cdp <=  BBO & bdo & ALO  |  bbo & BDO & ALO  |  bbo & bdo & alo  |  bbo & bdo & ALO  ;
 EDP <=  BBP & bdp  |  bbp & BDP  ; 
 CFP <=  BBP & bdp & AJP  |  bbp & BDP & AJP  |  bbp & bdp & ajp  |  BBP & BDP & ajp  ;
 CBP <=  BBP & bdp & ALP  |  bbp & BDP & ALP  |  bbp & bdp & alp  |  BBP & BDP & alp  ;
 HAU <=  FCU & gaf & tma  |  SJU & TMA  |  FDU & GAF  ; 
 OEU <=  FCU & gaf & tma  |  SJU & TMA  |  FDU & GAF  ; 
 MBD <=  LCM & LDN & LDO & LDP  |  LCN & LDO & LDP  |  LCO & LDP  |  LCP  ; 
 HAV <=  QRB & tmb  |  SJV & TMB  ; 
 OEV <=  QRB & tmb  |  SJV & TMB  ; 
 nbd <=  ldm  |  ldn  |  ldo  |  ldp  ; 
 HAW <=  XAA & tmc  |  xab & tmc  |  KAB & tmc  ; 
 oex <=  XAA & tmc  |  xab & tmc  |  KAB & tmc  |  sjw & TMC  ; 
 HAX <=  KAB & xaa & tmd  |  SJX & TMD  ; 
 oew <=  XAA & tmd  |  xab & tmd  |  kab & tmd  |  sjx & TMD  ; 
 ABM <=  IBM & TAA  |  BDM & TAC  |  ABM & TAE  ; 
 ABN <=  IBN & TAA  |  BDN & TAC  |  ABN & TAE  ; 
 AHM <=  IBM & TDA  |  IFM & TDC  |  AHM & TDE  ; 
 AHN <=  IBN & TDA  |  IFN & TDC  |  AHN & TDE  ; 
 ajm <=  ifm & TEA  |  ajm & tea  ; 
 ajn <=  ifn & TEA  |  ajn & tea  ; 
 ADM <=  IHM & TBA  |  BBM & TBC  |  ADM & TBE  ; 
 ADN <=  IHN & TBA  |  BBN & TBC  |  ADN & TBE  ; 
 AFM <=  IDM & TCA  |  AHM & TCC  |  AJM & TCE  ; 
 AFN <=  IDN & TCA  |  AHN & TCC  |  AJN & TCE  ; 
 alm <=  ifm & TFA  |  alm & tfa  ; 
 aln <=  ifn & TFA  |  aln & tfa  ; 
 ABO <=  IBO & TAB  |  BDO & TAD  |  ABO & TAF  ; 
 ABP <=  IBP & TAB  |  BDP & TAD  |  ABP & TAF  ; 
 AHO <=  IBO & TDB  |  IFO & TDD  |  AHO & TDF  ; 
 AHP <=  IBP & TDB  |  IFP & TDD  |  AHP & TDF  ; 
 CAO <=  BAO & bco & AKO  |  bao & BCO & AKO  |  bao & bco & ako  |  BAO & BCO & ako  ;
 ccp <=  BAO & bco & AKO  |  bao & BCO & AKO  |  bao & bco & ako  |  bao & bco & AKO  ;
 ADO <=  IHO & TBB  |  BBO & TBD  |  ADO & TBF  ; 
 ADP <=  IHP & TBB  |  BBP & TBD  |  ADP & TBF  ; 
 AFO <=  IDO & TCB  |  AHO & TCD  |  AJO & TCF  ; 
 AFP <=  IDP & TCB  |  AHP & TCD  |  AJP & TCF  ; 
 alo <=  ifo & TFB  |  alo & tfb  ; 
 alp <=  ifp & TFB  |  alp & tfb  ; 
 OID <= QDH ; 
 QEA <= IKC ; 
 QEC <= IKC ; 
 ofd <= kbh ; 
 OKA <=  XAA  |  xab & QEC  ; 
 ODN <=  WDN & tld & tlf  |  PCR & TLD  |  JFB & TLB  ; 
 WDN <=  WDN & tld & tlf  |  PCR & TLD  |  JFB & TLB  ; 
 OIH <=  QCD & ijg & ijh  |  QDD  |  KBH  ; 
 OLD <=  QCD & ijg & ijh  |  QDD  |  KBH  ; 
 QCD <=  QCD & ijg & ijh  |  QDD  |  KBH  ; 
 ODG <=  WDG & tld & tlf  |  PCG & TLD  |  FAG & TLB  ; 
 WDG <=  WDG & tld & tlf  |  PCG & TLD  |  FAG & TLB  ; 
 ODH <=  WDH & tld & tlf  |  PCH & TLD  |  FAH & TLB  ; 
 WDH <=  WDH & tld & tlf  |  PCH & TLD  |  FAH & TLB  ; 
 qdd <=  qdd & kbh  |  qdd & qcd  |  IJG  |  IJH  ; 
 qdh <=  qdd & kbh  |  qdd & qcd  |  IJG  |  IJH  ; 
 ODI <=  WDI & tld & tlf  |  PCI & TLD  |  FAI & TLB  ; 
 WDI <=  WDI & tld & tlf  |  PCI & TLD  |  FAI & TLB  ; 
 ODJ <=  WDJ & tld & tlf  |  PCJ & TLD  |  FAJ & TLB  ; 
 WDJ <=  WDJ & tld & tlf  |  PCJ & TLD  |  FAJ & TLB  ; 
 ajo <=  ifo & TEB  |  ajo & teb  ; 
 ajp <=  ifp & TEB  |  ajp & teb  ; 
 QFD <=  KCD & WDK  |  KCD & WDL  ; 
 ODK <=  WDK & tld & tlf  |  pck & TLD  |  fal & TLB  ; 
 WDK <=  WDK & tld & tlf  |  pck & TLD  |  fal & TLB  ; 
 ODL <=  WDL & tld & tlf  |  PCK & TLD  |  FAL & TLB  ; 
 WDL <=  WDL & tld & tlf  |  PCK & TLD  |  FAL & TLB  ; 
end 
endmodule;
