module ka( IZZ,
 IAA, 
 IAB, 
 IAC, 
 IAD, 
 IAE, 
 IAF, 
 IAG, 
 IAH, 
 IAI, 
 IAJ, 
 IAK, 
 IAL, 
 IAM, 
 IAN, 
 IAO, 
 IAP, 
 IBA, 
 IBB, 
 IBC, 
 IBD, 
 IBE, 
 IBF, 
 IBG, 
 IBH, 
 IBI, 
 IBJ, 
 IBK, 
 IBL, 
 IBM, 
 IBN, 
 IBO, 
 IBP, 
 ICA, 
 ICB, 
 ICC, 
 ICD, 
 ICE, 
 IDA, 
 IDB, 
 IDC, 
 IFA, 
 IFB, 
 IFC, 
 IFD, 
 IFE, 
 IFFF , 
 IFG, 
 IFH, 
 IFI, 
 IFJ, 
 IFK, 
 IFL, 
 IGA, 
 IGB, 
 OAA, 
 OAB, 
 OAC, 
 OAD, 
 OAE, 
 OAF, 
 OAG, 
 OAH, 
 OAI, 
 OAJ, 
 OAK, 
 OAL, 
 OAM, 
 OAN, 
 OAO, 
 OAP, 
 OBA, 
 OBB, 
 OBC, 
 OBD, 
 OBE, 
 OBF, 
 OBG, 
 OBH, 
 OBI, 
 OBJ, 
 OBK, 
 OBL, 
 OBM, 
 OBN, 
 OBO, 
 OBP, 
 OCA, 
 OCB, 
 OCC, 
 OCD, 
 OCE, 
 OCF, 
 OCG, 
 OCH, 
 OCI, 
 OCJ, 
 OCK, 
 OCL, 
 ODA, 
 ODB, 
 ODC, 
 ODD, 
 ODE, 
 ODF, 
 ODG, 
 ODH, 
 ODI, 
 ODJ, 
 ODK, 
 ODL, 
 OEA, 
 OEB, 
 OEC, 
 OED, 
 OEE, 
 OEF, 
 OEG, 
 OEH, 
 OEI, 
 OEJ, 
 OEK, 
 OEL, 
 OEM, 
 OFA, 
 OFB, 
 OFC, 
 OFD, 
 OFE, 
 OFF, 
 OFG, 
 OFH, 
 OFI, 
 OFJ, 
 OFK, 
 OFL, 
 OGA, 
 OGB, 
 OGC, 
 OGD, 
 OGE, 
 OHA, 
 OHB, 
 OHC, 
 OHD, 
 OHE, 
 OHF, 
 OHG, 
 OHH, 
 OJA, 
 OJB, 
 OJC, 
 OJD, 
 OJE, 
 OJF, 
 OJG, 
 OJH, 
 OJI, 
 OJJ, 
 OJK, 
 OJL, 
 OJM, 
 OJN, 
OJO ); 
    
 input IZZ; 
 input IAA; 
 input IAB; 
 input IAC; 
 input IAD; 
 input IAE; 
 input IAF; 
 input IAG; 
 input IAH; 
 input IAI; 
 input IAJ; 
 input IAK; 
 input IAL; 
 input IAM; 
 input IAN; 
 input IAO; 
 input IAP; 
 input IBA; 
 input IBB; 
 input IBC; 
 input IBD; 
 input IBE; 
 input IBF; 
 input IBG; 
 input IBH; 
 input IBI; 
 input IBJ; 
 input IBK; 
 input IBL; 
 input IBM; 
 input IBN; 
 input IBO; 
 input IBP; 
 input ICA; 
 input ICB; 
 input ICC; 
 input ICD; 
 input ICE; 
 input IDA; 
 input IDB; 
 input IDC; 
 input IFA; 
 input IFB; 
 input IFC; 
 input IFD; 
 input IFE; 
 input IFFF ; 
 input IFG; 
 input IFH; 
 input IFI; 
 input IFJ; 
 input IFK; 
 input IFL; 
 input IGA; 
 input IGB; 
 output OAA; 
 output OAB; 
 output OAC; 
 output OAD; 
 output OAE; 
 output OAF; 
 output OAG; 
 output OAH; 
 output OAI; 
 output OAJ; 
 output OAK; 
 output OAL; 
 output OAM; 
 output OAN; 
 output OAO; 
 output OAP; 
 output OBA; 
 output OBB; 
 output OBC; 
 output OBD; 
 output OBE; 
 output OBF; 
 output OBG; 
 output OBH; 
 output OBI; 
 output OBJ; 
 output OBK; 
 output OBL; 
 output OBM; 
 output OBN; 
 output OBO; 
 output OBP; 
 output OCA; 
 output OCB; 
 output OCC; 
 output OCD; 
 output OCE; 
 output OCF; 
 output OCG; 
 output OCH; 
 output OCI; 
 output OCJ; 
 output OCK; 
 output OCL; 
 output ODA; 
 output ODB; 
 output ODC; 
 output ODD; 
 output ODE; 
 output ODF; 
 output ODG; 
 output ODH; 
 output ODI; 
 output ODJ; 
 output ODK; 
 output ODL; 
 output OEA; 
 output OEB; 
 output OEC; 
 output OED; 
 output OEE; 
 output OEF; 
 output OEG; 
 output OEH; 
 output OEI; 
 output OEJ; 
 output OEK; 
 output OEL; 
 output OEM; 
 output OFA; 
 output OFB; 
 output OFC; 
 output OFD; 
 output OFE; 
 output OFF; 
 output OFG; 
 output OFH; 
 output OFI; 
 output OFJ; 
 output OFK; 
 output OFL; 
 output OGA; 
 output OGB; 
 output OGC; 
 output OGD; 
 output OGE; 
 output OHA; 
 output OHB; 
 output OHC; 
 output OHD; 
 output OHE; 
 output OHF; 
 output OHG; 
 output OHH; 
 output OJA; 
 output OJB; 
 output OJC; 
 output OJD; 
 output OJE; 
 output OJF; 
 output OJG; 
 output OJH; 
 output OJI; 
 output OJJ; 
 output OJK; 
 output OJL; 
 output OJM; 
 output OJN; 
 output OJO; 
  
  
reg  AAA ;
reg  AAB ;
reg  AAC ;
reg  AAD ;
reg  AAE ;
reg  AAF ;
reg  AAG ;
reg  AAH ;
reg  AAI ;
reg  AAJ ;
reg  AAK ;
reg  AAL ;
reg  ABA ;
reg  ABB ;
reg  ABC ;
reg  ABD ;
reg  ABE ;
reg  ABF ;
reg  ABG ;
reg  ABH ;
reg  ABI ;
reg  ABJ ;
reg  ABK ;
reg  ABL ;
reg  ACA ;
reg  ACB ;
reg  ACC ;
reg  ACD ;
reg  ACE ;
reg  ACF ;
reg  ACG ;
reg  ACH ;
reg  ACI ;
reg  ACJ ;
reg  ACK ;
reg  ACL ;
reg  bab ;
reg  bac ;
reg  bad ;
reg  bae ;
reg  baf ;
reg  bag ;
reg  bah ;
reg  bai ;
reg  baj ;
reg  bak ;
reg  bal ;
reg  CAA ;
reg  CAB ;
reg  CAC ;
reg  CAD ;
reg  CAE ;
reg  CAF ;
reg  CAG ;
reg  CAH ;
reg  CBA ;
reg  CBB ;
reg  CBC ;
reg  CBD ;
reg  CBE ;
reg  CBF ;
reg  CBG ;
reg  CBH ;
reg  DBA ;
reg  DBB ;
reg  DBC ;
reg  DBD ;
reg  DBE ;
reg  DBF ;
reg  DBG ;
reg  DBH ;
reg  DCA ;
reg  DCB ;
reg  DCC ;
reg  DCD ;
reg  DCE ;
reg  DCF ;
reg  DCG ;
reg  DCH ;
reg  gaa ;
reg  gab ;
reg  gac ;
reg  gad ;
reg  gae ;
reg  gaf ;
reg  gag ;
reg  gah ;
reg  gai ;
reg  gba ;
reg  gbb ;
reg  gbc ;
reg  gbd ;
reg  gbe ;
reg  gbf ;
reg  gbg ;
reg  gbh ;
reg  gcf ;
reg  gcg ;
reg  gci ;
reg  gcj ;
reg  HAA ;
reg  HAB ;
reg  HAC ;
reg  HAD ;
reg  HAE ;
reg  HAF ;
reg  HAG ;
reg  HAH ;
reg  HAI ;
reg  HAJ ;
reg  HAK ;
reg  HAL ;
reg  HAM ;
reg  HAN ;
reg  HAO ;
reg  KAA ;
reg  KAB ;
reg  KAC ;
reg  KAD ;
reg  KAE ;
reg  KAF ;
reg  KAG ;
reg  KAH ;
reg  KAI ;
reg  KAJ ;
reg  KAK ;
reg  KAL ;
reg  KAM ;
reg  KAN ;
reg  KAO ;
reg  KAP ;
reg  KBA ;
reg  KBB ;
reg  KBC ;
reg  KBD ;
reg  KBE ;
reg  KBF ;
reg  KBG ;
reg  KBH ;
reg  KBI ;
reg  KBJ ;
reg  KBK ;
reg  KBL ;
reg  KBM ;
reg  KBN ;
reg  KBO ;
reg  KBP ;
reg  NAA ;
reg  NAB ;
reg  NAC ;
reg  NAD ;
reg  NAE ;
reg  NAF ;
reg  NAG ;
reg  NAH ;
reg  NAI ;
reg  NAJ ;
reg  NAK ;
reg  NAL ;
reg  NAM ;
reg  NAN ;
reg  NAO ;
reg  NAP ;
reg  NBA ;
reg  NBB ;
reg  NBC ;
reg  NBD ;
reg  NBE ;
reg  NBF ;
reg  NBG ;
reg  NBH ;
reg  NBI ;
reg  NBJ ;
reg  NBK ;
reg  NBL ;
reg  NBM ;
reg  NBN ;
reg  NBO ;
reg  NBP ;
reg  OAA ;
reg  OAB ;
reg  OAC ;
reg  OAD ;
reg  OAE ;
reg  OAF ;
reg  OAG ;
reg  OAH ;
reg  OAI ;
reg  OAJ ;
reg  OAK ;
reg  OAL ;
reg  OAM ;
reg  OAN ;
reg  OAO ;
reg  OAP ;
reg  OBA ;
reg  OBB ;
reg  OBC ;
reg  OBD ;
reg  OBE ;
reg  OBF ;
reg  OBG ;
reg  OBH ;
reg  OBI ;
reg  OBJ ;
reg  OBK ;
reg  OBL ;
reg  OBM ;
reg  OBN ;
reg  OBO ;
reg  OBP ;
reg  OCA ;
reg  OCB ;
reg  OCC ;
reg  OCD ;
reg  OCE ;
reg  OCF ;
reg  OCG ;
reg  OCH ;
reg  OCI ;
reg  OCJ ;
reg  OCK ;
reg  OCL ;
reg  ODA ;
reg  ODB ;
reg  ODC ;
reg  ODD ;
reg  ODE ;
reg  ODF ;
reg  ODG ;
reg  ODH ;
reg  ODI ;
reg  ODJ ;
reg  ODK ;
reg  ODL ;
reg  OEA ;
reg  OEB ;
reg  OEC ;
reg  OED ;
reg  OEE ;
reg  OEF ;
reg  OEG ;
reg  OEH ;
reg  OEI ;
reg  OEJ ;
reg  OEK ;
reg  OEL ;
reg  oem ;
reg  OFA ;
reg  OFB ;
reg  OFC ;
reg  OFD ;
reg  OFE ;
reg  OFF ;
reg  OFG ;
reg  OFH ;
reg  OFI ;
reg  OFJ ;
reg  OFK ;
reg  OFL ;
reg  OGA ;
reg  OGB ;
reg  OGC ;
reg  OGD ;
reg  OGE ;
reg  OHA ;
reg  OHB ;
reg  OHC ;
reg  OHD ;
reg  OHE ;
reg  OHF ;
reg  OHG ;
reg  OHH ;
reg  ohi ;
reg  OJA ;
reg  OJB ;
reg  OJC ;
reg  OJD ;
reg  OJE ;
reg  OJF ;
reg  OJG ;
reg  OJH ;
reg  OJI ;
reg  OJJ ;
reg  OJK ;
reg  OJL ;
reg  OJM ;
reg  OJN ;
reg  OJO ;
reg  PAA ;
reg  PAB ;
reg  PAC ;
reg  PAD ;
reg  PAE ;
reg  PAF ;
reg  PAG ;
reg  PAH ;
reg  PAJ ;
reg  PAK ;
reg  PAL ;
reg  PAM ;
reg  PAN ;
reg  PAO ;
reg  PAP ;
reg  PBA ;
reg  PBB ;
reg  PBC ;
reg  PBD ;
reg  PBE ;
reg  PBF ;
reg  PBG ;
reg  PBH ;
reg  PCA ;
reg  PCB ;
reg  PCC ;
reg  PCD ;
reg  PDA ;
reg  PDB ;
reg  PDC ;
reg  PDD ;
reg  PEA ;
reg  PEB ;
reg  PEC ;
reg  PED ;
reg  PFA ;
reg  PFB ;
reg  PFC ;
reg  PFD ;
reg  QAA ;
reg  QAB ;
reg  QAC ;
reg  QAD ;
reg  QAE ;
reg  QBA ;
reg  QBB ;
reg  QBC ;
reg  QBD ;
reg  QBE ;
reg  QBF ;
reg  QBG ;
reg  QBH ;
reg  qbi ;
reg  qbj ;
reg  qbk ;
reg  QBL ;
reg  qca ;
reg  QCB ;
reg  QCC ;
reg  qcd ;
reg  QCE ;
reg  QCF ;
reg  QCG ;
reg  QCI ;
reg  QCJ ;
reg  QDA ;
reg  QDB ;
reg  QDC ;
reg  QDE ;
reg  qdf ;
reg  qdg ;
reg  qdi ;
reg  qdj ;
reg  qdk ;
reg  qdl ;
reg  qea ;
reg  QEB ;
reg  QEI ;
reg  QEJ ;
reg  QEK ;
reg  QEL ;
reg  qfa ;
reg  QFB ;
reg  QFC ;
reg  qfd ;
reg  QFI ;
reg  qga ;
reg  QGB ;
reg  QGC ;
reg  qha ;
reg  QHB ;
reg  QHC ;
reg  QHD ;
reg  QHI ;
reg  qhj ;
reg  QHK ;
reg  qhl ;
reg  qia ;
reg  QIB ;
reg  QIC ;
reg  QID ;
reg  QIE ;
reg  QIF ;
reg  QIG ;
reg  qii ;
reg  qij ;
reg  qik ;
reg  qil ;
reg  qja ;
reg  QJB ;
reg  QJC ;
reg  QJD ;
reg  QJE ;
reg  QJF ;
reg  QJG ;
reg  QJH ;
reg  QJI ;
reg  qjj ;
reg  qjk ;
reg  qjl ;
reg  qka ;
reg  QKB ;
reg  QKC ;
reg  qkd ;
reg  qla ;
reg  QLB ;
reg  QLC ;
reg  qma ;
reg  QMB ;
reg  QMC ;
reg  QMD ;
reg  QME ;
reg  QMF ;
reg  QMI ;
reg  qmj ;
reg  qmk ;
reg  qna ;
reg  qnb ;
reg  qnc ;
reg  qnd ;
reg  qne ;
reg  QNF ;
reg  QNG ;
reg  qnh ;
reg  QNI ;
reg  QNJ ;
reg  QNK ;
reg  QNL ;
reg  QNM ;
reg  QNN ;
reg  QNO ;
reg  QNP ;
reg  qnq ;
reg  QNR ;
reg  qoa ;
reg  qob ;
reg  qoc ;
reg  qod ;
reg  QQA ;
reg  QQB ;
reg  QQC ;
reg  qqd ;
reg  qqe ;
reg  qqf ;
reg  QRA ;
reg  QRB ;
reg  QRC ;
reg  QRD ;
reg  QRE ;
reg  QRF ;
reg  QRG ;
reg  QRH ;
reg  QRI ;
reg  QRJ ;
reg  QRK ;
reg  QRL ;
reg  QRM ;
reg  QRN ;
reg  QRO ;
reg  QRP ;
reg  QRQ ;
reg  qrr ;
reg  QSA ;
reg  QSB ;
reg  QSC ;
reg  QSD ;
reg  QSI ;
reg  QSJ ;
reg  QSK ;
reg  QSL ;
reg  QSM ;
reg  QSN ;
reg  QSO ;
reg  QSP ;
reg  QSQ ;
reg  QTA ;
reg  QTB ;
reg  QTC ;
reg  QUA ;
reg  QUB ;
reg  QUC ;
reg  QVA ;
reg  QVB ;
reg  QVC ;
reg  RAA ;
reg  RAB ;
reg  RAC ;
reg  RAD ;
reg  RAE ;
reg  RAF ;
reg  RAG ;
reg  RAH ;
reg  RAI ;
reg  RAJ ;
reg  RAK ;
reg  RAL ;
reg  RAM ;
reg  RAN ;
reg  RAO ;
reg  RAP ;
reg  RBA ;
reg  RBB ;
reg  RBC ;
reg  RBD ;
reg  RBE ;
reg  RBF ;
reg  RBG ;
reg  RBH ;
reg  rbi ;
reg  rbj ;
reg  rbk ;
reg  rbl ;
reg  rbm ;
reg  RCA ;
reg  RCB ;
reg  RCC ;
reg  RCD ;
reg  RCE ;
reg  RCF ;
reg  RCG ;
reg  RCH ;
reg  RDA ;
reg  RDB ;
reg  RDC ;
reg  RDD ;
reg  RDE ;
reg  RDF ;
reg  RDG ;
reg  RDH ;
reg  REA ;
reg  RED ;
reg  REE ;
reg  REG ;
reg  RFA ;
reg  RFD ;
reg  RFE ;
reg  RFG ;
reg  RGA ;
reg  RGD ;
reg  RGE ;
reg  RGG ;
reg  RHA ;
reg  RHD ;
reg  RIA ;
reg  RID ;
reg  VAA ;
reg  VAB ;
reg  VAC ;
reg  VAD ;
reg  VAE ;
reg  VAF ;
reg  VAG ;
reg  VAH ;
reg  VBA ;
reg  VBB ;
reg  VBC ;
reg  VBD ;
reg  VBE ;
reg  VBF ;
reg  VBG ;
reg  VBH ;
wire  aaa ;
wire  aab ;
wire  aac ;
wire  aad ;
wire  aae ;
wire  aaf ;
wire  aag ;
wire  aah ;
wire  aai ;
wire  aaj ;
wire  aak ;
wire  aal ;
wire  aba ;
wire  abb ;
wire  abc ;
wire  abd ;
wire  abe ;
wire  abf ;
wire  abg ;
wire  abh ;
wire  abi ;
wire  abj ;
wire  abk ;
wire  abl ;
wire  aca ;
wire  acb ;
wire  acc ;
wire  acd ;
wire  ace ;
wire  acf ;
wire  acg ;
wire  ach ;
wire  aci ;
wire  acj ;
wire  ack ;
wire  acl ;
wire  BAB ;
wire  BAC ;
wire  BAD ;
wire  BAE ;
wire  BAF ;
wire  BAG ;
wire  BAH ;
wire  BAI ;
wire  BAJ ;
wire  BAK ;
wire  BAL ;
wire  caa ;
wire  cab ;
wire  cac ;
wire  cad ;
wire  cae ;
wire  caf ;
wire  cag ;
wire  cah ;
wire  cba ;
wire  cbb ;
wire  cbc ;
wire  cbd ;
wire  cbe ;
wire  cbf ;
wire  cbg ;
wire  cbh ;
wire  dba ;
wire  dbb ;
wire  dbc ;
wire  dbd ;
wire  dbe ;
wire  dbf ;
wire  dbg ;
wire  dbh ;
wire  dca ;
wire  dcb ;
wire  dcc ;
wire  dcd ;
wire  dce ;
wire  dcf ;
wire  dcg ;
wire  dch ;
wire  eaa ;
wire  EAA ;
wire  eab ;
wire  EAB ;
wire  eac ;
wire  EAC ;
wire  ead ;
wire  EAD ;
wire  eae ;
wire  EAE ;
wire  eaf ;
wire  EAF ;
wire  eag ;
wire  EAG ;
wire  eah ;
wire  EAH ;
wire  eai ;
wire  EAI ;
wire  eaj ;
wire  EAJ ;
wire  eak ;
wire  EAK ;
wire  eal ;
wire  EAL ;
wire  eba ;
wire  EBA ;
wire  ebb ;
wire  EBB ;
wire  ebc ;
wire  EBC ;
wire  ebd ;
wire  EBD ;
wire  ebe ;
wire  EBE ;
wire  ebf ;
wire  EBF ;
wire  ebg ;
wire  EBG ;
wire  ebh ;
wire  EBH ;
wire  faa ;
wire  FAA ;
wire  fab ;
wire  FAB ;
wire  fac ;
wire  FAC ;
wire  fad ;
wire  FAD ;
wire  fae ;
wire  FAE ;
wire  faf ;
wire  FAF ;
wire  fag ;
wire  FAG ;
wire  fah ;
wire  FAH ;
wire  fai ;
wire  FAI ;
wire  faj ;
wire  FAJ ;
wire  fak ;
wire  FAK ;
wire  fal ;
wire  FAL ;
wire  fba ;
wire  FBA ;
wire  fbb ;
wire  FBB ;
wire  fbc ;
wire  FBC ;
wire  fbd ;
wire  FBD ;
wire  fbe ;
wire  FBE ;
wire  fbf ;
wire  FBF ;
wire  fbg ;
wire  FBG ;
wire  fbh ;
wire  FBH ;
wire  fbi ;
wire  FBI ;
wire  fbj ;
wire  FBJ ;
wire  fbk ;
wire  FBK ;
wire  fbl ;
wire  FBL ;
wire  fca ;
wire  FCA ;
wire  fcb ;
wire  FCB ;
wire  fcc ;
wire  FCC ;
wire  fcd ;
wire  FCD ;
wire  fce ;
wire  FCE ;
wire  fcf ;
wire  FCF ;
wire  fcg ;
wire  FCG ;
wire  fch ;
wire  FCH ;
wire  fci ;
wire  FCI ;
wire  fcj ;
wire  FCJ ;
wire  fck ;
wire  FCK ;
wire  fcl ;
wire  FCL ;
wire  fda ;
wire  FDA ;
wire  fdb ;
wire  FDB ;
wire  fdc ;
wire  FDC ;
wire  fdd ;
wire  FDD ;
wire  fde ;
wire  FDE ;
wire  fdf ;
wire  FDF ;
wire  fdg ;
wire  FDG ;
wire  fdh ;
wire  FDH ;
wire  fdi ;
wire  FDI ;
wire  fdj ;
wire  FDJ ;
wire  fdk ;
wire  FDK ;
wire  fdl ;
wire  FDL ;
wire  fea ;
wire  FEA ;
wire  feb ;
wire  FEB ;
wire  fec ;
wire  FEC ;
wire  fed ;
wire  FED ;
wire  fee ;
wire  FEE ;
wire  fef ;
wire  FEF ;
wire  feg ;
wire  FEG ;
wire  feh ;
wire  FEH ;
wire  fei ;
wire  FEI ;
wire  fej ;
wire  FEJ ;
wire  fek ;
wire  FEK ;
wire  fel ;
wire  FEL ;
wire  ffa ;
wire  FFA ;
wire  ffb ;
wire  FFB ;
wire  ffc ;
wire  FFC ;
wire  ffd ;
wire  FFD ;
wire  ffe ;
wire  FFE ;
wire  fff ;
wire  FFF ;
wire  ffg ;
wire  FFG ;
wire  ffh ;
wire  FFH ;
wire  ffi ;
wire  FFI ;
wire  ffj ;
wire  FFJ ;
wire  ffk ;
wire  FFK ;
wire  ffl ;
wire  FFL ;
wire  fga ;
wire  FGA ;
wire  fgb ;
wire  FGB ;
wire  fgc ;
wire  FGC ;
wire  fgd ;
wire  FGD ;
wire  fge ;
wire  FGE ;
wire  fgf ;
wire  FGF ;
wire  fgg ;
wire  FGG ;
wire  fgh ;
wire  FGH ;
wire  fgi ;
wire  FGI ;
wire  fgj ;
wire  FGJ ;
wire  fgk ;
wire  FGK ;
wire  fgl ;
wire  FGL ;
wire  fha ;
wire  FHA ;
wire  fhb ;
wire  FHB ;
wire  fhc ;
wire  FHC ;
wire  fhd ;
wire  FHD ;
wire  fhe ;
wire  FHE ;
wire  fhf ;
wire  FHF ;
wire  fhg ;
wire  FHG ;
wire  fhh ;
wire  FHH ;
wire  fhi ;
wire  FHI ;
wire  fhj ;
wire  FHJ ;
wire  fhk ;
wire  FHK ;
wire  fhl ;
wire  FHL ;
wire  GAA ;
wire  GAB ;
wire  GAC ;
wire  GAD ;
wire  GAE ;
wire  GAF ;
wire  GAG ;
wire  GAH ;
wire  GAI ;
wire  GBA ;
wire  GBB ;
wire  GBC ;
wire  GBD ;
wire  GBE ;
wire  GBF ;
wire  GBG ;
wire  GBH ;
wire  GCF ;
wire  GCG ;
wire  GCI ;
wire  GCJ ;
wire  haa ;
wire  hab ;
wire  hac ;
wire  had ;
wire  hae ;
wire  haf ;
wire  hag ;
wire  hah ;
wire  hai ;
wire  haj ;
wire  hak ;
wire  hal ;
wire  ham ;
wire  han ;
wire  hao ;
wire  iaa ;
wire  iab ;
wire  iac ;
wire  iad ;
wire  iae ;
wire  iaf ;
wire  iag ;
wire  iah ;
wire  iai ;
wire  iaj ;
wire  iak ;
wire  ial ;
wire  iam ;
wire  ian ;
wire  iao ;
wire  iap ;
wire  iba ;
wire  ibb ;
wire  ibc ;
wire  ibd ;
wire  ibe ;
wire  ibf ;
wire  ibg ;
wire  ibh ;
wire  ibi ;
wire  ibj ;
wire  ibk ;
wire  ibl ;
wire  ibm ;
wire  ibn ;
wire  ibo ;
wire  ibp ;
wire  ica ;
wire  icb ;
wire  icc ;
wire  icd ;
wire  ice ;
wire  ida ;
wire  idb ;
wire  idc ;
wire  ifa ;
wire  ifb ;
wire  ifc ;
wire  ifd ;
wire  ife ;
wire  ifff  ;
wire  ifg ;
wire  ifh ;
wire  ifi ;
wire  ifj ;
wire  ifk ;
wire  ifl ;
wire  iga ;
wire  igb ;
wire  jaa ;
wire  JAA ;
wire  jab ;
wire  JAB ;
wire  jac ;
wire  JAC ;
wire  jak ;
wire  JAK ;
wire  jba ;
wire  JBA ;
wire  jbb ;
wire  JBB ;
wire  jbc ;
wire  JBC ;
wire  jbd ;
wire  JBD ;
wire  jbe ;
wire  JBE ;
wire  jbf ;
wire  JBF ;
wire  jbg ;
wire  JBG ;
wire  JCA ;
wire  JCB ;
wire  JCC ;
wire  JCD ;
wire  JCE ;
wire  JCF ;
wire  JCG ;
wire  JCH ;
wire  JCI ;
wire  jda ;
wire  JDA ;
wire  jea ;
wire  JEA ;
wire  jeb ;
wire  JEB ;
wire  jec ;
wire  JEC ;
wire  jed ;
wire  JED ;
wire  jfa ;
wire  JFA ;
wire  jfb ;
wire  JFB ;
wire  jfc ;
wire  JFC ;
wire  jfd ;
wire  JFD ;
wire  jfe ;
wire  JFE ;
wire  jff ;
wire  JFF ;
wire  jfg ;
wire  JFG ;
wire  jfh ;
wire  JFH ;
wire  jfi ;
wire  JFI ;
wire  jfj ;
wire  JFJ ;
wire  JGA ;
wire  JGB ;
wire  JGC ;
wire  JGD ;
wire  JGE ;
wire  JGF ;
wire  JGG ;
wire  JGH ;
wire  JGI ;
wire  jgj ;
wire  JGJ ;
wire  jgk ;
wire  JGK ;
wire  jha ;
wire  JHA ;
wire  jhb ;
wire  JHB ;
wire  jhc ;
wire  JHC ;
wire  jhd ;
wire  JHD ;
wire  jhe ;
wire  JHE ;
wire  jhf ;
wire  JHF ;
wire  jhg ;
wire  JHG ;
wire  jhh ;
wire  JHH ;
wire  jhi ;
wire  JHI ;
wire  jhj ;
wire  JHJ ;
wire  jhk ;
wire  JHK ;
wire  jia ;
wire  JIA ;
wire  jib ;
wire  JIB ;
wire  jma ;
wire  JMA ;
wire  jmb ;
wire  JMB ;
wire  jmc ;
wire  JMC ;
wire  jmd ;
wire  JMD ;
wire  jme ;
wire  JME ;
wire  jmf ;
wire  JMF ;
wire  jmg ;
wire  JMG ;
wire  jmh ;
wire  JMH ;
wire  jmi ;
wire  JMI ;
wire  jna ;
wire  JNA ;
wire  jnb ;
wire  JNB ;
wire  jnc ;
wire  JNC ;
wire  jnd ;
wire  JND ;
wire  jne ;
wire  JNE ;
wire  jnf ;
wire  JNF ;
wire  jng ;
wire  JNG ;
wire  jnh ;
wire  JNH ;
wire  jni ;
wire  JNI ;
wire  jqc ;
wire  JQC ;
wire  kaa ;
wire  kab ;
wire  kac ;
wire  kad ;
wire  kae ;
wire  kaf ;
wire  kag ;
wire  kah ;
wire  kai ;
wire  kaj ;
wire  kak ;
wire  kal ;
wire  kam ;
wire  kan ;
wire  kao ;
wire  kap ;
wire  kba ;
wire  kbb ;
wire  kbc ;
wire  kbd ;
wire  kbe ;
wire  kbf ;
wire  kbg ;
wire  kbh ;
wire  kbi ;
wire  kbj ;
wire  kbk ;
wire  kbl ;
wire  kbm ;
wire  kbn ;
wire  kbo ;
wire  kbp ;
wire  laa ;
wire  LAA ;
wire  lab ;
wire  LAB ;
wire  lac ;
wire  LAC ;
wire  lad ;
wire  LAD ;
wire  lae ;
wire  LAE ;
wire  laf ;
wire  LAF ;
wire  lag ;
wire  LAG ;
wire  lah ;
wire  LAH ;
wire  laq ;
wire  LAQ ;
wire  naa ;
wire  nab ;
wire  nac ;
wire  nad ;
wire  nae ;
wire  naf ;
wire  nag ;
wire  nah ;
wire  nai ;
wire  naj ;
wire  nak ;
wire  nal ;
wire  nam ;
wire  nan ;
wire  nao ;
wire  nap ;
wire  nba ;
wire  nbb ;
wire  nbc ;
wire  nbd ;
wire  nbe ;
wire  nbf ;
wire  nbg ;
wire  nbh ;
wire  nbi ;
wire  nbj ;
wire  nbk ;
wire  nbl ;
wire  nbm ;
wire  nbn ;
wire  nbo ;
wire  nbp ;
wire  oaa ;
wire  oab ;
wire  oac ;
wire  oad ;
wire  oae ;
wire  oaf ;
wire  oag ;
wire  oah ;
wire  oai ;
wire  oaj ;
wire  oak ;
wire  oal ;
wire  oam ;
wire  oan ;
wire  oao ;
wire  oap ;
wire  oba ;
wire  obb ;
wire  obc ;
wire  obd ;
wire  obe ;
wire  obf ;
wire  obg ;
wire  obh ;
wire  obi ;
wire  obj ;
wire  obk ;
wire  obl ;
wire  obm ;
wire  obn ;
wire  obo ;
wire  obp ;
wire  oca ;
wire  ocb ;
wire  occ ;
wire  ocd ;
wire  oce ;
wire  ocf ;
wire  ocg ;
wire  och ;
wire  oci ;
wire  ocj ;
wire  ock ;
wire  ocl ;
wire  oda ;
wire  odb ;
wire  odc ;
wire  odd ;
wire  ode ;
wire  odf ;
wire  odg ;
wire  odh ;
wire  odi ;
wire  odj ;
wire  odk ;
wire  odl ;
wire  oea ;
wire  oeb ;
wire  oec ;
wire  oed ;
wire  oee ;
wire  oef ;
wire  oeg ;
wire  oeh ;
wire  oei ;
wire  oej ;
wire  oek ;
wire  oel ;
wire  OEM ;
wire  ofa ;
wire  ofb ;
wire  ofc ;
wire  ofd ;
wire  ofe ;
wire  off ;
wire  ofg ;
wire  ofh ;
wire  ofi ;
wire  ofj ;
wire  ofk ;
wire  ofl ;
wire  oga ;
wire  ogb ;
wire  ogc ;
wire  ogd ;
wire  oge ;
wire  oha ;
wire  ohb ;
wire  ohc ;
wire  ohd ;
wire  ohe ;
wire  ohf ;
wire  ohg ;
wire  ohh ;
wire  OHI ;
wire  oja ;
wire  ojb ;
wire  ojc ;
wire  ojd ;
wire  oje ;
wire  ojf ;
wire  ojg ;
wire  ojh ;
wire  oji ;
wire  ojj ;
wire  ojk ;
wire  ojl ;
wire  ojm ;
wire  ojn ;
wire  ojo ;
wire  paa ;
wire  pab ;
wire  pac ;
wire  pad ;
wire  pae ;
wire  paf ;
wire  pag ;
wire  pah ;
wire  paj ;
wire  pak ;
wire  pal ;
wire  pam ;
wire  pan ;
wire  pao ;
wire  pap ;
wire  pba ;
wire  pbb ;
wire  pbc ;
wire  pbd ;
wire  pbe ;
wire  pbf ;
wire  pbg ;
wire  pbh ;
wire  pca ;
wire  pcb ;
wire  pcc ;
wire  pcd ;
wire  pda ;
wire  pdb ;
wire  pdc ;
wire  pdd ;
wire  pea ;
wire  peb ;
wire  pec ;
wire  ped ;
wire  pfa ;
wire  pfb ;
wire  pfc ;
wire  pfd ;
wire  qaa ;
wire  qab ;
wire  qac ;
wire  qad ;
wire  qae ;
wire  qba ;
wire  qbb ;
wire  qbc ;
wire  qbd ;
wire  qbe ;
wire  qbf ;
wire  qbg ;
wire  qbh ;
wire  QBI ;
wire  QBJ ;
wire  QBK ;
wire  qbl ;
wire  QCA ;
wire  qcb ;
wire  qcc ;
wire  QCD ;
wire  qce ;
wire  qcf ;
wire  qcg ;
wire  qci ;
wire  qcj ;
wire  qda ;
wire  qdb ;
wire  qdc ;
wire  qde ;
wire  QDF ;
wire  QDG ;
wire  QDI ;
wire  QDJ ;
wire  QDK ;
wire  QDL ;
wire  QEA ;
wire  qeb ;
wire  qei ;
wire  qej ;
wire  qek ;
wire  qel ;
wire  QFA ;
wire  qfb ;
wire  qfc ;
wire  QFD ;
wire  qfi ;
wire  QGA ;
wire  qgb ;
wire  qgc ;
wire  QHA ;
wire  qhb ;
wire  qhc ;
wire  qhd ;
wire  qhi ;
wire  QHJ ;
wire  qhk ;
wire  QHL ;
wire  QIA ;
wire  qib ;
wire  qic ;
wire  qid ;
wire  qie ;
wire  qif ;
wire  qig ;
wire  QII ;
wire  QIJ ;
wire  QIK ;
wire  QIL ;
wire  QJA ;
wire  qjb ;
wire  qjc ;
wire  qjd ;
wire  qje ;
wire  qjf ;
wire  qjg ;
wire  qjh ;
wire  qji ;
wire  QJJ ;
wire  QJK ;
wire  QJL ;
wire  QKA ;
wire  qkb ;
wire  qkc ;
wire  QKD ;
wire  QLA ;
wire  qlb ;
wire  qlc ;
wire  QMA ;
wire  qmb ;
wire  qmc ;
wire  qmd ;
wire  qme ;
wire  qmf ;
wire  qmi ;
wire  QMJ ;
wire  QMK ;
wire  QNA ;
wire  QNB ;
wire  QNC ;
wire  QND ;
wire  QNE ;
wire  qnf ;
wire  qng ;
wire  QNH ;
wire  qni ;
wire  qnj ;
wire  qnk ;
wire  qnl ;
wire  qnm ;
wire  qnn ;
wire  qno ;
wire  qnp ;
wire  QNQ ;
wire  qnr ;
wire  QOA ;
wire  QOB ;
wire  QOC ;
wire  QOD ;
wire  qqa ;
wire  qqb ;
wire  qqc ;
wire  QQD ;
wire  QQE ;
wire  QQF ;
wire  qra ;
wire  qrb ;
wire  qrc ;
wire  qrd ;
wire  qre ;
wire  qrf ;
wire  qrg ;
wire  qrh ;
wire  qri ;
wire  qrj ;
wire  qrk ;
wire  qrl ;
wire  qrm ;
wire  qrn ;
wire  qro ;
wire  qrp ;
wire  qrq ;
wire  QRR ;
wire  qsa ;
wire  qsb ;
wire  qsc ;
wire  qsd ;
wire  qsi ;
wire  qsj ;
wire  qsk ;
wire  qsl ;
wire  qsm ;
wire  qsn ;
wire  qso ;
wire  qsp ;
wire  qsq ;
wire  qta ;
wire  qtb ;
wire  qtc ;
wire  qua ;
wire  qub ;
wire  quc ;
wire  qva ;
wire  qvb ;
wire  qvc ;
wire  raa ;
wire  rab ;
wire  rac ;
wire  rad ;
wire  rae ;
wire  raf ;
wire  rag ;
wire  rah ;
wire  rai ;
wire  raj ;
wire  rak ;
wire  ral ;
wire  ram ;
wire  ran ;
wire  rao ;
wire  rap ;
wire  rba ;
wire  rbb ;
wire  rbc ;
wire  rbd ;
wire  rbe ;
wire  rbf ;
wire  rbg ;
wire  rbh ;
wire  RBI ;
wire  RBJ ;
wire  RBK ;
wire  RBL ;
wire  RBM ;
wire  rca ;
wire  rcb ;
wire  rcc ;
wire  rcd ;
wire  rce ;
wire  rcf ;
wire  rcg ;
wire  rch ;
wire  rda ;
wire  rdb ;
wire  rdc ;
wire  rdd ;
wire  rde ;
wire  rdf ;
wire  rdg ;
wire  rdh ;
wire  rea ;
wire  red ;
wire  ree ;
wire  regg ;
wire  rfa ;
wire  rfd ;
wire  rfe ;
wire  rfg ;
wire  rga ;
wire  rgd ;
wire  rge ;
wire  rgg ;
wire  rha ;
wire  rhd ;
wire  ria ;
wire  rid ;
wire  taa ;
wire  taa ;
wire  TAA ;
wire  tab ;
wire  tab ;
wire  TAB ;
wire  tac ;
wire  tac ;
wire  TAC ;
wire  tad ;
wire  TAD ;
wire  TAE ;
wire  TAF ;
wire  TAG ;
wire  tah ;
wire  TAH ;
wire  tai ;
wire  TAI ;
wire  taj ;
wire  TAJ ;
wire  tba ;
wire  TBA ;
wire  tbb ;
wire  TBB ;
wire  tbc ;
wire  TBC ;
wire  tbd ;
wire  TBD ;
wire  tca ;
wire  TCA ;
wire  tcb ;
wire  TCB ;
wire  tcc ;
wire  TCC ;
wire  tcd ;
wire  TCD ;
wire  tda ;
wire  TDA ;
wire  tdb ;
wire  TDB ;
wire  tdc ;
wire  TDC ;
wire  tdd ;
wire  TDD ;
wire  tea ;
wire  TEA ;
wire  teb ;
wire  TEB ;
wire  tec ;
wire  TEC ;
wire  ted ;
wire  TED ;
wire  tee ;
wire  TEE ;
wire  tef ;
wire  TEF ;
wire  teg ;
wire  TEG ;
wire  tfa ;
wire  TFA ;
wire  tfb ;
wire  TFB ;
wire  tga ;
wire  TGA ;
wire  tgb ;
wire  TGB ;
wire  tja ;
wire  TJA ;
wire  tjb ;
wire  TJB ;
wire  tjc ;
wire  TJC ;
wire  tjd ;
wire  TJD ;
wire  tje ;
wire  TJE ;
wire  tjf ;
wire  TJF ;
wire  tka ;
wire  TKA ;
wire  tkb ;
wire  TKB ;
wire  tkc ;
wire  TKC ;
wire  tkd ;
wire  TKD ;
wire  tke ;
wire  TKE ;
wire  tkf ;
wire  TKF ;
wire  tle ;
wire  TLE ;
wire  tlf ;
wire  TLF ;
wire  uaa ;
wire  UAA ;
wire  uab ;
wire  UAB ;
wire  uac ;
wire  UAC ;
wire  uad ;
wire  UAD ;
wire  uae ;
wire  UAE ;
wire  uaf ;
wire  UAF ;
wire  uag ;
wire  UAG ;
wire  uah ;
wire  UAH ;
wire  vaa ;
wire  vab ;
wire  vac ;
wire  vad ;
wire  vae ;
wire  vaf ;
wire  vag ;
wire  vah ;
wire  vba ;
wire  vbb ;
wire  vbc ;
wire  vbd ;
wire  vbe ;
wire  vbf ;
wire  vbg ;
wire  vbh ;
wire  ZZI ;
wire  zzo ;
wire  zzo ;
wire  zzo ;
wire  zzo ;
wire  zzo ;
wire  zzo ;
wire  zzo ;
wire  zzo ;
wire  ZZO ;
wire  ZZO ;
wire  ZZO ;
wire  ZZO ;
wire  ZZO ;
wire  ZZO ;
wire  ZZO ;
wire  ZZO ;
wire  ZZO ;
assign ZZI = 1'b1;
assign ZZO = 1'b0;
assign faa =  aaa  ; 
assign FAA = ~faa;  //complement 
assign fab =  aab  ; 
assign FAB = ~fab;  //complement 
assign JHA =  AAA  ; 
assign jha = ~JHA;  //complement  
assign JHE =  AAE  ; 
assign jhe = ~JHE;  //complement 
assign BAB = ~bab;  //complement 
assign fac =  aac  ; 
assign FAC = ~fac;  //complement 
assign fad =  aad  ; 
assign FAD = ~fad;  //complement 
assign aca = ~ACA;  //complement 
assign acb = ~ACB;  //complement 
assign EAA =  aca  ; 
assign eaa = ~EAA;  //complement 
assign EAB =  ACB & bab  |  acb & BAB  ; 
assign eab = ~EAB;  //complement 
assign fae =  aae  ; 
assign FAE = ~fae;  //complement 
assign faf =  aaf  ; 
assign FAF = ~faf;  //complement 
assign aba = ~ABA;  //complement 
assign abb = ~ABB;  //complement 
assign aaa = ~AAA;  //complement 
assign aab = ~AAB;  //complement 
assign fag =  aag  ; 
assign FAG = ~fag;  //complement 
assign fah =  aah  ; 
assign FAH = ~fah;  //complement 
assign jma = caa; 
assign JMA = ~jma; //complement 
assign jna = caa; 
assign JNA = ~jna;  //complement 
assign fai =  aai  ; 
assign FAI = ~fai;  //complement 
assign faj =  aaj  ; 
assign FAJ = ~faj;  //complement 
assign vaa = ~VAA;  //complement 
assign vba = ~VBA;  //complement 
assign fak =  aak  ; 
assign FAK = ~fak;  //complement 
assign fal =  aal  ; 
assign FAL = ~fal;  //complement 
assign haa = ~HAA;  //complement 
assign hai = ~HAI;  //complement 
assign naa = ~NAA;  //complement 
assign nai = ~NAI;  //complement 
assign nba = ~NBA;  //complement 
assign nbi = ~NBI;  //complement 
assign JCA = ~HAC & ~HAB & ~HAA  ; 
assign JCB = ~HAC & ~HAB &  HAA  ; 
assign JCC = ~HAC &  HAB & ~HAA  ; 
assign JCD = ~HAC &  HAB &  HAA  ; 
assign JCE =  HAC & ~HAB & ~HAA  ; 
assign JCF =  HAC & ~HAB &  HAA ; 
assign JCG =  HAC &  HAB & ~HAA  ; 
assign JCH =  HAC &  HAB &  HAA ; 
assign JCI = ZZI ; 
assign uaa =  paf & pag & pah & paa  ; 
assign UAA = ~uaa;  //complement  
assign zzo =  ZZI  ; 
assign ZZO = ~zzo;  //complement 
assign paa = ~PAA;  //complement 
assign pba = ~PBA;  //complement 
assign raa = ~RAA;  //complement 
assign rai = ~RAI;  //complement 
assign JAA =  QAB & rap & rao  ; 
assign jaa = ~JAA;  //complement 
assign JBA =  ran & ram  ; 
assign jba = ~JBA;  //complement 
assign TAJ =  qae  ; 
assign taj = ~TAJ;  //complement 
assign qci = ~QCI;  //complement 
assign rba = ~RBA;  //complement 
assign rca = ~RCA;  //complement 
assign rda = ~RDA;  //complement 
assign rea = ~REA;  //complement 
assign taa =  QAA  |  pba & pbe  ; 
assign TAA = ~taa; //complement 
assign taa =  QAA  |  pba & pbe  ; 
assign TAE = ~tae;  //complement 
assign qaa = ~QAA;  //complement 
assign qae = ~QAE;  //complement 
assign jfa =  qac & qad & qcd & qcj & qha & qhi  ; 
assign JFA = ~jfa;  //complement  
assign GAA = ~gaa;  //complement 
assign RBI = ~rbi;  //complement 
assign laa =  qaa  |  raa  ; 
assign LAA = ~laa; //complement 
assign QCA = ~qca;  //complement 
assign QCD = ~qcd;  //complement 
assign QBI = ~qbi;  //complement 
assign QBJ = ~qbj;  //complement 
assign qcb = ~QCB;  //complement 
assign qcc = ~QCC;  //complement 
assign qce = ~QCE;  //complement 
assign qcf = ~QCF;  //complement 
assign qcj = ~QCJ;  //complement 
assign qcg = ~QCG;  //complement 
assign qbg = ~QBG;  //complement 
assign qta = ~QTA;  //complement 
assign kaa = ~KAA;  //complement 
assign tca = qic; 
assign TCA = ~tca; //complement 
assign tcb = qic; 
assign TCB = ~tcb;  //complement 
assign tcd = qic; 
assign TCD = ~tcd;  //complement 
assign tcc = qic; 
assign TCC = ~tcc;  //complement 
assign dba = ~DBA;  //complement 
assign dca = ~DCA;  //complement 
assign oaa = ~OAA;  //complement 
assign kai = ~KAI;  //complement 
assign pca = ~PCA;  //complement 
assign pda = ~PDA;  //complement 
assign oai = ~OAI;  //complement 
assign kba = ~KBA;  //complement 
assign EBA =  KBI & PFA  |  KBA & PFB  |  KAI & PFC  |  KAA & PFD  ; 
assign eba = ~EBA;  //complement 
assign caa = ~CAA;  //complement 
assign cba = ~CBA;  //complement 
assign oba = ~OBA;  //complement 
assign kbi = ~KBI;  //complement 
assign jda =  qbj & qnb  ; 
assign JDA = ~jda;  //complement 
assign TKD =  PCA & QNQ  ; 
assign tkd = ~TKD;  //complement 
assign tba =  qqa & qlc  ; 
assign TBA = ~tba;  //complement 
assign tda =  qkc  ; 
assign TDA = ~tda;  //complement 
assign obi = ~OBI;  //complement 
assign GBA = ~gba;  //complement 
assign GBB = ~gbb;  //complement 
assign JEA =  GBA  |  GBB  |  GBC & QDE  |  GBD & qde  ; 
assign jea = ~JEA;  //complement 
assign QDI = ~qdi;  //complement 
assign ofa = ~OFA;  //complement 
assign oha = ~OHA;  //complement 
assign ojd = ~OJD;  //complement 
assign oje = ~OJE;  //complement 
assign QBK = ~qbk;  //complement 
assign qde = ~QDE;  //complement 
assign oee = ~OEE;  //complement 
assign oef = ~OEF;  //complement 
assign oeg = ~OEG;  //complement 
assign oeh = ~OEH;  //complement 
assign rfa = ~RFA;  //complement 
assign rga = ~RGA;  //complement 
assign rha = ~RHA;  //complement 
assign ria = ~RIA;  //complement 
assign oda = ~ODA;  //complement 
assign odb = ~ODB;  //complement 
assign odc = ~ODC;  //complement 
assign odd = ~ODD;  //complement 
assign oei = ~OEI;  //complement 
assign QOA = ~qoa;  //complement 
assign QOB = ~qob;  //complement 
assign oca = ~OCA;  //complement 
assign oci = ~OCI;  //complement 
assign fba =  aaa  ; 
assign FBA = ~fba;  //complement 
assign fbb =  aab  ; 
assign FBB = ~fbb;  //complement 
assign JHB =  AAA & AAB  ; 
assign jhb = ~JHB;  //complement  
assign JHF =  AAE & AAF  ; 
assign jhf = ~JHF;  //complement 
assign BAC = ~bac;  //complement 
assign BAD = ~bad;  //complement 
assign fbc =  aac  ; 
assign FBC = ~fbc;  //complement 
assign fbd =  aad  ; 
assign FBD = ~fbd;  //complement 
assign acc = ~ACC;  //complement 
assign acd = ~ACD;  //complement 
assign EAC =  ACC & bac  |  acc & BAC  ; 
assign eac = ~EAC;  //complement 
assign EAD =  ACD & bad  |  acd & BAD  ; 
assign ead = ~EAD;  //complement 
assign fbe =  aae  ; 
assign FBE = ~fbe;  //complement 
assign fbf =  aaf  ; 
assign FBF = ~fbf;  //complement 
assign abc = ~ABC;  //complement 
assign abd = ~ABD;  //complement 
assign aac = ~AAC;  //complement 
assign aad = ~AAD;  //complement 
assign fbg =  aag  ; 
assign FBG = ~fbg;  //complement 
assign fbh =  aah  ; 
assign FBH = ~fbh;  //complement 
assign jmb = cab; 
assign JMB = ~jmb; //complement 
assign jnb = cab; 
assign JNB = ~jnb;  //complement 
assign fbi =  aai  ; 
assign FBI = ~fbi;  //complement 
assign fbj =  aaj  ; 
assign FBJ = ~fbj;  //complement 
assign vab = ~VAB;  //complement 
assign vbb = ~VBB;  //complement 
assign fbk =  aak  ; 
assign FBK = ~fbk;  //complement 
assign fbl =  aal  ; 
assign FBL = ~fbl;  //complement 
assign hab = ~HAB;  //complement 
assign haj = ~HAJ;  //complement 
assign nab = ~NAB;  //complement 
assign naj = ~NAJ;  //complement 
assign nbb = ~NBB;  //complement 
assign nbj = ~NBJ;  //complement 
assign uab =  pag & pah & paa & pab  ; 
assign UAB = ~uab;  //complement  
assign zzo =  ; 
assign ZZO = ~zzo;  //complement 
assign pab = ~PAB;  //complement 
assign paj = ~PAJ;  //complement 
assign pbb = ~PBB;  //complement 
assign rab = ~RAB;  //complement 
assign raj = ~RAJ;  //complement 
assign JAB =  QAB & rap & RAO  ; 
assign jab = ~JAB;  //complement 
assign JBB =  ran & RAM  ; 
assign jbb = ~JBB;  //complement 
assign rbb = ~RBB;  //complement 
assign rcb = ~RCB;  //complement 
assign rdb = ~RDB;  //complement 
assign tab =  QAA  |  pbb & pbf  ; 
assign TAB = ~tab; //complement 
assign tab =  QAA  |  pbb & pbf  ; 
assign TAF = ~taf;  //complement 
assign qab = ~QAB;  //complement 
assign jfb =  qea & qja & qji & qka & qmi & qbe  ; 
assign JFB = ~jfb;  //complement  
assign jfc =  qac & qad & qkd  ; 
assign JFC = ~jfc;  //complement 
assign GAB = ~gab;  //complement 
assign QKD = ~qkd;  //complement 
assign RBJ = ~rbj;  //complement 
assign RBM = ~rbm;  //complement 
assign lab =  qaa  |  rab  ; 
assign LAB = ~lab; //complement 
assign QEA = ~qea;  //complement 
assign QHA = ~qha;  //complement 
assign JGA = ~rbk & ~rbj & ~rbi & QEA & rbg ; 
assign JGB = ~rbk & ~rbj &  rbi & QEA & rbg ; 
assign JGC = ~rbk &  rbj & ~rbi & QEA & rbg ; 
assign JGD = ~rbk &  rbj &  rbi & QEA & rbg ; 
assign JGE =  rbk & ~rbj & ~rbi & QEA & rbg ; 
assign JGF =  rbk & ~rbj &  rbi & QEA & rbg ; 
assign JGG =  rbk &  rbj & ~rbi & QEA & rbg ; 
assign JGH =  rbk &  rbj &  rbi & QEA & rbg ; 
assign JGI = ZZI ; 
assign qeb = ~QEB;  //complement 
assign QHJ = ~qhj;  //complement 
assign qhi = ~QHI;  //complement 
assign qhk = ~QHK;  //complement 
assign qhb = ~QHB;  //complement 
assign qhc = ~QHC;  //complement 
assign qhd = ~QHD;  //complement 
assign QHL = ~qhl;  //complement 
assign qtb = ~QTB;  //complement 
assign qtc = ~QTC;  //complement 
assign kab = ~KAB;  //complement 
assign ocb = ~OCB;  //complement 
assign ocj = ~OCJ;  //complement 
assign dbb = ~DBB;  //complement 
assign dcb = ~DCB;  //complement 
assign oab = ~OAB;  //complement 
assign kaj = ~KAJ;  //complement 
assign pcb = ~PCB;  //complement 
assign pdb = ~PDB;  //complement 
assign oaj = ~OAJ;  //complement 
assign kbb = ~KBB;  //complement 
assign EBB =  KBJ & PFA  |  KBB & PFB  |  KAJ & PFC  |  KAB & PFD  ; 
assign ebb = ~EBB;  //complement 
assign cab = ~CAB;  //complement 
assign cbb = ~CBB;  //complement 
assign obb = ~OBB;  //complement 
assign kbj = ~KBJ;  //complement 
assign TKC =  PCB & QNQ  ; 
assign tkc = ~TKC;  //complement 
assign tbb =  qqa  ; 
assign TBB = ~tbb;  //complement 
assign tdb =  qlc  ; 
assign TDB = ~tdb;  //complement 
assign obj = ~OBJ;  //complement 
assign JEB =  GBA & QDF  |  GBB & qdf  |  GBC & QDG  |  GBD & qdg  ; 
assign jeb = ~JEB;  //complement 
assign QDJ = ~qdj;  //complement 
assign ofb = ~OFB;  //complement 
assign ohb = ~OHB;  //complement 
assign ojf = ~OJF;  //complement 
assign ojg = ~OJG;  //complement 
assign JGJ =  QEA & GCG & gcf  ; 
assign jgj = ~JGJ;  //complement 
assign JGK =  QEA & GCG & GCF  ; 
assign jgk = ~JGK;  //complement 
assign QDF = ~qdf;  //complement 
assign QDG = ~qdg;  //complement 
assign oea = ~OEA;  //complement 
assign oeb = ~OEB;  //complement 
assign oec = ~OEC;  //complement 
assign oed = ~OED;  //complement 
assign qei = ~QEI;  //complement 
assign qej = ~QEJ;  //complement 
assign qek = ~QEK;  //complement 
assign qel = ~QEL;  //complement 
assign oej = ~OEJ;  //complement 
assign QOC = ~qoc;  //complement 
assign QOD = ~qod;  //complement 
assign fca =  aaa  ; 
assign FCA = ~fca;  //complement 
assign fcb =  aab  ; 
assign FCB = ~fcb;  //complement 
assign JHC =  AAA & AAB & AAC  ; 
assign jhc = ~JHC;  //complement  
assign JHG =  AAE & AAF & AAG  ; 
assign jhg = ~JHG;  //complement 
assign BAE = ~bae;  //complement 
assign BAF = ~baf;  //complement 
assign fcc =  aac  ; 
assign FCC = ~fcc;  //complement 
assign fcd =  aad  ; 
assign FCD = ~fcd;  //complement 
assign ace = ~ACE;  //complement 
assign acf = ~ACF;  //complement 
assign EAE =  ACE & bae  |  ace & BAE  ; 
assign eae = ~EAE;  //complement 
assign EAF =  ACF & baf  |  acf & BAF  ; 
assign eaf = ~EAF;  //complement 
assign fce =  aae  ; 
assign FCE = ~fce;  //complement 
assign fcf =  aaf  ; 
assign FCF = ~fcf;  //complement 
assign abe = ~ABE;  //complement 
assign abf = ~ABF;  //complement 
assign aae = ~AAE;  //complement 
assign aaf = ~AAF;  //complement 
assign fcg =  aag  ; 
assign FCG = ~fcg;  //complement 
assign fch =  aah  ; 
assign FCH = ~fch;  //complement 
assign jmc = cac; 
assign JMC = ~jmc; //complement 
assign jnc = cac; 
assign JNC = ~jnc;  //complement 
assign fci =  aai  ; 
assign FCI = ~fci;  //complement 
assign fcj =  aaj  ; 
assign FCJ = ~fcj;  //complement 
assign vac = ~VAC;  //complement 
assign vbc = ~VBC;  //complement 
assign qua = ~QUA;  //complement 
assign fck =  aak  ; 
assign FCK = ~fck;  //complement 
assign fcl =  aal  ; 
assign FCL = ~fcl;  //complement 
assign jib =  zza & ZZA & qjg & qme  ; 
assign JIB = ~jib;  //complement  
assign hac = ~HAC;  //complement 
assign hak = ~HAK;  //complement 
assign nac = ~NAC;  //complement 
assign nak = ~NAK;  //complement 
assign nbc = ~NBC;  //complement 
assign nbk = ~NBK;  //complement 
assign uac =  pag & paa & pab & pac  ; 
assign UAC = ~uac;  //complement  
assign zzo =  ; 
assign ZZO = ~zzo;  //complement 
assign pac = ~PAC;  //complement 
assign pak = ~PAK;  //complement 
assign pbc = ~PBC;  //complement 
assign rac = ~RAC;  //complement 
assign rak = ~RAK;  //complement 
assign JBC =  RAN & ram & ral  ; 
assign jbc = ~JBC;  //complement 
assign JAC =  QAB & RAP  ; 
assign jac = ~JAC;  //complement 
assign JAK =  RAK  ; 
assign jak = ~JAK;  //complement 
assign rbc = ~RBC;  //complement 
assign rcc = ~RCC;  //complement 
assign rdc = ~RDC;  //complement 
assign tac =  QAA  |  pbc & pbg  ; 
assign TAC = ~tac; //complement 
assign tac =  QAA  |  pbc & pbg  ; 
assign TAG = ~tag;  //complement 
assign qac = ~QAC;  //complement 
assign jfe =  qja & qjb & qjc & qjd & qje  ; 
assign JFE = ~jfe;  //complement  
assign jia =  qfc & qia & qka & qla  ; 
assign JIA = ~jia;  //complement 
assign GAC = ~gac;  //complement 
assign RBK = ~rbk;  //complement 
assign lac =  qaa  |  rac  ; 
assign LAC = ~lac; //complement 
assign QFA = ~qfa;  //complement 
assign QJA = ~qja;  //complement 
assign qjb = ~QJB;  //complement 
assign qjc = ~QJC;  //complement 
assign qjd = ~QJD;  //complement 
assign qje = ~QJE;  //complement 
assign qfb = ~QFB;  //complement 
assign qfc = ~QFC;  //complement 
assign qjf = ~QJF;  //complement 
assign qjg = ~QJG;  //complement 
assign qjh = ~QJH;  //complement 
assign qji = ~QJI;  //complement 
assign QFD = ~qfd;  //complement 
assign QJL = ~qjl;  //complement 
assign kac = ~KAC;  //complement 
assign dbc = ~DBC;  //complement 
assign dcc = ~DCC;  //complement 
assign oac = ~OAC;  //complement 
assign kak = ~KAK;  //complement 
assign pcc = ~PCC;  //complement 
assign pdc = ~PDC;  //complement 
assign oak = ~OAK;  //complement 
assign kbc = ~KBC;  //complement 
assign EBC =  KBK & PFA  |  KBC & PFB  |  KAK & PFC  |  KAC & PFD  ; 
assign ebc = ~EBC;  //complement 
assign cac = ~CAC;  //complement 
assign cbc = ~CBC;  //complement 
assign obc = ~OBC;  //complement 
assign kbk = ~KBK;  //complement 
assign TKB =  PCC & QNQ  ; 
assign tkb = ~TKB;  //complement 
assign tbc =  qqb  ; 
assign TBC = ~tbc;  //complement 
assign tdc =  qqc  ; 
assign TDC = ~tdc;  //complement 
assign obk = ~OBK;  //complement 
assign GBE = ~gbe;  //complement 
assign GBF = ~gbf;  //complement 
assign JEC =  GBA & QDI  |  GBB & QDJ  |  GBC & QDK  |  GBD & QDL  ; 
assign jec = ~JEC;  //complement 
assign QDK = ~qdk;  //complement 
assign ofc = ~OFC;  //complement 
assign ohc = ~OHC;  //complement 
assign ojh = ~OJH;  //complement 
assign oji = ~OJI;  //complement 
assign GCI = ~gci;  //complement 
assign GCJ = ~gcj;  //complement 
assign qqa = ~QQA;  //complement 
assign qqb = ~QQB;  //complement 
assign ode = ~ODE;  //complement 
assign odi = ~ODI;  //complement 
assign odj = ~ODJ;  //complement 
assign QJJ = ~qjj;  //complement 
assign QJK = ~qjk;  //complement 
assign qfi = ~QFI;  //complement 
assign qqc = ~QQC;  //complement 
assign oek = ~OEK;  //complement 
assign odl = ~ODL;  //complement 
assign occ = ~OCC;  //complement 
assign ock = ~OCK;  //complement 
assign fda =  aaa  ; 
assign FDA = ~fda;  //complement 
assign fdb =  aab  ; 
assign FDB = ~fdb;  //complement 
assign JHD =  AAA & AAB & AAC & AAD  ; 
assign jhd = ~JHD;  //complement  
assign JHH =  AAE & AAF & AAG & AAH  ; 
assign jhh = ~JHH;  //complement 
assign BAG = ~bag;  //complement 
assign BAH = ~bah;  //complement 
assign fdc =  aac  ; 
assign FDC = ~fdc;  //complement 
assign fdd =  aad  ; 
assign FDD = ~fdd;  //complement 
assign acg = ~ACG;  //complement 
assign ach = ~ACH;  //complement 
assign EAG =  ACG & bag  |  acg & BAG  ; 
assign eag = ~EAG;  //complement 
assign EAH =  ACH & bah  |  ach & BAH  ; 
assign eah = ~EAH;  //complement 
assign fde =  aae  ; 
assign FDE = ~fde;  //complement 
assign fdf =  aaf  ; 
assign FDF = ~fdf;  //complement 
assign abg = ~ABG;  //complement 
assign abh = ~ABH;  //complement 
assign aag = ~AAG;  //complement 
assign aah = ~AAH;  //complement 
assign fdg =  aag  ; 
assign FDG = ~fdg;  //complement 
assign fdh =  aah  ; 
assign FDH = ~fdh;  //complement 
assign jmd = cad; 
assign JMD = ~jmd; //complement 
assign jnd = cad; 
assign JND = ~jnd;  //complement 
assign fdi =  aai  ; 
assign FDI = ~fdi;  //complement 
assign fdj =  aaj  ; 
assign FDJ = ~fdj;  //complement 
assign vad = ~VAD;  //complement 
assign vbd = ~VBD;  //complement 
assign qub = ~QUB;  //complement 
assign fdk =  aak  ; 
assign FDK = ~fdk;  //complement 
assign fdl =  aal  ; 
assign FDL = ~fdl;  //complement 
assign JMI =  QUA & qub & quc  |  qua & QUB & quc  |  qua & qub & QUC  |  QUA & QUB & QUC  ; 
assign jmi = ~JMI; //complement 
assign had = ~HAD;  //complement 
assign hal = ~HAL;  //complement 
assign nad = ~NAD;  //complement 
assign nal = ~NAL;  //complement 
assign nbd = ~NBD;  //complement 
assign nbl = ~NBL;  //complement 
assign uad =  paa & pab & pac & pad  ; 
assign UAD = ~uad;  //complement  
assign zzo =  ; 
assign ZZO = ~zzo;  //complement 
assign pad = ~PAD;  //complement 
assign pal = ~PAL;  //complement 
assign pbd = ~PBD;  //complement 
assign rad = ~RAD;  //complement 
assign ral = ~RAL;  //complement 
assign JBD =  RAN & ram & RAL  ; 
assign jbd = ~JBD;  //complement 
assign JBG =  QBG & ran & ram  ; 
assign jbg = ~JBG;  //complement 
assign tad =  QAA  |  pbd & pbh  |  pbd  |  QAA & pbh  ; 
assign TAD = ~tad; //complement 
assign rbd = ~RBD;  //complement 
assign rcd = ~RCD;  //complement 
assign rdd = ~RDD;  //complement 
assign red = ~RED;  //complement 
assign tah =  QAA  |  pbc & pbh  ; 
assign TAH = ~tah; //complement 
assign qad = ~QAD;  //complement 
assign jfd =  qcg & qea & qfd & qjf & qmd & qnl  ; 
assign JFD = ~jfd;  //complement  
assign GAD = ~gad;  //complement 
assign RBL = ~rbl;  //complement 
assign lad =  qaa  |  rad  ; 
assign LAD = ~lad; //complement 
assign QGA = ~qga;  //complement 
assign QIA = ~qia;  //complement 
assign qie = ~QIE;  //complement 
assign qif = ~QIF;  //complement 
assign qig = ~QIG;  //complement 
assign qgb = ~QGB;  //complement 
assign qgc = ~QGC;  //complement 
assign qib = ~QIB;  //complement 
assign qid = ~QID;  //complement 
assign kad = ~KAD;  //complement 
assign qic = ~QIC;  //complement 
assign dbd = ~DBD;  //complement 
assign dcd = ~DCD;  //complement 
assign oad = ~OAD;  //complement 
assign kal = ~KAL;  //complement 
assign pcd = ~PCD;  //complement 
assign pdd = ~PDD;  //complement 
assign oal = ~OAL;  //complement 
assign kbd = ~KBD;  //complement 
assign EBD =  KBL & PFA  |  KBD & PFB  |  KAL & PFC  |  KAD & PFD  ; 
assign ebd = ~EBD;  //complement 
assign cad = ~CAD;  //complement 
assign cbd = ~CBD;  //complement 
assign obd = ~OBD;  //complement 
assign kbl = ~KBL;  //complement 
assign TKA =  PCD & QNQ  ; 
assign tka = ~TKA;  //complement 
assign tbd =  qqb  ; 
assign TBD = ~tbd;  //complement 
assign tdd =  qqc  ; 
assign TDD = ~tdd;  //complement 
assign obl = ~OBL;  //complement 
assign GBG = ~gbg;  //complement 
assign GBH = ~gbh;  //complement 
assign JED =  GBA & qdi  |  GBB & qdj  |  GBC & qdk  |  GBD & qdl  ; 
assign jed = ~JED;  //complement 
assign QDL = ~qdl;  //complement 
assign ofd = ~OFD;  //complement 
assign ohd = ~OHD;  //complement 
assign ojj = ~OJJ;  //complement 
assign ojk = ~OJK;  //complement 
assign TJA = QIF; 
assign tja = ~TJA; //complement 
assign TJB = QIF; 
assign tjb = ~TJB;  //complement 
assign rfd = ~RFD;  //complement 
assign rgd = ~RGD;  //complement 
assign rhd = ~RHD;  //complement 
assign rid = ~RID;  //complement 
assign oja = ~OJA;  //complement 
assign odf = ~ODF;  //complement 
assign QII = ~qii;  //complement 
assign QIJ = ~qij;  //complement 
assign QIK = ~qik;  //complement 
assign QIL = ~qil;  //complement 
assign ojb = ~OJB;  //complement 
assign oel = ~OEL;  //complement 
assign ojc = ~OJC;  //complement 
assign ocd = ~OCD;  //complement 
assign ocl = ~OCL;  //complement 
assign fea =  aba  ; 
assign FEA = ~fea;  //complement 
assign feb =  abb  ; 
assign FEB = ~feb;  //complement 
assign JHI =  AAI  ; 
assign jhi = ~JHI;  //complement  
assign BAI = ~bai;  //complement 
assign BAJ = ~baj;  //complement 
assign fec =  abc  ; 
assign FEC = ~fec;  //complement 
assign fed =  abd  ; 
assign FED = ~fed;  //complement 
assign aci = ~ACI;  //complement 
assign acj = ~ACJ;  //complement 
assign EAI =  ACI & bai  |  aci & BAI  ; 
assign eai = ~EAI;  //complement 
assign EAJ =  ACJ & baj  |  acj & BAJ  ; 
assign eaj = ~EAJ;  //complement 
assign fee =  abe  ; 
assign FEE = ~fee;  //complement 
assign fef =  abf  ; 
assign FEF = ~fef;  //complement 
assign abi = ~ABI;  //complement 
assign abj = ~ABJ;  //complement 
assign aai = ~AAI;  //complement 
assign aaj = ~AAJ;  //complement 
assign feg =  abg  ; 
assign FEG = ~feg;  //complement 
assign feh =  abh  ; 
assign FEH = ~feh;  //complement 
assign jme = cae; 
assign JME = ~jme; //complement 
assign jne = cae; 
assign JNE = ~jne;  //complement 
assign TEB =  QBB & qba  ; 
assign teb = ~TEB;  //complement 
assign TEE =  QBC & qba  ; 
assign tee = ~TEE;  //complement 
assign fei =  abi  ; 
assign FEI = ~fei;  //complement 
assign fej =  abj  ; 
assign FEJ = ~fej;  //complement 
assign vae = ~VAE;  //complement 
assign vbe = ~VBE;  //complement 
assign TEA = qba & qbb ; 
assign tea = ~TEA ; //complement 
assign tec = qba & qba ; 
assign TEC = ~tec ;  //complement 
assign TED = qba & qbc ; 
assign ted = ~TED ;  //complement 
assign tef = qba & qba; 
assign TEF = ~tef; 
assign fek =  abk  ; 
assign FEK = ~fek;  //complement 
assign fel =  abl  ; 
assign FEL = ~fel;  //complement 
assign hae = ~HAE;  //complement 
assign ham = ~HAM;  //complement 
assign nae = ~NAE;  //complement 
assign nam = ~NAM;  //complement 
assign nbe = ~NBE;  //complement 
assign nbm = ~NBM;  //complement 
assign TGA = QCI & gci ; 
assign tga = ~TGA ; //complement 
assign TGB = QCI & GCI ; 
assign tgb = ~TGB ;  //complement 
assign TEG = QBA; 
assign teg = ~TEG;  //complement 
assign uae =  pab & pac & pad & pae  ; 
assign UAE = ~uae;  //complement  
assign zzo =  ; 
assign ZZO = ~zzo;  //complement 
assign pae = ~PAE;  //complement 
assign pam = ~PAM;  //complement 
assign pbe = ~PBE;  //complement 
assign rae = ~RAE;  //complement 
assign ram = ~RAM;  //complement 
assign JBE =  RAN & RAM & rak  ; 
assign jbe = ~JBE;  //complement 
assign rbe = ~RBE;  //complement 
assign rce = ~RCE;  //complement 
assign rde = ~RDE;  //complement 
assign ree = ~REE;  //complement 
assign qbb = ~QBB;  //complement 
assign qbc = ~QBC;  //complement 
assign qba = ~QBA;  //complement 
assign GAE = ~gae;  //complement 
assign rfe = ~RFE;  //complement 
assign rge = ~RGE;  //complement 
assign lae =  qaa  |  rae  ; 
assign LAE = ~lae; //complement 
assign QKA = ~qka;  //complement 
assign QLA = ~qla;  //complement 
assign jfj =  qkb & qlb  ; 
assign JFJ = ~jfj;  //complement 
assign QQD = ~qqd;  //complement 
assign QQE = ~qqe;  //complement 
assign QQF = ~qqf;  //complement 
assign qkb = ~QKB;  //complement 
assign qkc = ~QKC;  //complement 
assign kae = ~KAE;  //complement 
assign dbe = ~DBE;  //complement 
assign dce = ~DCE;  //complement 
assign oae = ~OAE;  //complement 
assign kam = ~KAM;  //complement 
assign pea = ~PEA;  //complement 
assign pfa = ~PFA;  //complement 
assign oam = ~OAM;  //complement 
assign kbe = ~KBE;  //complement 
assign EBE =  KBM & PFA  |  KBE & PFB  |  KAM & PFC  |  KAE & PFD  ; 
assign ebe = ~EBE;  //complement 
assign cae = ~CAE;  //complement 
assign cbe = ~CBE;  //complement 
assign obe = ~OBE;  //complement 
assign kbm = ~KBM;  //complement 
assign TFA = QNA; 
assign tfa = ~TFA; //complement 
assign tkf = qnq; 
assign TKF = ~tkf;  //complement 
assign QNA = ~qna;  //complement 
assign QNQ = ~qnq;  //complement 
assign obm = ~OBM;  //complement 
assign qda = ~QDA;  //complement 
assign qlb = ~QLB;  //complement 
assign qlc = ~QLC;  //complement 
assign ofe = ~OFE;  //complement 
assign ohe = ~OHE;  //complement 
assign ojl = ~OJL;  //complement 
assign ojm = ~OJM;  //complement 
assign TJC = QIF; 
assign tjc = ~TJC; //complement 
assign TJD = QIF; 
assign tjd = ~TJD;  //complement 
assign TJE = QIF; 
assign tje = ~TJE;  //complement 
assign TJF = QIF; 
assign tjf = ~TJF;  //complement 
assign qsa = ~QSA;  //complement 
assign qsi = ~QSI;  //complement 
assign qsm = ~QSM;  //complement 
assign OEM = ~oem;  //complement 
assign ofj = ~OFJ;  //complement 
assign oce = ~OCE;  //complement 
assign ffa =  aba  ; 
assign FFA = ~ffa;  //complement 
assign ffb =  abb  ; 
assign FFB = ~ffb;  //complement 
assign JHJ =  AAI & AAJ  ; 
assign jhj = ~JHJ;  //complement  
assign BAK = ~bak;  //complement 
assign BAL = ~bal;  //complement 
assign ffc =  abc  ; 
assign FFC = ~ffc;  //complement 
assign ffd =  abd  ; 
assign FFD = ~ffd;  //complement 
assign ack = ~ACK;  //complement 
assign acl = ~ACL;  //complement 
assign EAK =  ACK & bak  |  ack & BAK  ; 
assign eak = ~EAK;  //complement 
assign EAL =  ACL & bal  |  acl & BAL  ; 
assign eal = ~EAL;  //complement 
assign ffe =  abe  ; 
assign FFE = ~ffe;  //complement 
assign fff =  abf  ; 
assign FFF = ~fff;  //complement 
assign abk = ~ABK;  //complement 
assign abl = ~ABL;  //complement 
assign aak = ~AAK;  //complement 
assign aal = ~AAL;  //complement 
assign ffg =  abg  ; 
assign FFG = ~ffg;  //complement 
assign ffh =  abh  ; 
assign FFH = ~ffh;  //complement 
assign jmf = caf; 
assign JMF = ~jmf; //complement 
assign jnf = caf; 
assign JNF = ~jnf;  //complement 
assign GBC = ~gbc;  //complement 
assign GBD = ~gbd;  //complement 
assign ffi =  abi  ; 
assign FFI = ~ffi;  //complement 
assign ffj =  abj  ; 
assign FFJ = ~ffj;  //complement 
assign vaf = ~VAF;  //complement 
assign vbf = ~VBF;  //complement 
assign quc = ~QUC;  //complement 
assign ffk =  abk  ; 
assign FFK = ~ffk;  //complement 
assign ffl =  abl  ; 
assign FFL = ~ffl;  //complement 
assign haf = ~HAF;  //complement 
assign han = ~HAN;  //complement 
assign naf = ~NAF;  //complement 
assign nan = ~NAN;  //complement 
assign nbf = ~NBF;  //complement 
assign nbn = ~NBN;  //complement 
assign uaf =  pac & pad & pae & paf  ; 
assign UAF = ~uaf;  //complement  
assign zzo =  ; 
assign ZZO = ~zzo;  //complement 
assign paf = ~PAF;  //complement 
assign pan = ~PAN;  //complement 
assign pbf = ~PBF;  //complement 
assign raf = ~RAF;  //complement 
assign ran = ~RAN;  //complement 
assign JBF =  RAN & RAM & RAK  ; 
assign jbf = ~JBF;  //complement 
assign rbf = ~RBF;  //complement 
assign rcf = ~RCF;  //complement 
assign rdf = ~RDF;  //complement 
assign GAF = ~gaf;  //complement 
assign GCF = ~gcf;  //complement 
assign laf =  qaa  |  raf  ; 
assign LAF = ~laf; //complement 
assign QMA = ~qma;  //complement 
assign qmi = ~QMI;  //complement 
assign qmb = ~QMB;  //complement 
assign qmc = ~QMC;  //complement 
assign qmd = ~QMD;  //complement 
assign qme = ~QME;  //complement 
assign qmf = ~QMF;  //complement 
assign kaf = ~KAF;  //complement 
assign dbf = ~DBF;  //complement 
assign dcf = ~DCF;  //complement 
assign oaf = ~OAF;  //complement 
assign kan = ~KAN;  //complement 
assign peb = ~PEB;  //complement 
assign pfb = ~PFB;  //complement 
assign oan = ~OAN;  //complement 
assign kbf = ~KBF;  //complement 
assign EBF =  KBN & PFA  |  KBF & PFB  |  KAN & PFC  |  KAF & PFD  ; 
assign ebf = ~EBF;  //complement 
assign caf = ~CAF;  //complement 
assign cbf = ~CBF;  //complement 
assign obf = ~OBF;  //complement 
assign kbn = ~KBN;  //complement 
assign tfb = qnh & qig ; 
assign TFB = ~tfb ; //complement 
assign tlf = qnh & qig ; 
assign TLF = ~tlf ;  //complement 
assign obn = ~OBN;  //complement 
assign qva = ~QVA;  //complement 
assign off = ~OFF;  //complement 
assign ohf = ~OHF;  //complement 
assign ojn = ~OJN;  //complement 
assign ojo = ~OJO;  //complement 
assign QNB = ~qnb;  //complement 
assign QNH = ~qnh;  //complement 
assign qsb = ~QSB;  //complement 
assign qsj = ~QSJ;  //complement 
assign QMJ = ~qmj;  //complement 
assign QMK = ~qmk;  //complement 
assign qsn = ~QSN;  //complement 
assign ofi = ~OFI;  //complement 
assign qbh = ~QBH;  //complement 
assign odg = ~ODG;  //complement 
assign odh = ~ODH;  //complement 
assign ocf = ~OCF;  //complement 
assign fga =  aba  ; 
assign FGA = ~fga;  //complement 
assign fgb =  abb  ; 
assign FGB = ~fgb;  //complement 
assign JHK =  AAI & AAJ & AAK  ; 
assign jhk = ~JHK;  //complement  
assign fgc =  abc  ; 
assign FGC = ~fgc;  //complement 
assign fgd =  abd  ; 
assign FGD = ~fgd;  //complement 
assign fge =  abe  ; 
assign FGE = ~fge;  //complement 
assign fgf =  abf  ; 
assign FGF = ~fgf;  //complement 
assign fgg =  abg  ; 
assign FGG = ~fgg;  //complement 
assign fgh =  abh  ; 
assign FGH = ~fgh;  //complement 
assign jmg = cag; 
assign JMG = ~jmg; //complement 
assign jng = cag; 
assign JNG = ~jng;  //complement 
assign fgi =  abi  ; 
assign FGI = ~fgi;  //complement 
assign fgj =  abj  ; 
assign FGJ = ~fgj;  //complement 
assign vag = ~VAG;  //complement 
assign vbg = ~VBG;  //complement 
assign fgk =  abk  ; 
assign FGK = ~fgk;  //complement 
assign fgl =  abl  ; 
assign FGL = ~fgl;  //complement 
assign hag = ~HAG;  //complement 
assign hao = ~HAO;  //complement 
assign nag = ~NAG;  //complement 
assign nao = ~NAO;  //complement 
assign nbg = ~NBG;  //complement 
assign nbo = ~NBO;  //complement 
assign uag =  pad & pae & paf & pag  ; 
assign UAG = ~uag;  //complement  
assign zzo =  ; 
assign ZZO = ~zzo;  //complement 
assign pag = ~PAG;  //complement 
assign pao = ~PAO;  //complement 
assign pbg = ~PBG;  //complement 
assign rag = ~RAG;  //complement 
assign rao = ~RAO;  //complement 
assign rbg = ~RBG;  //complement 
assign rcg = ~RCG;  //complement 
assign rdg = ~RDG;  //complement 
assign regg = ~REG;  //complement 
assign tai =  QAE  ; 
assign TAI = ~tai;  //complement 
assign GAG = ~gag;  //complement 
assign GCG = ~gcg;  //complement 
assign rfg = ~RFG;  //complement 
assign rgg = ~RGG;  //complement 
assign lag =  qaa  |  rag  ; 
assign LAG = ~lag; //complement 
assign qbe = ~QBE;  //complement 
assign kag = ~KAG;  //complement 
assign dbg = ~DBG;  //complement 
assign dcg = ~DCG;  //complement 
assign oag = ~OAG;  //complement 
assign kao = ~KAO;  //complement 
assign pec = ~PEC;  //complement 
assign pfc = ~PFC;  //complement 
assign oao = ~OAO;  //complement 
assign kbg = ~KBG;  //complement 
assign EBG =  KBO & PFA  |  KBG & PFB  |  KAO & PFC  |  KAG & PFD  ; 
assign ebg = ~EBG;  //complement 
assign cag = ~CAG;  //complement 
assign cbg = ~CBG;  //complement 
assign obg = ~OBG;  //complement 
assign kbo = ~KBO;  //complement 
assign obo = ~OBO;  //complement 
assign qvb = ~QVB;  //complement 
assign JQC =  QSQ & QSC  ; 
assign jqc = ~JQC;  //complement 
assign ofg = ~OFG;  //complement 
assign ohg = ~OHG;  //complement 
assign qsq = ~QSQ;  //complement 
assign QNC = ~qnc;  //complement 
assign qsc = ~QSC;  //complement 
assign qsk = ~QSK;  //complement 
assign qbf = ~QBF;  //complement 
assign qbl = ~QBL;  //complement 
assign qnr = ~QNR;  //complement 
assign qsp = ~QSP;  //complement 
assign odk = ~ODK;  //complement 
assign oge = ~OGE;  //complement 
assign qbd = ~QBD;  //complement 
assign qso = ~QSO;  //complement 
assign oga = ~OGA;  //complement 
assign ogb = ~OGB;  //complement 
assign ogc = ~OGC;  //complement 
assign ogd = ~OGD;  //complement 
assign ocg = ~OCG;  //complement 
assign fha =  aba  ; 
assign FHA = ~fha;  //complement 
assign fhb =  abb  ; 
assign FHB = ~fhb;  //complement 
assign fhc =  abc  ; 
assign FHC = ~fhc;  //complement 
assign fhd =  abd  ; 
assign FHD = ~fhd;  //complement 
assign fhe =  abe  ; 
assign FHE = ~fhe;  //complement 
assign fhf =  abf  ; 
assign FHF = ~fhf;  //complement 
assign fhg =  abg  ; 
assign FHG = ~fhg;  //complement 
assign fhh =  abh  ; 
assign FHH = ~fhh;  //complement 
assign jmh = cah; 
assign JMH = ~jmh; //complement 
assign jnh = cah; 
assign JNH = ~jnh;  //complement 
assign fhi =  abi  ; 
assign FHI = ~fhi;  //complement 
assign fhj =  abj  ; 
assign FHJ = ~fhj;  //complement 
assign vah = ~VAH;  //complement 
assign vbh = ~VBH;  //complement 
assign qra = ~QRA;  //complement 
assign qrb = ~QRB;  //complement 
assign qrc = ~QRC;  //complement 
assign qrd = ~QRD;  //complement 
assign fhk =  abk  ; 
assign FHK = ~fhk;  //complement 
assign fhl =  abl  ; 
assign FHL = ~fhl;  //complement 
assign qre = ~QRE;  //complement 
assign qrf = ~QRF;  //complement 
assign qrg = ~QRG;  //complement 
assign qrh = ~QRH;  //complement 
assign qri = ~QRI;  //complement 
assign qrj = ~QRJ;  //complement 
assign qrk = ~QRK;  //complement 
assign qrl = ~QRL;  //complement 
assign qrm = ~QRM;  //complement 
assign qrn = ~QRN;  //complement 
assign qro = ~QRO;  //complement 
assign hah = ~HAH;  //complement 
assign nah = ~NAH;  //complement 
assign nap = ~NAP;  //complement 
assign nbh = ~NBH;  //complement 
assign nbp = ~NBP;  //complement 
assign QRR = ~qrr;  //complement 
assign uah =  pae & paf & pag & pah  ; 
assign UAH = ~uah;  //complement  
assign zzo =  ; 
assign ZZO = ~zzo;  //complement 
assign pah = ~PAH;  //complement 
assign pap = ~PAP;  //complement 
assign pbh = ~PBH;  //complement 
assign rah = ~RAH;  //complement 
assign rap = ~RAP;  //complement 
assign rbh = ~RBH;  //complement 
assign rch = ~RCH;  //complement 
assign rdh = ~RDH;  //complement 
assign LAQ =  QAE & RAQ  ; 
assign laq = ~LAQ;  //complement 
assign GAH = ~gah;  //complement 
assign GAI = ~gai;  //complement 
assign lah =  qaa  |  rah  ; 
assign LAH = ~lah; //complement 
assign qnm = ~QNM;  //complement 
assign qnn = ~QNN;  //complement 
assign qno = ~QNO;  //complement 
assign qnp = ~QNP;  //complement 
assign jfg =  qre & qrf & qrg & qrh & qri  ; 
assign JFG = ~jfg;  //complement  
assign jff =  qra & qrb & qrc & qrd  ; 
assign JFF = ~jff;  //complement 
assign qni = ~QNI;  //complement 
assign qnj = ~QNJ;  //complement 
assign qnk = ~QNK;  //complement 
assign qnl = ~QNL;  //complement 
assign jfh =  qrj & qrk & qrl & qrm & qrn & qro  ; 
assign JFH = ~jfh;  //complement  
assign jfi =  qnd & qni & qnj  ; 
assign JFI = ~jfi;  //complement 
assign kah = ~KAH;  //complement 
assign qrp = ~QRP;  //complement 
assign qrq = ~QRQ;  //complement 
assign dbh = ~DBH;  //complement 
assign dch = ~DCH;  //complement 
assign oah = ~OAH;  //complement 
assign kap = ~KAP;  //complement 
assign ped = ~PED;  //complement 
assign pfd = ~PFD;  //complement 
assign oap = ~OAP;  //complement 
assign kbh = ~KBH;  //complement 
assign EBH =  KBP & PFA  |  KBH & PFB  |  KAP & PFC  |  KAH & PFD  ; 
assign ebh = ~EBH;  //complement 
assign cah = ~CAH;  //complement 
assign cbh = ~CBH;  //complement 
assign obh = ~OBH;  //complement 
assign kbp = ~KBP;  //complement 
assign tke = qnk; 
assign TKE = ~tke; //complement 
assign tle = qnk; 
assign TLE = ~tle;  //complement 
assign obp = ~OBP;  //complement 
assign qvc = ~QVC;  //complement 
assign ofl = ~OFL;  //complement 
assign qdc = ~QDC;  //complement 
assign ofh = ~OFH;  //complement 
assign ohh = ~OHH;  //complement 
assign JNI =  QVA & qvb & qvc  |  qva & QVB & qvc  |  qva & qvb & QVC  |  QVA & QVB & QVC  ; 
assign jni = ~JNI; //complement 
assign QND = ~qnd;  //complement 
assign qng = ~QNG;  //complement 
assign qsd = ~QSD;  //complement 
assign qsl = ~QSL;  //complement 
assign qnf = ~QNF;  //complement 
assign och = ~OCH;  //complement 
assign OHI = ~ohi;  //complement 
assign QNE = ~qne;  //complement 
assign ofk = ~OFK;  //complement 
assign qdb = ~QDB;  //complement 
assign iaa = ~IAA; //complement 
assign iab = ~IAB; //complement 
assign iac = ~IAC; //complement 
assign iad = ~IAD; //complement 
assign iae = ~IAE; //complement 
assign iaf = ~IAF; //complement 
assign iag = ~IAG; //complement 
assign iah = ~IAH; //complement 
assign iai = ~IAI; //complement 
assign iaj = ~IAJ; //complement 
assign iak = ~IAK; //complement 
assign ial = ~IAL; //complement 
assign iam = ~IAM; //complement 
assign ian = ~IAN; //complement 
assign iao = ~IAO; //complement 
assign iap = ~IAP; //complement 
assign iba = ~IBA; //complement 
assign ibb = ~IBB; //complement 
assign ibc = ~IBC; //complement 
assign ibd = ~IBD; //complement 
assign ibe = ~IBE; //complement 
assign ibf = ~IBF; //complement 
assign ibg = ~IBG; //complement 
assign ibh = ~IBH; //complement 
assign ibi = ~IBI; //complement 
assign ibj = ~IBJ; //complement 
assign ibk = ~IBK; //complement 
assign ibl = ~IBL; //complement 
assign ibm = ~IBM; //complement 
assign ibn = ~IBN; //complement 
assign ibo = ~IBO; //complement 
assign ibp = ~IBP; //complement 
assign ica = ~ICA; //complement 
assign icb = ~ICB; //complement 
assign icc = ~ICC; //complement 
assign icd = ~ICD; //complement 
assign ice = ~ICE; //complement 
assign ida = ~IDA; //complement 
assign idb = ~IDB; //complement 
assign idc = ~IDC; //complement 
assign ifa = ~IFA; //complement 
assign ifb = ~IFB; //complement 
assign ifc = ~IFC; //complement 
assign ifd = ~IFD; //complement 
assign ife = ~IFE; //complement 
assign ifff  = ~IFFF ; //complement 
assign ifg = ~IFG; //complement 
assign ifh = ~IFH; //complement 
assign ifi = ~IFI; //complement 
assign ifj = ~IFJ; //complement 
assign ifk = ~IFK; //complement 
assign ifl = ~IFL; //complement 
assign iga = ~IGA; //complement 
assign igb = ~IGB; //complement 
always@(posedge IZZ )
   begin 
 bab <=  jha  ; 
 ACA <= AAA ; 
 ACB <= AAB ; 
 ABA <=  ABA & TED  |  AAA & TEE  |  HAD & TEF  ; 
 ABB <=  ABB & TED  |  AAB & TEE  |  HAE & TEF  ; 
 AAA <=  AAA & TEA  |  EAA & TEB  |  HAD & TEC  ; 
 AAB <=  AAB & TEA  |  EAB & TEB  |  HAE & TEC  ; 
 VAA <=  QNG & PBA  ; 
 VBA <=  QNG & PBA  ; 
 HAA <=  RAA & TGA  |  IAA & TGB  ; 
 HAI <=  RAI & TGA  |  IAI & TGB  ; 
 NAA <= IAA ; 
 NAI <= IAI ; 
 NBA <= IBA ; 
 NBI <= IBI ; 
 PAA <=  PAA & taj & teg  |  PAH & TAJ  |  JCA & TEG  ; 
 PBA <=  PAA & taj & teg  |  PAH & TAJ  |  JCA & TEG  ; 
 RAA <=  MAA & TAA  |  MBA & TAB  |  MCA & TAC  |  MDA & TAD  |  LAA  ; 
 RAI <=  MAA & TAA  |  MBA & TAB  |  MCA & TAC  |  MDA & TAD  |  LAA  ; 
 QCI <= QCB ; 
 RBA <= RAA ; 
 RCA <= RBA ; 
 RDA <= RCA ; 
 REA <= RDA ; 
 QAA <=  JAA & JBG  |  JAC & JBB  |  JFA  |  JFB  |  QKD  ; 
 QAE <=  JAA & JBG  |  JAC & JBB  |  JFA  |  JFB  |  QKD  ; 
 gaa <= raa ; 
 rbi <= raa ; 
 qca <=  jaa  |  jba  |  QBG  ; 
 qcd <=  qcc  |  qda  ; 
 qbi <=  qib  |  RBJ  |  rba  ; 
 qbj <=  qib  |  RBJ  |  RBI  ; 
 QCB <= QCA ; 
 QCC <= QCB ; 
 QCE <= QCD ; 
 QCF <= QCE ; 
 QCJ <=  QCB  |  QCD  |  QCE  ; 
 QCG <= QCF ; 
 QBG <=  JIB  |  JIA  |  QTA  ; 
 QTA <=  JIB  |  JIA  |  QTB  ; 
 KAA <=  KAA & tka & tja  |  CBA & TKA  |  NAA & TJA  ; 
 DBA <=  DBA & qrq  |  DAA & QRQ  ; 
 DCA <=  DCA & qrq  |  DBA & QRQ  ; 
 OAA <=  RAA & TBA  |  KAA & TCA  |  RCA & TDA  ; 
 KAI <=  KAI & tkb & tjb  |  CBA & TKB  |  NAI & TJB  ; 
 PCA <=  PDA & tkf  |  PDD & TKF  |  TKE  ; 
 PDA <=  PDA & tkf  |  PDD & TKF  |  TKE  ; 
 OAI <=  RBA & TBB  |  KAI & TCB  |  RBA & TDB  ; 
 KBA <=  KBA & tkc & tjc  |  CBA & TKC  |  NBA & TJC  ; 
 CAA <=  CAA & tfa & tfb  |  DCA & TFA  |  EBA & TFB  ; 
 CBA <=  CAA & tfa & tfb  |  DCA & TFA  |  EBA & TFB  ; 
 OBA <=  RCA & TBC  |  KBA & TCC  |  RAA & TDC  ; 
 KBI <=  KBI & tkd & tjd  |  CBA & TKD  |  NBI & TJD  ; 
 OBI <=  RDA & TBD  |  KBI & TCD  |  RBA & TDD  ; 
 gba <=  GAB  |  GAA  ; 
 gbb <=  GAB  |  gaa  ; 
 qdi <=  qdi & qoa  |  ICA  |  QSP  ; 
 OFA <= CAA ; 
 OHA <= CAA ; 
 OJD <= ABA ; 
 OJE <= ABB ; 
 qbk <=  pcd  |  qnq  ; 
 QDE <=  QDE & jda & qnj  |  QBI  |  QBK  ; 
 OEE <= QEI ; 
 OEF <= QEJ ; 
 OEG <= QEK ; 
 OEH <= QEL ; 
 RFA <= REA ; 
 RGA <= RFA ; 
 RHA <= RGA ; 
 RIA <= RHA ; 
 ODA <=  RBI & QGA  |  RDA & QHC  ; 
 ODB <=  RBJ & QGA  |  RDB & QHC  ; 
 ODC <=  RDC & QHC  ; 
 ODD <=  rdc & QHC  ; 
 OEI <=  QFI & rcd  |  QFD & red  |  QII & rca  |  JFJ & rcg  ; 
 qoa <=  qhb  |  gba  ; 
 qob <=  qhb  |  gbb  ; 
 OCA <= RBA ; 
 OCI <= RCA ; 
 bac <=  jhb  ; 
 bad <=  jhc  ; 
 ACC <= AAC ; 
 ACD <= AAD ; 
 ABC <=  ABC & TED  |  AAC & TEE  |  HAF & TEF  ; 
 ABD <=  ABD & TED  |  AAD & TEE  |  HAG & TEF  ; 
 AAC <=  AAC & TEA  |  EAC & TEB  |  HAF & TEC  ; 
 AAD <=  AAD & TEA  |  EAD & TEB  |  HAG & TEC  ; 
 VAB <=  QNG & PBB  ; 
 VBB <=  QNG & PBB  ; 
 HAB <=  RAB & TGA  |  IAB & TGB  ; 
 HAJ <=  RAJ & TGA  |  IAJ & TGB  ; 
 NAB <= IAB ; 
 NAJ <= IAJ ; 
 NBB <= IBB ; 
 NBJ <= IBJ ; 
 PAB <=  PAB & taj & teg  |  PAA & TAJ  |  JCB & TEG  ; 
 PAJ <=  PAB & taj & teg  |  PAA & TAJ  |  JCB & TEG  ; 
 PBB <=  PAB & taj & teg  |  PAA & TAJ  |  JCB & TEG  ; 
 RAB <=  MAB & TAA  |  MBB & TAB  |  MCB & TAC  |  MDB & TAD  |  LAB  ; 
 RAJ <=  MAB & TAA  |  MBB & TAB  |  MCB & TAC  |  MDB & TAD  |  LAB  ; 
 RBB <= RAB ; 
 RCB <= RBB ; 
 RDB <= RCB ; 
 QAB <=  JAA & JBG  |  QCC & qda  |  JFC & qsc  ; 
 gab <= rab ; 
 qkd <= qka ; 
 rbj <= rab ; 
 rbm <= rab ; 
 qea <=  jab & jaa  |  jbc & jab  ; 
 qha <=  jaa & jaa  |  jbd & jab  ; 
 QEB <= QEA ; 
 qhj <= qhi ; 
 QHI <=  QHA  |  QHB  ; 
 QHK <=  QHC  |  QHD  ; 
 QHB <= QHA ; 
 QHC <= QHB ; 
 QHD <= QHC ; 
 qhl <= qhk ; 
 QTB <=  JIB  |  JIA  |  QTC  ; 
 QTC <=  JIB  ; 
 KAB <=  KAB & tka & tja  |  CBB & TKA  |  NAB & TJA  ; 
 OCB <= RBB ; 
 OCJ <= RCB ; 
 DBB <=  DBB & qrq  |  DAB & QRQ  ; 
 DCB <=  DCB & qrq  |  DBB & QRQ  ; 
 OAB <=  RAB & TBA  |  KAB & TCA  |  RCB & TDA  ; 
 KAJ <=  KAJ & tkb & tjb  |  CBB & TKB  |  NAJ & TJB  ; 
 PCB <=  PDB & tkf & tke  |  PDA & TKF  ; 
 PDB <=  PDB & tkf & tke  |  PDA & TKF  ; 
 OAJ <=  RBB & TBB  |  KAJ & TCB  |  RBB & TDB  ; 
 KBB <=  KBB & tkc & tjc  |  CBB & TKC  |  NBB & TJC  ; 
 CAB <=  CAB & tfa & tfb  |  DCB & TFA  |  EBB & TFB  ; 
 CBB <=  CAB & tfa & tfb  |  DCB & TFA  |  EBB & TFB  ; 
 OBB <=  RCB & TBC  |  KBB & TCC  |  RAB & TDC  ; 
 KBJ <=  KBJ & tkd & tjd  |  CBB & TKD  |  NBJ & TJD  ; 
 OBJ <=  RDB & TBD  |  KBJ & TCD  |  RBB & TDD  ; 
 qdj <=  qdj & qob  |  ICB  |  QSP  ; 
 OFB <= CAB ; 
 OHB <= CAB ; 
 OJF <= ABC ; 
 OJG <= ABD ; 
 qdf <=  IDA  |  IDB  ; 
 qdg <=  IDC  ; 
 OEA <= JGA ; 
 OEB <= JGB ; 
 OEC <= JGJ ; 
 OED <= JGK ; 
 QEI <= JGE ; 
 QEJ <= JGF ; 
 QEK <= JGG ; 
 QEL <= JGH ; 
 OEJ <=  QFI & RCD  |  QFD & RED  |  QIJ & rca  |  JFJ & RCG  ; 
 qoc <=  qhb  |  gbc  ; 
 qod <=  qhb  |  gbd  ; 
 bae <=  jhd  ; 
 baf <=  jhd  |  jhe  ; 
 ACE <= AAE ; 
 ACF <= AAF ; 
 ABE <=  ABE & TED  |  AAE & TEE  |  HAH & TEF  ; 
 ABF <=  ABF & TED  |  AAF & TEE  |  HAI & TEF  ; 
 AAE <=  AAE & TEA  |  EAE & TEB  |  HAH & TEC  ; 
 AAF <=  AAF & TEA  |  EAF & TEB  |  HAI & TEC  ; 
 VAC <=  QNG & PBC  ; 
 VBC <=  QNG & PBC  ; 
 QUA <=  JNA & jnb & jnc  |  jna & JNB & jnc  |  jna & jnb & JNC  |  JNA & JNB & JNC  ;
 HAC <=  RAC & TGA  |  IAC & TGB  ; 
 HAK <=  RAK & TGA  |  IAK & TGB  ; 
 NAC <= IAC ; 
 NAK <= IAK ; 
 NBC <= IBC ; 
 NBK <= IBK ; 
 PAC <=  PAC & taj & teg  |  PAB & TAJ  |  JCC & TEG  ; 
 PAK <=  PAC & taj & teg  |  PAB & TAJ  |  JCC & TEG  ; 
 PBC <=  PAC & taj & teg  |  PAB & TAJ  |  JCC & TEG  ; 
 RAC <=  MAC & TAA  |  MBC & TAB  |  MCC & TAC  |  MDC & TAD  |  LAC  ; 
 RAK <=  MAC & TAA  |  MBC & TAB  |  MCC & TAC  |  MDC & TAD  |  LAC  ; 
 RBC <= RAC ; 
 RCC <= RBC ; 
 RDC <= RCC ; 
 QAC <=  JAA & JBB & JAK  |  QHC  |  JAA & JBE  ; 
 gac <= rac ; 
 rbk <= rac ; 
 qfa <=  jaa  |  jbb  |  JAK  ; 
 qja <=  jaa  |  jbf  ; 
 QJB <= QJA ; 
 QJC <= QJB ; 
 QJD <= QJC ; 
 QJE <= QJD ; 
 QFB <= QFA ; 
 QFC <= QFB ; 
 QJF <= QJE ; 
 QJG <= QJF ; 
 QJH <= QJG ; 
 QJI <= JFE ; 
 qfd <=  qfc  |  rdb  ; 
 qjl <=  qjd  |  rea  ; 
 KAC <=  KAC & tka & tja  |  CBC & TKA  |  NAC & TJA  ; 
 DBC <=  DBC & qrq  |  DAC & QRQ  ; 
 DCC <=  DCC & qrq  |  DBC & QRQ  ; 
 OAC <=  RAC & TBA  |  KAC & TCA  |  RCC & TDA  ; 
 KAK <=  KAK & tkb & tjb  |  CBC & TKB  |  NAK & TJB  ; 
 PCC <=  PDC & tkf & tke  |  PDB & TKF  ; 
 PDC <=  PDC & tkf & tke  |  PDB & TKF  ; 
 OAK <=  RBC & TBB  |  KAK & TCB  |  RBC & TDB  ; 
 KBC <=  KBC & tkc & tjc  |  CBC & TKC  |  NBC & TJC  ; 
 CAC <=  CAC & tfa & tfb  |  DCC & TFA  |  EBC & TFB  ; 
 CBC <=  CAC & tfa & tfb  |  DCC & TFA  |  EBC & TFB  ; 
 OBC <=  RCC & TBC  |  KBC & TCC  |  RAC & TDC  ; 
 KBK <=  KBK & tkd & tjd  |  CBC & TKD  |  NBK & TJD  ; 
 OBK <=  RDC & TBD  |  KBK & TCD  |  RBC & TDD  ; 
 gbe <=  GAD  |  GAC  ; 
 gbf <=  GAD  |  gac  ; 
 qdk <=  qdk & qoc  |  ICC  |  QSP  ; 
 OFC <= CAC ; 
 OHC <= CAC ; 
 OJH <= ABE ; 
 OJI <= ABF ; 
 gci <=  gbb  |  gbe  ; 
 gcj <=  gbb  ; 
 QQA <=  QFI & RCA  |  QFD  |  JAB  ; 
 QQB <=  QFD & RCA  ; 
 ODE <= QGA ; 
 ODI <= QMB ; 
 ODJ <= QJD ; 
 qjj <=  qjh  |  RID  |  RIA  ; 
 qjk <=  qjh  |  rid  |  RIA  ; 
 QFI <=  QFA & rbb  ; 
 QQC <=  QFI & rca  ; 
 OEK <=  QGC & rcd  |  QJJ  |  QMJ  |  QIK & rca  ; 
 ODL <=  QHJ  |  QHL  |  QJC  |  QJE  |  QMC  ; 
 OCC <= RBC ; 
 OCK <= RCC ; 
 bag <=  jhd  |  jhf  ; 
 bah <=  jhd  |  jhg  ; 
 ACG <= AAG ; 
 ACH <= AAH ; 
 ABG <=  ABG & TED  |  AAG & TEE  |  HAJ & TEF  ; 
 ABH <=  ABH & TED  |  AAH & TEE  |  HAK & TEF  ; 
 AAG <=  AAG & TEA  |  EAG & TEB  |  HAJ & TEC  ; 
 AAH <=  AAH & TEA  |  EAH & TEB  |  HAK & TEC  ; 
 VAD <=  QNG & PBD  ; 
 VBD <=  QNG & PBD  ; 
 QUB <=  JND & jne  |  jnd & JNE  |  jnd & jne  |  JND & JNE  ;
 HAD <=  RAD & TGA  |  IAD & TGB  ; 
 HAL <=  RAL & TGA  |  IAL & TGB  ; 
 NAD <= IAD ; 
 NAL <= IAL ; 
 NBD <= IBD ; 
 NBL <= IBL ; 
 PAD <=  PAD & taj & teg  |  PAC & TAJ  |  JCD & TEG  ; 
 PAL <=  PAD & taj & teg  |  PAC & TAJ  |  JCD & TEG  ; 
 PBD <=  PAD & taj & teg  |  PAC & TAJ  |  JCD & TEG  ; 
 RAD <=  MAD & TAA  |  MBD & TAB  |  MCD & TAC  |  MDD & TAD  |  LAD  ; 
 RAL <=  MAD & TAA  |  MBD & TAB  |  MCD & TAC  |  MDD & TAD  |  LAD  ; 
 RBD <= RAD ; 
 RCD <= RBD ; 
 RDD <= RCD ; 
 RED <= RDD ; 
 QAD <=  QFB & rcb  |  QLB  |  JFD  ; 
 gad <= rad ; 
 rbl <= rad ; 
 qga <=  jaa  |  jbb  |  jak  ; 
 qia <=  jaa  |  jbe  ; 
 QIE <= QID ; 
 QIF <= QIE ; 
 QIG <= QIF ; 
 QGB <= QGA ; 
 QGC <= QGB ; 
 QIB <= QIA ; 
 QID <=  QIC & QCJ  ; 
 KAD <=  KAD & tka & tja  |  CBD & TKA  |  NAD & TJA  ; 
 QIC <= QIB ; 
 DBD <=  DBD & qrq  |  DAD & QRQ  ; 
 DCD <=  DCD & qrq  |  DBD & QRQ  ; 
 OAD <=  RAD & TBA  |  KAD & TCA  |  RCD & TDA  ; 
 KAL <=  KAL & tkb & tjb  |  CBD & TKB  |  NAL & TJB  ; 
 PCD <=  PDD & tkf & tke  |  PDC & TKF  ; 
 PDD <=  PDD & tkf & tke  |  PDC & TKF  ; 
 OAL <=  RBD & TBB  |  KAL & TCB  |  RBD & TDB  ; 
 KBD <=  KBD & tkc & tjc  |  CBD & TKC  |  NBD & TJC  ; 
 CAD <=  CAD & tfa & tfb  |  DCD & TFA  |  EBD & TFB  ; 
 CBD <=  CAD & tfa & tfb  |  DCD & TFA  |  EBD & TFB  ; 
 OBD <=  RCD & TBC  |  KBD & TCC  |  RAD & TDC  ; 
 KBL <=  KBL & tkd & tjd  |  CBD & TKD  |  NBL & TJD  ; 
 OBL <=  RDD & TBD  |  KBL & TCD  |  RBD & TDD  ; 
 gbg <=  gad  |  GAC  ; 
 gbh <=  gad  |  gac  ; 
 qdl <=  qdl & qod  |  ICD  |  QSP  ; 
 OFD <= CAD ; 
 OHD <= CAD ; 
 OJJ <= ABG ; 
 OJK <= ABH ; 
 RFD <= RED ; 
 RGD <= RFD ; 
 RHD <= RGD ; 
 RID <= RHD ; 
 OJA <=  PAJ  |  PAL  |  PAN  |  PAP  ; 
 ODF <= QIA ; 
 qii <=  qia  |  RBL  |  RBM  ; 
 qij <=  qia  |  rbl  |  RBM  ; 
 qik <=  qia  |  RBL  |  rbj  ; 
 qil <=  qia  |  rbl  |  rbj  ; 
 OJB <=  PAK  |  PAL  |  PAO  |  PAP  ; 
 OEL <=  QGC & RCD  |  QJK  |  QMK  |  QIL & rca  ; 
 OJC <=  PAM  |  PAN  |  PAO  |  PAP  ; 
 OCD <= RBD ; 
 OCL <= RCD ; 
 bai <=  jhd  |  jhh  ; 
 baj <=  jhd  |  jhh  |  jhi  ; 
 ACI <= AAI ; 
 ACJ <= AAJ ; 
 ABI <=  ABI & TED  |  AAI & TEE  |  HAL & TEF  ; 
 ABJ <=  ABJ & TED  |  AAJ & TEE  |  HAM & TEF  ; 
 AAI <=  AAI & TEA  |  EAI & TEB  |  HAH & TEC  ; 
 AAJ <=  AAJ & TEA  |  EAJ & TEB  |  HAI & TEC  ; 
 VAE <=  QNG & PBE  ; 
 VBE <=  QNG & PBE  ; 
 HAE <=  RAE & TGA  |  IAE & TGB  ; 
 HAM <=  RAM & TGA  |  IAM & TGB  ; 
 NAE <= IAE ; 
 NAM <= IAM ; 
 NBE <= IBE ; 
 NBM <= IBM ; 
 PAE <=  PAE & taj & teg  |  PAD & TAJ  |  JCE & TEG  ; 
 PAM <=  PAE & taj & teg  |  PAD & TAJ  |  JCE & TEG  ; 
 PBE <=  PAE & taj & teg  |  PAD & TAJ  |  JCE & TEG  ; 
 RAE <=  MAE & TAA  |  MBE & TAB  |  MCE & TAC  |  MDE & TAD  |  LAE  ; 
 RAM <=  MAE & TAA  |  MBE & TAB  |  MCE & TAC  |  MDE & TAD  |  LAE  ; 
 RBE <= RAE ; 
 RCE <= RBE ; 
 RDE <= RCE ; 
 REE <= RDE ; 
 QBB <=  PAD & TAI  |  QCE & uad  ; 
 QBC <=  PAH & TAI  ; 
 QBA <=  QCC & QDA  |  QBF  |  QND  ; 
 gae <= rae ; 
 RFE <= REE ; 
 RGE <= RFE ; 
 qka <=  jac  |  jba  ; 
 qla <=  jac  |  jbb  ; 
 qqd <= tai ; 
 qqe <= qqd ; 
 qqf <= qqe ; 
 QKB <= QKA ; 
 QKC <= QKB ; 
 KAE <=  KAE & tka & tja  |  CBE & TKA  |  NAE & TJA  ; 
 DBE <=  DBE & qrq  |  DAE & QRQ  ; 
 DCE <=  DCE & qrq  |  DBE & QRQ  ; 
 OAE <=  RAE & TBA  |  KAE & TCA  ; 
 KAM <=  KAM & tkb & tjb  |  CBE & TKB  |  NAM & TJB  ; 
 PEA <=  PEA & tlf  |  PED & TLF  |  TLE  ; 
 PFA <=  PEA & tlf  |  PED & TLF  |  TLE  ; 
 OAM <=  RBE & TBB  |  KAM & TCB  ; 
 KBE <=  KBE & tkc & tjc  |  CBE & TKC  |  NBE & TJC  ; 
 CAE <=  CAE & tfa & tfb  |  DCE & TFA  |  EBE & TFB  ; 
 CBE <=  CAE & tfa & tfb  |  DCE & TFA  |  EBE & TFB  ; 
 OBE <=  RCE & TBC  |  KBE & TCC  |  RAE & TDC  ; 
 KBM <=  KBM & tkd & tjf  |  CBE & TKD  |  NBM & TJF  ; 
 qna <=  QSM  |  qsi  ; 
 qnq <=  qna  |  QSK  ; 
 OBM <=  RDE & TBD  |  KBM & TCD  |  RBE & TDD  ; 
 QDA <=  JEA & GBE  |  JEB & GBF  |  JEC & GBG  |  JED & GBH  ; 
 QLB <= QLA ; 
 QLC <= QLB ; 
 OFE <= CAE ; 
 OHE <= CAE ; 
 OJL <= ABI ; 
 OJM <= ABJ ; 
 QSA <=  QSA & qrp  |  DAI & QRP  ; 
 QSI <=  QSI & qrp  |  QSA & QRP  ; 
 QSM <= QSI ; 
 oem <=  QIB & rcd  |  QJB & rcb  |  QJD & red  |  QMB & rcg  |  QMI  ; 
 OFJ <= QSI ; 
 OCE <= RBE ; 
 bak <=  jhd  |  jhh  |  jhj  ; 
 bal <=  jhd  |  jhh  |  jhk  ; 
 ACK <= AAK ; 
 ACL <= AAL ; 
 ABK <=  ABK & TED  |  AAK & TEE  |  HAN & TEF  ; 
 ABL <=  ABL & TED  |  AAL & TEE  |  HAO & TEF  ; 
 AAK <=  AAK & TEA  |  EAK & TEB  |  HAJ & TEC  ; 
 AAL <=  AAL & TEA  |  EAL & TEB  |  HAK & TEC  ; 
 gbc <=  gab  |  GAA  |  MBE  ; 
 gbd <=  gab  |  gaa  ; 
 VAF <=  QNG & PBF  ; 
 VBF <=  QNG & PBF  ; 
 QUC <=  JNF & jng & jnh  |  jnf & JNG & jnh  |  jnf & jng & JNH  |  JNF & JNG & JNH  ;
 HAF <=  RAF & TGA  |  IAF & TGB  ; 
 HAN <=  RAN & TGA  |  IAN & TGB  ; 
 NAF <= IAF ; 
 NAN <= IAN ; 
 NBF <= IBF ; 
 NBN <= IBN ; 
 PAF <=  PAF & taj & teg  |  PAE & TAJ  |  JCF & TEG  ; 
 PAN <=  PAF & taj & teg  |  PAE & TAJ  |  JCF & TEG  ; 
 PBF <=  PAF & taj & teg  |  PAE & TAJ  |  JCF & TEG  ; 
 RAF <=  MAF & TAA  |  MBF & TAB  |  MCF & TAC  |  MDF & TAD  |  LAF  ; 
 RAN <=  MAF & TAA  |  MBF & TAB  |  MCF & TAC  |  MDF & TAD  |  LAF  ; 
 RBF <= RAF ; 
 RCF <= RBF ; 
 RDF <= RCF ; 
 gaf <= raf ; 
 gcf <= raf ; 
 qma <=  jac  |  raf  ; 
 QMI <=  QMA  |  QMB  |  QMC  ; 
 QMB <= QMA ; 
 QMC <= QMB ; 
 QMD <= QMC ; 
 QME <= QMD ; 
 QMF <= QME ; 
 KAF <=  KAF & tka & tja  |  CBF & TKA  |  NAF & TJA  ; 
 DBF <=  DBF & qrq  |  DAF & QRQ  ; 
 DCF <=  DCF & qrq  |  DBF & QRQ  ; 
 OAF <=  RAF & TBA  |  KAF & TCA  ; 
 KAN <=  KAN & tkb & tjb  |  CBF & TKB  |  NAN & TJB  ; 
 PEB <=  PEB & tlf & tle  |  PEA & TLF  ; 
 PFB <=  PEB & tlf & tle  |  PEA & TLF  ; 
 OAN <=  RBF & TBB  |  KAN & TCB  ; 
 KBF <=  KBF & tkc & tjc  |  CBF & TKC  |  NBF & TJC  ; 
 CAF <=  CAF & tfa & tfb  |  DCF & TFA  |  EBF & TFB  ; 
 CBF <=  CAF & tfa & tfb  |  DCF & TFA  |  EBF & TFB  ; 
 OBF <=  RCF & TBC  |  KBF & TCC  |  RAF & TDC  ; 
 KBN <=  KBN & tkd & tjf  |  CBF & TKD  |  NBN & TJF  ; 
 OBN <=  RDF & TBD  |  KBN & TCD  |  RBF & TDD  ; 
 QVA <=  GAA & gab & gac  |  gaa & GAB & gac  |  gaa & gab & GAC  |  GAA & GAB & GAC  ;
 OFF <= CAF ; 
 OHF <= CAF ; 
 OJN <= ABK ; 
 OJO <= ABL ; 
 qnb <=  qsn  |  QSJ  |  pea  ; 
 qnh <=  qsn  |  QSJ  |  PEA  ; 
 QSB <=  QSB & qrp  |  DAJ & QRP  ; 
 QSJ <=  QSJ & qrp  |  QSB & QRP  ; 
 qmj <=  qmf  |  RGE  |  RGG  ; 
 qmk <=  qmf  |  RGE  |  rgg  ; 
 QSN <= QSJ ; 
 OFI <=  QBH & qsj & qso  |  QIG  |  QNH  ; 
 QBH <=  QBH & qsj & qso  |  QIG  |  QNH  ; 
 ODG <=  QJH  |  QMF & RDE  ; 
 ODH <=  QJL  |  QMC & RDE  ; 
 OCF <= RBF ; 
 VAG <=  QNG & PBG  ; 
 VBG <=  QNG & PBG  ; 
 HAG <=  RAG & TGA  |  IAG & TGB  ; 
 HAO <=  RAO & TGA  |  IAO & TGB  ; 
 NAG <= IAG ; 
 NAO <= IAO ; 
 NBG <= IBG ; 
 NBO <= IBO ; 
 PAG <=  PAG & taj & teg  |  PAF & TAJ  |  JCG & TEG  ; 
 PAO <=  PAG & taj & teg  |  PAF & TAJ  |  JCG & TEG  ; 
 PBG <=  PAG & taj & teg  |  PAF & TAJ  |  JCG & TEG  ; 
 RAG <=  MAG & TAA  |  MBG & TAB  |  MCG & TAC  |  MDG & TAD  |  LAG  ; 
 RAO <=  MAG & TAA  |  MBG & TAB  |  MCG & TAC  |  MDG & TAD  |  LAG  ; 
 RBG <= RAG ; 
 RCG <= RBG ; 
 RDG <= RCG ; 
 REG <= RDG ; 
 gag <= rag ; 
 gcg <= rag ; 
 RFG <= REG ; 
 RGG <= RFG ; 
 QBE <=  QSO & qnf  |  JFI  ; 
 KAG <=  KAG & tka & tja  |  CBG & TKA  |  NAG & TJA  ; 
 DBG <=  DBG & qrq  |  DAG & QRQ  ; 
 DCG <=  DCG & qrq  |  DBG & QRQ  ; 
 OAG <=  RAG & TBA  |  KAG & TCA  ; 
 KAO <=  KAO & tkb & tjb  |  CBG & TKB  |  NAO & TJB  ; 
 PEC <=  PEC & tlf & tle  |  PEB & TLF  ; 
 PFC <=  PEC & tlf & tle  |  PEB & TLF  ; 
 OAO <=  RBG & TBB  |  KAO & TCB  ; 
 KBG <=  KBG & tkc & tjc  |  CBG & TKC  |  NBG & TJC  ; 
 CAG <=  CAG & tfa & tfb  |  DCG & TFA  |  EBG & TFB  ; 
 CBG <=  CAG & tfa & tfb  |  DCG & TFA  |  EBG & TFB  ; 
 OBG <=  RCG & TBC  |  KBG & TCC  |  RAG & TDC  ; 
 KBO <=  KBO & tkd & tjf  |  CBG & TKD  |  NBO & TJF  ; 
 OBO <=  RDG & TBD  |  KBO & TCD  |  RBG & TDD  ; 
 QVB <=  GAD & gae & gaf  |  gad & GAE & gaf  |  gad & gae & GAF  |  GAD & GAE & GAF  ;
 OFG <= CAG ; 
 OHG <= CAG ; 
 QSQ <= IGB ; 
 qnc <=  QSO  |  qsk  ; 
 QSC <=  QSC & qrp  |  DAK & QRP  ; 
 QSK <=  QSK & qrp  |  JQC & QRP  ; 
 QBF <= QNR ; 
 QBL <= QBD ; 
 QNR <= QNC ; 
 QSP <= QSO ; 
 ODK <= QBD ; 
 OGE <= QBL ; 
 QBD <= QSO ; 
 QSO <= QSK ; 
 OGA <= QSK ; 
 OGB <= QSK ; 
 OGC <= QSK ; 
 OGD <= QSK ; 
 OCG <= RBG ; 
 VAH <=  QNG & PBH  ; 
 VBH <=  QNG & PBH  ; 
 QRA <= jff ; 
 QRB <= QRA ; 
 QRC <= QRB ; 
 QRD <= QRC ; 
 QRE <= jfg ; 
 QRF <= QRE ; 
 QRG <= QRF ; 
 QRH <= QRG ; 
 QRI <= QRH ; 
 QRJ <= jfh ; 
 QRK <= QRJ ; 
 QRL <= QRK ; 
 QRM <= QRL ; 
 QRN <= QRM ; 
 QRO <= QRN ; 
 HAH <=  RAH & TGA  |  IAH & TGB  ; 
 NAH <= IAH ; 
 NAP <= IAP ; 
 NBH <= IBH ; 
 NBP <= IBP ; 
 qrr <= iga ; 
 PAH <=  PAH & taj & teg  |  PAG & TAJ  |  JCH & TEG  ; 
 PAP <=  PAH & taj & teg  |  PAG & TAJ  |  JCH & TEG  ; 
 PBH <=  PAH & taj & teg  |  PAG & TAJ  |  JCH & TEG  ; 
 RAH <=  MAH & TAA  |  MBH & TAB  |  MCH & TAC  |  MDH & TAD  |  LAH  ; 
 RAP <=  MAH & TAA  |  MBH & TAB  |  MCH & TAC  |  MDH & TAD  |  LAH  ; 
 RBH <= RAH ; 
 RCH <= RBH ; 
 RDH <= RCH ; 
 gah <= rah ; 
 gai <= raq ; 
 QNM <= QNL ; 
 QNN <= QNM ; 
 QNO <= QNN ; 
 QNP <= QNO ; 
 QNI <= QND ; 
 QNJ <= QNI ; 
 QNK <= QNJ ; 
 QNL <= QNK ; 
 KAH <=  KAH & tka & tja  |  CBH & TKA  |  NAH & TJA  ; 
 QRP <=  QRA & QRE & QRJ  |  QRR  ; 
 QRQ <=  QRA & QRE & QRJ  |  QRR  ; 
 DBH <=  DBH & qrq  |  DAH & QRQ  ; 
 DCH <=  DCH & qrq  |  DBH & QRQ  ; 
 OAH <=  RAH & TBA  |  KAH & TCA  ; 
 KAP <=  KAP & tkb & tjb  |  CBH & TKB  |  NAP & TJB  ; 
 PED <=  PED & tlf & tle  |  PEC & TLF  ; 
 PFD <=  PED & tlf & tle  |  PEC & TLF  ; 
 OAP <=  RBH & TBB  |  KAP & TCB  ; 
 KBH <=  KBH & tkc & tjc  |  CBH & TKC  |  NBH & TJC  ; 
 CAH <=  CAH & tfa & tfb  |  DCH & TFA  |  EBH & TFB  ; 
 CBH <=  CAH & tfa & tfb  |  DCH & TFA  |  EBH & TFB  ; 
 OBH <=  RCH & TBC  |  KBH & TCC  |  RAH & TDC  ; 
 KBP <=  KBP & tkd & tjf  |  CBH & TKD  |  NBP & TJF  ; 
 OBP <=  RDH & TBD  |  KBP & TCD  |  RBH & TDD  ; 
 QVC <=  GAG & gah & gai  |  gag & GAH & gai  |  gag & gah & GAI  |  GAG & GAH & GAI  ;
 OFL <=  QDC & qnp & qsl  |  ICE  ; 
 QDC <=  QDC & qnp & qsl  |  ICE  ; 
 OFH <= CAH ; 
 OHH <= CAH ; 
 qnd <=  qso  |  QSK  ; 
 QNG <=  QNE  |  QNF  ; 
 QSD <=  QSD & qrp  |  DAL & QRP  ; 
 QSL <=  QSL & qrp  |  QSD & QRP  ; 
 QNF <= QNE ; 
 OCH <= RBH ; 
 ohi <=  qna  |  qsk  |  qsl  ; 
 qne <=  qna  |  qsk  |  QSL  ; 
 OFK <=  QDB & qnp & qsl  |  JNI & QQF  ; 
 QDB <=  QDB & qnp & qsl  |  JNI & QQF  ; 
end
ram_4096x1 sinst_000(MAA,JMA,{faa,fab,fac,fad,fae,faf,fag,fah,fai,faj,fak,fal}, UAA, VAA, IZZ); 
ram_4096x1 sinst_001(MAB,JMB,{faa,fab,fac,fad,fae,faf,fag,fah,fai,faj,fak,fal}, UAA, VAA, IZZ); 
ram_4096x1 sinst_002(MAC,JMC,{faa,fab,fac,fad,fae,faf,fag,fah,fai,faj,fak,fal}, UAA, VAA, IZZ); 
ram_4096x1 sinst_003(MAD,JMD,{faa,fab,fac,fad,fae,faf,fag,fah,fai,faj,fak,fal}, UAA, VAA, IZZ); 
ram_4096x1 sinst_004(MAE,JME,{FAA,FAB,FAC,FAD,FAE,FAF,FAG,FAG,FAI,FAJ,FAK,FAL}, UAA, VBA, IZZ); 
ram_4096x1 sinst_005(MAF,JMF,{FAA,FAB,FAC,FAD,FAE,FAF,FAG,FAG,FAI,FAJ,FAK,FAL}, UAA, VBA, IZZ); 
ram_4096x1 sinst_006(MAG,JMG,{FAA,FAB,FAC,FAD,FAE,FAF,FAG,FAG,FAI,FAJ,FAK,FAL}, UAA, VBA, IZZ); 
ram_4096x1 sinst_007(MAH,JMH,{FAA,FAB,FAC,FAD,FAE,FAF,FAG,FAG,FAI,FAJ,FAK,FAL}, UAA, VBA, IZZ); 
ram_4096x1 sinst_008(MAI,JMI,{FAA,FAB,FAC,FAD,FAE,FAF,FAG,FAG,FAI,FAJ,FAK,FAL}, UAA, VBA, IZZ); 
ram_4096x1 sinst_009(MBA,JMA,{fba,fbb,fbc,fbd,fbe,fbf,fbg,fbh,fbi,fbj,fbk,fbl}, UAA, VAA, IZZ); 
ram_4096x1 sinst_010(MBB,JMB,{fba,fbb,fbc,fbd,fbe,fbf,fbg,fbh,fbi,fbj,fbk,fbl}, UAA, VAA, IZZ); 
ram_4096x1 sinst_011(MBC,JMC,{fba,fbb,fbc,fbd,fbe,fbf,fbg,fbh,fbi,fbj,fbk,fbl}, UAA, VAA, IZZ); 
ram_4096x1 sinst_012(MBD,JMD,{fba,fbb,fbc,fbd,fbe,fbf,fbg,fbh,fbi,fbj,fbk,fbl}, UAA, VAA, IZZ); 
ram_4096x1 sinst_013(MBE,JME,{FBA,FBB,FBC,FBD,FBE,FBF,FBG,FBG,FBI,FBJ,FBK,FBL}, UAA, VBA, IZZ); 
ram_4096x1 sinst_014(MBF,JMF,{FBA,FBB,FBC,FBD,FBE,FBF,FBG,FBG,FBI,FBJ,FBK,FBL}, UAA, VBA, IZZ); 
ram_4096x1 sinst_015(MBG,JMG,{FBA,FBB,FBC,FBD,FBE,FBF,FBG,FBG,FBI,FBJ,FBK,FBL}, UAA, VBA, IZZ); 
ram_4096x1 sinst_016(MBH,JMH,{FBA,FBB,FBC,FBD,FBE,FBF,FBG,FBG,FBI,FBJ,FBK,FBL}, UAA, VBA, IZZ); 
ram_4096x1 sinst_017(MBI,JMI,{FBA,FBB,FBC,FBD,FBE,FBF,FBG,FBG,FBI,FBJ,FBK,FBL}, UAA, VBA, IZZ); 
ram_4096x1 sinst_018(MCA,JMA,{fca,fcb,fcc,fcd,fce,fcf,fcg,fch,fci,fcj,fck,fcl}, UAC, VAC, IZZ); 
ram_4096x1 sinst_019(MCB,JMB,{fca,fcb,fcc,fcd,fce,fcf,fcg,fch,fci,fcj,fck,fcl}, UAC, VAC, IZZ); 
ram_4096x1 sinst_020(MCC,JMC,{fca,fcb,fcc,fcd,fce,fcf,fcg,fch,fci,fcj,fck,fcl}, UAC, VAC, IZZ); 
ram_4096x1 sinst_021(MCD,JMD,{fca,fcb,fcc,fcd,fce,fcf,fcg,fch,fci,fcj,fck,fcl}, UAC, VAC, IZZ); 
ram_4096x1 sinst_022(MCE,JME,{FCA,FCB,FCC,FCD,FCE,FCF,FCG,FCG,FCI,FCJ,FCK,FCL}, UAC, VBC, IZZ); 
ram_4096x1 sinst_023(MCF,JMF,{FCA,FCB,FCC,FCD,FCE,FCF,FCG,FCG,FCI,FCJ,FCK,FCL}, UAC, VBC, IZZ); 
ram_4096x1 sinst_024(MCG,JMG,{FCA,FCB,FCC,FCD,FCE,FCF,FCG,FCG,FCI,FCJ,FCK,FCL}, UAC, VBC, IZZ); 
ram_4096x1 sinst_025(MCH,JMH,{FCA,FCB,FCC,FCD,FCE,FCF,FCG,FCG,FCI,FCJ,FCK,FCL}, UAC, VBC, IZZ); 
ram_4096x1 sinst_026(MCI,JMI,{FCA,FCB,FCC,FCD,FCE,FCF,FCG,FCG,FCI,FCJ,FCK,FCL}, UAC, VBC, IZZ); 
ram_4096x1 sinst_027(MDA,JMA,{fda,fdb,fdc,fdd,fde,fdf,fdg,fdh,fdi,fdj,fdk,fdl}, UAD, VAD, IZZ); 
ram_4096x1 sinst_028(MDB,JMB,{fda,fdb,fdc,fdd,fde,fdf,fdg,fdh,fdi,fdj,fdk,fdl}, UAD, VAD, IZZ); 
ram_4096x1 sinst_029(MDC,JMC,{fda,fdb,fdc,fdd,fde,fdf,fdg,fdh,fdi,fdj,fdk,fdl}, UAD, VAD, IZZ); 
ram_4096x1 sinst_030(MDD,JMD,{fda,fdb,fdc,fdd,fde,fdf,fdg,fdh,fdi,fdj,fdk,fdl}, UAD, VAD, IZZ); 
ram_4096x1 sinst_031(MDE,JME,{FDA,FDB,FDC,FDD,FDE,FDF,FDG,FDG,FDI,FDJ,FDK,FDL}, UAD, VBD, IZZ); 
ram_4096x1 sinst_032(MDF,JMF,{FDA,FDB,FDC,FDD,FDE,FDF,FDG,FDG,FDI,FDJ,FDK,FDL}, UAD, VBD, IZZ); 
ram_4096x1 sinst_033(MDG,JMG,{FDA,FDB,FDC,FDD,FDE,FDF,FDG,FDG,FDI,FDJ,FDK,FDL}, UAD, VBD, IZZ); 
ram_4096x1 sinst_034(MDH,JMH,{FDA,FDB,FDC,FDD,FDE,FDF,FDG,FDG,FDI,FDJ,FDK,FDL}, UAD, VBD, IZZ); 
ram_4096x1 sinst_035(MDI,JMI,{FDA,FDB,FDC,FDD,FDE,FDF,FDG,FDG,FDI,FDJ,FDK,FDL}, UAD, VBD, IZZ); 
ram_4096x1 sinst_036(MAA,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_037(MAB,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_038(MAC,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_039(MAD,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_040(MAE,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_041(MAF,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_042(MAG,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_043(MAH,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_044(MAI,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_045(MBA,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_046(MBB,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_047(MBC,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_048(MBD,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_049(MBF,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_050(MBG,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_051(MBH,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_052(MBI,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_053(MCA,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_054(MCB,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_055(MCC,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_056(MCD,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_057(MCE,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_058(MCF,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_059(MCG,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_060(MCH,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_061(MCI,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_062(MDA,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_063(MDB,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_064(MDC,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_065(MDD,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_066(MDE,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_067(MDF,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_068(MDG,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_069(MDH,,{,,,,,,,,,,,}, , , IZZ); 
ram_4096x1 sinst_070(MDI,,{,,,,,,,,,,,}, , , IZZ); 
endmodule;
