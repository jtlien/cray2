module jc( IZZ,
 IAA, 
 IAB, 
 IBA, 
 IBB, 
 IBC, 
 IBD, 
 IBE, 
 ICA, 
 ICB, 
 IDA, 
 IDB, 
 IDC, 
 IDD, 
 IEA, 
 IEB, 
 IEC, 
 IED, 
 IEE, 
 IFA, 
 IFB, 
 IFC, 
 IFD, 
 IFE, 
 IFFF , 
 IGA, 
 IHA, 
 IHB, 
 OAA, 
 OAB, 
 OAC, 
 OAD, 
 OAE, 
 OAF, 
 OAG, 
 OAH, 
 OAI, 
 OAJ, 
 OAK, 
 OAL, 
 OAM, 
 OAN, 
 OAO, 
 OAP, 
 OBA, 
 OBB, 
 OBC, 
 OBD, 
 OBE, 
 OBF, 
 OBG, 
 OBH, 
 OBI, 
 OBJ, 
 OBK, 
 OBL, 
 OBM, 
 OBN, 
 OBO, 
 OBP, 
 OCA, 
 OCB, 
 OCC, 
 OCD, 
 OCE, 
 OCF, 
 OCG, 
 OCH, 
 OCI, 
 OCJ, 
 OCK, 
 OCL, 
 OCM, 
 OCN, 
 OCO, 
 OCP, 
 ODA, 
 ODB, 
 ODC, 
 ODD, 
 ODE, 
 ODF, 
 ODG, 
 ODH, 
 ODI, 
 ODJ, 
 ODK, 
 ODL, 
 ODM, 
 ODN, 
 ODO, 
 ODP, 
 OEA, 
 OEB, 
 OEC, 
 OED, 
 OEE, 
 OEF, 
 OEG, 
 OEH, 
 OEI, 
 OEJ, 
 OEK, 
 OEL, 
 OEM, 
 OEN, 
 OEO, 
 OEP, 
 OFA, 
 OFB, 
 OFC, 
 OFD, 
 OFE, 
 OFF, 
 OFG, 
 OFH, 
 OFI, 
 OFJ, 
 OFK, 
 OFL, 
 OFM, 
 OFN, 
 OFO, 
 OFP, 
 OGA, 
 OGB, 
 OGC, 
 OGD, 
 OGE, 
 OGF, 
 OGG, 
 OGH, 
 OGI, 
 OGJ, 
 OGK, 
 OGL, 
 OGM, 
 OGN, 
 OGO, 
 OGP, 
 OHA, 
 OHB, 
 OHC, 
 OHD, 
 OHE, 
 OHF, 
 OHG, 
 OHH, 
 OHI, 
 OHJ, 
 OHK, 
 OHL, 
 OHM, 
 OHN, 
 OHO, 
 OHP, 
 OIA, 
 OIB, 
 OIC, 
 OID, 
 OIE, 
 OIF, 
 OIG, 
 OIH, 
 OII, 
 OIJ, 
 OIK, 
 OIL, 
 OIM, 
 OIN, 
 OIO, 
 OIP, 
 OJA, 
 OJB, 
 OJC, 
 OJD, 
 OJE, 
 OJF, 
 OJG, 
 OJH, 
 OJI, 
 OJJ, 
 OJK, 
 OJL, 
 OJM, 
 OJN, 
 OJO, 
 OJP, 
 OKA, 
 OKB, 
 OKC, 
 OKD, 
 OKE, 
 OKF, 
 OKG, 
 OKH, 
 OKI, 
 OKJ, 
 OKK, 
 OKL, 
 OKM, 
 OKN, 
 OKO, 
 OKP, 
 OLA, 
 OLB, 
 OLC, 
 OLD, 
 OLE, 
 OLF, 
 OLG, 
 OLH, 
 OLI, 
 OLJ, 
 OLK, 
 OLL, 
 OLM, 
 OLN, 
 OLO, 
 OLP, 
 OMA, 
 OMB, 
 OMC, 
 OMD, 
 OME, 
 OMF, 
 OMG, 
 OMH, 
 OMI, 
 OMJ, 
 OMK, 
 OML, 
 OMM, 
 OMN, 
 OMO, 
 OMP, 
 ONA, 
 ONB, 
 ONC, 
 OND, 
 ONE, 
 ONF, 
 ONG, 
 ONH, 
 ONI, 
 ONJ, 
 ONK, 
 ONL, 
 ONM, 
 ONN, 
 ONO, 
 ONP, 
 OOA, 
 OOB, 
 OOC, 
 OOD, 
 OOE, 
 OOF, 
 OOG, 
 OOH, 
 OOI, 
 OOJ, 
 OOK, 
 OOL, 
 OOM, 
 OON, 
 OOO, 
 OOP, 
 OPA, 
 OPB, 
 OPC, 
 OPD, 
 OPE, 
 OPF, 
 OPG, 
 OPH, 
 OPI, 
 OPJ, 
 OPK, 
 OPL, 
 OPM, 
 OPN, 
 OPO, 
 OPP, 
 OQA, 
 OQB, 
 OQC, 
OQD ); 
    
 input IZZ; 
 input IAA; 
 input IAB; 
 input IBA; 
 input IBB; 
 input IBC; 
 input IBD; 
 input IBE; 
 input ICA; 
 input ICB; 
 input IDA; 
 input IDB; 
 input IDC; 
 input IDD; 
 input IEA; 
 input IEB; 
 input IEC; 
 input IED; 
 input IEE; 
 input IFA; 
 input IFB; 
 input IFC; 
 input IFD; 
 input IFE; 
 input IFFF ; 
 input IGA; 
 input IHA; 
 input IHB; 

 output OAA; 
 output OAB; 
 output OAC; 
 output OAD; 
 output OAE; 
 output OAF; 
 output OAG; 
 output OAH; 
 output OAI; 
 output OAJ; 
 output OAK; 
 output OAL; 
 output OAM; 
 output OAN; 
 output OAO; 
 output OAP; 
 output OBA; 
 output OBB; 
 output OBC; 
 output OBD; 
 output OBE; 
 output OBF; 
 output OBG; 
 output OBH; 
 output OBI; 
 output OBJ; 
 output OBK; 
 output OBL; 
 output OBM; 
 output OBN; 
 output OBO; 
 output OBP; 
 output OCA; 
 output OCB; 
 output OCC; 
 output OCD; 
 output OCE; 
 output OCF; 
 output OCG; 
 output OCH; 
 output OCI; 
 output OCJ; 
 output OCK; 
 output OCL; 
 output OCM; 
 output OCN; 
 output OCO; 
 output OCP; 
 output ODA; 
 output ODB; 
 output ODC; 
 output ODD; 
 output ODE; 
 output ODF; 
 output ODG; 
 output ODH; 
 output ODI; 
 output ODJ; 
 output ODK; 
 output ODL; 
 output ODM; 
 output ODN; 
 output ODO; 
 output ODP; 
 output OEA; 
 output OEB; 
 output OEC; 
 output OED; 
 output OEE; 
 output OEF; 
 output OEG; 
 output OEH; 
 output OEI; 
 output OEJ; 
 output OEK; 
 output OEL; 
 output OEM; 
 output OEN; 
 output OEO; 
 output OEP; 
 output OFA; 
 output OFB; 
 output OFC; 
 output OFD; 
 output OFE; 
 output OFF; 
 output OFG; 
 output OFH; 
 output OFI; 
 output OFJ; 
 output OFK; 
 output OFL; 
 output OFM; 
 output OFN; 
 output OFO; 
 output OFP; 
 output OGA; 
 output OGB; 
 output OGC; 
 output OGD; 
 output OGE; 
 output OGF; 
 output OGG; 
 output OGH; 
 output OGI; 
 output OGJ; 
 output OGK; 
 output OGL; 
 output OGM; 
 output OGN; 
 output OGO; 
 output OGP; 
 output OHA; 
 output OHB; 
 output OHC; 
 output OHD; 
 output OHE; 
 output OHF; 
 output OHG; 
 output OHH; 
 output OHI; 
 output OHJ; 
 output OHK; 
 output OHL; 
 output OHM; 
 output OHN; 
 output OHO; 
 output OHP; 
 output OIA; 
 output OIB; 
 output OIC; 
 output OID; 
 output OIE; 
 output OIF; 
 output OIG; 
 output OIH; 
 output OII; 
 output OIJ; 
 output OIK; 
 output OIL; 
 output OIM; 
 output OIN; 
 output OIO; 
 output OIP; 
 output OJA; 
 output OJB; 
 output OJC; 
 output OJD; 
 output OJE; 
 output OJF; 
 output OJG; 
 output OJH; 
 output OJI; 
 output OJJ; 
 output OJK; 
 output OJL; 
 output OJM; 
 output OJN; 
 output OJO; 
 output OJP; 
 output OKA; 
 output OKB; 
 output OKC; 
 output OKD; 
 output OKE; 
 output OKF; 
 output OKG; 
 output OKH; 
 output OKI; 
 output OKJ; 
 output OKK; 
 output OKL; 
 output OKM; 
 output OKN; 
 output OKO; 
 output OKP; 
 output OLA; 
 output OLB; 
 output OLC; 
 output OLD; 
 output OLE; 
 output OLF; 
 output OLG; 
 output OLH; 
 output OLI; 
 output OLJ; 
 output OLK; 
 output OLL; 
 output OLM; 
 output OLN; 
 output OLO; 
 output OLP; 
 output OMA; 
 output OMB; 
 output OMC; 
 output OMD; 
 output OME; 
 output OMF; 
 output OMG; 
 output OMH; 
 output OMI; 
 output OMJ; 
 output OMK; 
 output OML; 
 output OMM; 
 output OMN; 
 output OMO; 
 output OMP; 
 output ONA; 
 output ONB; 
 output ONC; 
 output OND; 
 output ONE; 
 output ONF; 
 output ONG; 
 output ONH; 
 output ONI; 
 output ONJ; 
 output ONK; 
 output ONL; 
 output ONM; 
 output ONN; 
 output ONO; 
 output ONP; 
 output OOA; 
 output OOB; 
 output OOC; 
 output OOD; 
 output OOE; 
 output OOF; 
 output OOG; 
 output OOH; 
 output OOI; 
 output OOJ; 
 output OOK; 
 output OOL; 
 output OOM; 
 output OON; 
 output OOO; 
 output OOP; 
 output OPA; 
 output OPB; 
 output OPC; 
 output OPD; 
 output OPE; 
 output OPF; 
 output OPG; 
 output OPH; 
 output OPI; 
 output OPJ; 
 output OPK; 
 output OPL; 
 output OPM; 
 output OPN; 
 output OPO; 
 output OPP; 
 output OQA; 
 output OQB; 
 output OQC; 
 output OQD; 
  
  
reg  aaa ;
reg  aab ;
reg  aac ;
reg  aad ;
reg  aba ;
reg  abb ;
reg  abc ;
reg  abd ;
reg  haa ;
reg  hab ;
reg  hac ;
reg  had ;
reg  hae ;
reg  haf ;
reg  hag ;
reg  hah ;
reg  hai ;
reg  haj ;
reg  hak ;
reg  hal ;
reg  ham ;
reg  han ;
reg  hao ;
reg  hap ;
reg  hba ;
reg  hbb ;
reg  hbc ;
reg  hbd ;
reg  hbe ;
reg  hbf ;
reg  hbg ;
reg  hbh ;
reg  hbi ;
reg  hbj ;
reg  hbk ;
reg  hbl ;
reg  hbm ;
reg  hbn ;
reg  hbo ;
reg  hbp ;
reg  hca ;
reg  hcb ;
reg  hcc ;
reg  hcd ;
reg  hce ;
reg  hcf ;
reg  hcg ;
reg  hch ;
reg  hci ;
reg  hcj ;
reg  hck ;
reg  hcl ;
reg  hcm ;
reg  hcn ;
reg  hco ;
reg  hcp ;
reg  hda ;
reg  hdb ;
reg  hdc ;
reg  hdd ;
reg  hde ;
reg  hdf ;
reg  hdg ;
reg  hdh ;
reg  hdi ;
reg  hdj ;
reg  hdk ;
reg  hdl ;
reg  hdm ;
reg  hdn ;
reg  hdo ;
reg  hdp ;
reg  hea ;
reg  heb ;
reg  hec ;
reg  hed ;
reg  hee ;
reg  hef ;
reg  heg ;
reg  heh ;
reg  hei ;
reg  hej ;
reg  hek ;
reg  hel ;
reg  hem ;
reg  hen ;
reg  heo ;
reg  hep ;
reg  hfa ;
reg  hfb ;
reg  hfc ;
reg  hfd ;
reg  hfe ;
reg  hff ;
reg  hfg ;
reg  hfh ;
reg  hfi ;
reg  hfj ;
reg  hfk ;
reg  hfl ;
reg  hfm ;
reg  hfn ;
reg  hfo ;
reg  hfp ;
reg  hga ;
reg  hgb ;
reg  hgc ;
reg  hgd ;
reg  hge ;
reg  hgf ;
reg  hgg ;
reg  hgh ;
reg  hgi ;
reg  hgj ;
reg  hgk ;
reg  hgl ;
reg  hgm ;
reg  hgn ;
reg  hgo ;
reg  hgp ;
reg  hha ;
reg  hhb ;
reg  hhc ;
reg  hhd ;
reg  hhe ;
reg  hhf ;
reg  hhg ;
reg  hhh ;
reg  hhi ;
reg  hhj ;
reg  hhk ;
reg  hhl ;
reg  hhm ;
reg  hhn ;
reg  hho ;
reg  hhp ;
reg  KAC ;
reg  KAD ;
reg  KAE ;
reg  KAF ;
reg  KCC ;
reg  KCD ;
reg  KCE ;
reg  KCF ;
reg  KEC ;
reg  KED ;
reg  KEE ;
reg  KEF ;
reg  KGC ;
reg  KGD ;
reg  KGE ;
reg  KGF ;
reg  LAA ;
reg  LAB ;
reg  LAC ;
reg  LAD ;
reg  LAE ;
reg  LAF ;
reg  LBA ;
reg  LBB ;
reg  LBC ;
reg  LBD ;
reg  LBE ;
reg  LCA ;
reg  LCB ;
reg  LCC ;
reg  LCD ;
reg  LCE ;
reg  LCF ;
reg  LDA ;
reg  LDB ;
reg  LDC ;
reg  LDD ;
reg  LDE ;
reg  LEA ;
reg  LEB ;
reg  LEC ;
reg  LED ;
reg  LEE ;
reg  LEF ;
reg  LFA ;
reg  LFB ;
reg  LFC ;
reg  LFD ;
reg  LFE ;
reg  LGA ;
reg  LGB ;
reg  LGC ;
reg  LGD ;
reg  LGE ;
reg  LGF ;
reg  LHA ;
reg  LHB ;
reg  LHC ;
reg  LHD ;
reg  LHE ;
reg  OAA ;
reg  OAB ;
reg  OAC ;
reg  OAD ;
reg  OAE ;
reg  OAF ;
reg  OAG ;
reg  OAH ;
reg  OAI ;
reg  OAJ ;
reg  OAK ;
reg  OAL ;
reg  OAM ;
reg  OAN ;
reg  OAO ;
reg  OAP ;
reg  OBA ;
reg  OBB ;
reg  OBC ;
reg  OBD ;
reg  OBE ;
reg  OBF ;
reg  OBG ;
reg  OBH ;
reg  OBI ;
reg  OBJ ;
reg  OBK ;
reg  OBL ;
reg  OBM ;
reg  OBN ;
reg  OBO ;
reg  OBP ;
reg  OCA ;
reg  OCB ;
reg  OCC ;
reg  OCD ;
reg  OCE ;
reg  OCF ;
reg  OCG ;
reg  OCH ;
reg  OCI ;
reg  OCJ ;
reg  OCK ;
reg  OCL ;
reg  OCM ;
reg  OCN ;
reg  OCO ;
reg  OCP ;
reg  ODA ;
reg  ODB ;
reg  ODC ;
reg  ODD ;
reg  ODE ;
reg  ODF ;
reg  ODG ;
reg  ODH ;
reg  ODI ;
reg  ODJ ;
reg  ODK ;
reg  ODL ;
reg  ODM ;
reg  ODN ;
reg  ODO ;
reg  ODP ;
reg  OEA ;
reg  OEB ;
reg  OEC ;
reg  OED ;
reg  OEE ;
reg  OEF ;
reg  OEG ;
reg  OEH ;
reg  OEI ;
reg  OEJ ;
reg  OEK ;
reg  OEL ;
reg  OEM ;
reg  OEN ;
reg  OEO ;
reg  OEP ;
reg  OFA ;
reg  OFB ;
reg  OFC ;
reg  OFD ;
reg  OFE ;
reg  OFF ;
reg  OFG ;
reg  OFH ;
reg  OFI ;
reg  OFJ ;
reg  OFK ;
reg  OFL ;
reg  OFM ;
reg  OFN ;
reg  OFO ;
reg  OFP ;
reg  OGA ;
reg  OGB ;
reg  OGC ;
reg  OGD ;
reg  OGE ;
reg  OGF ;
reg  OGG ;
reg  OGH ;
reg  OGI ;
reg  OGJ ;
reg  OGK ;
reg  OGL ;
reg  OGM ;
reg  OGN ;
reg  OGO ;
reg  OGP ;
reg  OHA ;
reg  OHB ;
reg  OHC ;
reg  OHD ;
reg  OHE ;
reg  OHF ;
reg  OHG ;
reg  OHH ;
reg  OHI ;
reg  OHJ ;
reg  OHK ;
reg  OHL ;
reg  OHM ;
reg  OHN ;
reg  OHO ;
reg  OHP ;
reg  OIA ;
reg  OIB ;
reg  OIC ;
reg  OID ;
reg  OIE ;
reg  OIF ;
reg  OIG ;
reg  OIH ;
reg  OII ;
reg  OIJ ;
reg  OIK ;
reg  OIL ;
reg  OIM ;
reg  OIN ;
reg  OIO ;
reg  OIP ;
reg  OJA ;
reg  OJB ;
reg  OJC ;
reg  OJD ;
reg  OJE ;
reg  OJF ;
reg  OJG ;
reg  OJH ;
reg  OJI ;
reg  OJJ ;
reg  OJK ;
reg  OJL ;
reg  OJM ;
reg  OJN ;
reg  OJO ;
reg  OJP ;
reg  OKA ;
reg  OKB ;
reg  OKC ;
reg  OKD ;
reg  OKE ;
reg  OKF ;
reg  OKG ;
reg  OKH ;
reg  OKI ;
reg  OKJ ;
reg  OKK ;
reg  OKL ;
reg  OKM ;
reg  OKN ;
reg  OKO ;
reg  OKP ;
reg  OLA ;
reg  OLB ;
reg  OLC ;
reg  OLD ;
reg  OLE ;
reg  OLF ;
reg  OLG ;
reg  OLH ;
reg  OLI ;
reg  OLJ ;
reg  OLK ;
reg  OLL ;
reg  OLM ;
reg  OLN ;
reg  OLO ;
reg  OLP ;
reg  OMA ;
reg  OMB ;
reg  OMC ;
reg  OMD ;
reg  OME ;
reg  OMF ;
reg  OMG ;
reg  OMH ;
reg  OMI ;
reg  OMJ ;
reg  OMK ;
reg  OML ;
reg  OMM ;
reg  OMN ;
reg  OMO ;
reg  OMP ;
reg  ONA ;
reg  ONB ;
reg  ONC ;
reg  OND ;
reg  ONE ;
reg  ONF ;
reg  ONG ;
reg  ONH ;
reg  ONI ;
reg  ONJ ;
reg  ONK ;
reg  ONL ;
reg  ONM ;
reg  ONN ;
reg  ONO ;
reg  ONP ;
reg  OOA ;
reg  OOB ;
reg  OOC ;
reg  OOD ;
reg  OOE ;
reg  OOF ;
reg  OOG ;
reg  OOH ;
reg  OOI ;
reg  OOJ ;
reg  OOK ;
reg  OOL ;
reg  OOM ;
reg  OON ;
reg  OOO ;
reg  OOP ;
reg  OPA ;
reg  OPB ;
reg  OPC ;
reg  OPD ;
reg  OPE ;
reg  OPF ;
reg  OPG ;
reg  OPH ;
reg  OPI ;
reg  OPJ ;
reg  OPK ;
reg  OPL ;
reg  OPM ;
reg  OPN ;
reg  OPO ;
reg  OPP ;
reg  OQA ;
reg  OQB ;
reg  OQC ;
reg  OQD ;
reg  PAA ;
reg  PAB ;
reg  PAC ;
reg  PAD ;
reg  PBA ;
reg  PBB ;
reg  PBC ;
reg  PBD ;
reg  PCA ;
reg  PCB ;
reg  PCC ;
reg  PCD ;
reg  PDA ;
reg  PDB ;
reg  PDC ;
reg  PDD ;
reg  PEA ;
reg  PEB ;
reg  PEC ;
reg  PED ;
reg  PFA ;
reg  PFB ;
reg  PFC ;
reg  PFD ;
reg  PGA ;
reg  PGB ;
reg  PGC ;
reg  PGD ;
reg  PHA ;
reg  PHB ;
reg  PHC ;
reg  PHD ;
reg  qaa ;
reg  QAB ;
reg  QAC ;
reg  QAD ;
reg  qae ;
reg  qaf ;
reg  qag ;
reg  qah ;
reg  QAI ;
reg  QAJ ;
reg  QAK ;
reg  QAL ;
reg  QAM ;
reg  qan ;
reg  QAP ;
reg  qba ;
reg  QBB ;
reg  qca ;
reg  QCB ;
reg  QCC ;
reg  QCD ;
reg  qce ;
reg  qcf ;
reg  qcg ;
reg  qch ;
reg  QCI ;
reg  QCJ ;
reg  QCK ;
reg  QCL ;
reg  QCM ;
reg  qcn ;
reg  QCP ;
reg  qda ;
reg  QDB ;
reg  qea ;
reg  QEB ;
reg  QEC ;
reg  QED ;
reg  qee ;
reg  qef ;
reg  qeg ;
reg  qeh ;
reg  QEI ;
reg  QEJ ;
reg  QEK ;
reg  QEL ;
reg  QEM ;
reg  qen ;
reg  QEP ;
reg  qfa ;
reg  QFB ;
reg  qga ;
reg  QGB ;
reg  QGC ;
reg  QGD ;
reg  qge ;
reg  qgf ;
reg  qgg ;
reg  qgh ;
reg  QGI ;
reg  QGJ ;
reg  QGK ;
reg  QGL ;
reg  QGM ;
reg  qgn ;
reg  QGP ;
reg  qha ;
reg  QHB ;
reg  QIA ;
reg  qja ;
reg  QKA ;
reg  qkb ;
reg  qla ;
reg  qlb ;
reg  QNA ;
reg  QNB ;
wire  AAA ;
wire  AAB ;
wire  AAC ;
wire  AAD ;
wire  ABA ;
wire  ABB ;
wire  ABC ;
wire  ABD ;
wire  eaa ;
wire  EAA ;
wire  eab ;
wire  EAB ;
wire  eac ;
wire  EAC ;
wire  ead ;
wire  EAD ;
wire  eae ;
wire  EAE ;
wire  eaf ;
wire  EAF ;
wire  eag ;
wire  EAG ;
wire  eah ;
wire  EAH ;
wire  eai ;
wire  EAI ;
wire  eaj ;
wire  EAJ ;
wire  eak ;
wire  EAK ;
wire  eal ;
wire  EAL ;
wire  eam ;
wire  EAM ;
wire  ean ;
wire  EAN ;
wire  eao ;
wire  EAO ;
wire  eap ;
wire  EAP ;
wire  eaq ;
wire  EAQ ;
wire  ear ;
wire  EAR ;
wire  eca ;
wire  ECA ;
wire  ecb ;
wire  ECB ;
wire  ecc ;
wire  ECC ;
wire  ecd ;
wire  ECD ;
wire  ece ;
wire  ECE ;
wire  ecf ;
wire  ECF ;
wire  ecg ;
wire  ECG ;
wire  ech ;
wire  ECH ;
wire  eci ;
wire  ECI ;
wire  ecj ;
wire  ECJ ;
wire  eck ;
wire  ECK ;
wire  ecl ;
wire  ECL ;
wire  ecm ;
wire  ECM ;
wire  ecn ;
wire  ECN ;
wire  eco ;
wire  ECO ;
wire  ecp ;
wire  ECP ;
wire  ecq ;
wire  ECQ ;
wire  ecr ;
wire  ECR ;
wire  eea ;
wire  EEA ;
wire  eeb ;
wire  EEB ;
wire  eec ;
wire  EEC ;
wire  eed ;
wire  EED ;
wire  eee ;
wire  EEE ;
wire  eef ;
wire  EEF ;
wire  eeg ;
wire  EEG ;
wire  eeh ;
wire  EEH ;
wire  eei ;
wire  EEI ;
wire  eej ;
wire  EEJ ;
wire  eek ;
wire  EEK ;
wire  eel ;
wire  EEL ;
wire  eem ;
wire  EEM ;
wire  een ;
wire  EEN ;
wire  eeo ;
wire  EEO ;
wire  eep ;
wire  EEP ;
wire  eeq ;
wire  EEQ ;
wire  eer ;
wire  EER ;
wire  ega ;
wire  EGA ;
wire  egb ;
wire  EGB ;
wire  egc ;
wire  EGC ;
wire  egd ;
wire  EGD ;
wire  ege ;
wire  EGE ;
wire  egf ;
wire  EGF ;
wire  egg ;
wire  EGG ;
wire  egh ;
wire  EGH ;
wire  egi ;
wire  EGI ;
wire  egj ;
wire  EGJ ;
wire  egk ;
wire  EGK ;
wire  egl ;
wire  EGL ;
wire  egm ;
wire  EGM ;
wire  egn ;
wire  EGN ;
wire  ego ;
wire  EGO ;
wire  egp ;
wire  EGP ;
wire  egq ;
wire  EGQ ;
wire  egr ;
wire  EGR ;
wire  gaa ;
wire  GAA ;
wire  gab ;
wire  GAB ;
wire  gac ;
wire  GAC ;
wire  gad ;
wire  GAD ;
wire  gae ;
wire  GAE ;
wire  gaf ;
wire  GAF ;
wire  gag ;
wire  GAG ;
wire  gah ;
wire  GAH ;
wire  gai ;
wire  GAI ;
wire  gaj ;
wire  GAJ ;
wire  gak ;
wire  GAK ;
wire  gal ;
wire  GAL ;
wire  gam ;
wire  GAM ;
wire  gan ;
wire  GAN ;
wire  gao ;
wire  GAO ;
wire  gap ;
wire  GAP ;
wire  gca ;
wire  GCA ;
wire  gcb ;
wire  GCB ;
wire  gcc ;
wire  GCC ;
wire  gcd ;
wire  GCD ;
wire  gce ;
wire  GCE ;
wire  gcf ;
wire  GCF ;
wire  gcg ;
wire  GCG ;
wire  gch ;
wire  GCH ;
wire  gci ;
wire  GCI ;
wire  gcj ;
wire  GCJ ;
wire  gck ;
wire  GCK ;
wire  gcl ;
wire  GCL ;
wire  gcm ;
wire  GCM ;
wire  gcn ;
wire  GCN ;
wire  gco ;
wire  GCO ;
wire  gcp ;
wire  GCP ;
wire  gea ;
wire  GEA ;
wire  geb ;
wire  GEB ;
wire  gec ;
wire  GEC ;
wire  ged ;
wire  GED ;
wire  gee ;
wire  GEE ;
wire  gef ;
wire  GEF ;
wire  geg ;
wire  GEG ;
wire  geh ;
wire  GEH ;
wire  gei ;
wire  GEI ;
wire  gej ;
wire  GEJ ;
wire  gek ;
wire  GEK ;
wire  gel ;
wire  GEL ;
wire  gem ;
wire  GEM ;
wire  gen ;
wire  GEN ;
wire  geo ;
wire  GEO ;
wire  gep ;
wire  GEP ;
wire  gga ;
wire  GGA ;
wire  ggb ;
wire  GGB ;
wire  ggc ;
wire  GGC ;
wire  ggd ;
wire  GGD ;
wire  gge ;
wire  GGE ;
wire  ggf ;
wire  GGF ;
wire  ggg ;
wire  GGG ;
wire  ggh ;
wire  GGH ;
wire  ggi ;
wire  GGI ;
wire  ggj ;
wire  GGJ ;
wire  ggk ;
wire  GGK ;
wire  ggl ;
wire  GGL ;
wire  ggm ;
wire  GGM ;
wire  ggn ;
wire  GGN ;
wire  ggo ;
wire  GGO ;
wire  ggp ;
wire  GGP ;
wire  HAA ;
wire  HAB ;
wire  HAC ;
wire  HAD ;
wire  HAE ;
wire  HAF ;
wire  HAG ;
wire  HAH ;
wire  HAI ;
wire  HAJ ;
wire  HAK ;
wire  HAL ;
wire  HAM ;
wire  HAN ;
wire  HAO ;
wire  HAP ;
wire  HBA ;
wire  HBB ;
wire  HBC ;
wire  HBD ;
wire  HBE ;
wire  HBF ;
wire  HBG ;
wire  HBH ;
wire  HBI ;
wire  HBJ ;
wire  HBK ;
wire  HBL ;
wire  HBM ;
wire  HBN ;
wire  HBO ;
wire  HBP ;
wire  HCA ;
wire  HCB ;
wire  HCC ;
wire  HCD ;
wire  HCE ;
wire  HCF ;
wire  HCG ;
wire  HCH ;
wire  HCI ;
wire  HCJ ;
wire  HCK ;
wire  HCL ;
wire  HCM ;
wire  HCN ;
wire  HCO ;
wire  HCP ;
wire  HDA ;
wire  HDB ;
wire  HDC ;
wire  HDD ;
wire  HDE ;
wire  HDF ;
wire  HDG ;
wire  HDH ;
wire  HDI ;
wire  HDJ ;
wire  HDK ;
wire  HDL ;
wire  HDM ;
wire  HDN ;
wire  HDO ;
wire  HDP ;
wire  HEA ;
wire  HEB ;
wire  HEC ;
wire  HED ;
wire  HEE ;
wire  HEF ;
wire  HEG ;
wire  HEH ;
wire  HEI ;
wire  HEJ ;
wire  HEK ;
wire  HEL ;
wire  HEM ;
wire  HEN ;
wire  HEO ;
wire  HEP ;
wire  HFA ;
wire  HFB ;
wire  HFC ;
wire  HFD ;
wire  HFE ;
wire  HFF ;
wire  HFG ;
wire  HFH ;
wire  HFI ;
wire  HFJ ;
wire  HFK ;
wire  HFL ;
wire  HFM ;
wire  HFN ;
wire  HFO ;
wire  HFP ;
wire  HGA ;
wire  HGB ;
wire  HGC ;
wire  HGD ;
wire  HGE ;
wire  HGF ;
wire  HGG ;
wire  HGH ;
wire  HGI ;
wire  HGJ ;
wire  HGK ;
wire  HGL ;
wire  HGM ;
wire  HGN ;
wire  HGO ;
wire  HGP ;
wire  HHA ;
wire  HHB ;
wire  HHC ;
wire  HHD ;
wire  HHE ;
wire  HHF ;
wire  HHG ;
wire  HHH ;
wire  HHI ;
wire  HHJ ;
wire  HHK ;
wire  HHL ;
wire  HHM ;
wire  HHN ;
wire  HHO ;
wire  HHP ;
wire  iaa ;
wire  iab ;
wire  iba ;
wire  ibb ;
wire  ibc ;
wire  ibd ;
wire  ibe ;
wire  ica ;
wire  icb ;
wire  ida ;
wire  idb ;
wire  idc ;
wire  idd ;
wire  iea ;
wire  ieb ;
wire  iec ;
wire  ied ;
wire  iee ;
wire  ifa ;
wire  ifb ;
wire  ifc ;
wire  ifd ;
wire  ife ;
wire  ifff  ;
wire  iga ;
wire  iha ;
wire  ihb ;
wire  izz ;
wire  jaa ;
wire  JAA ;
wire  jab ;
wire  JAB ;
wire  jac ;
wire  JAC ;
wire  jad ;
wire  JAD ;
wire  jae ;
wire  JAE ;
wire  jaf ;
wire  JAF ;
wire  jag ;
wire  JAG ;
wire  jah ;
wire  JAH ;
wire  jba ;
wire  JBA ;
wire  jbb ;
wire  JBB ;
wire  jbc ;
wire  JBC ;
wire  jbd ;
wire  JBD ;
wire  jbe ;
wire  JBE ;
wire  jbf ;
wire  JBF ;
wire  jbg ;
wire  JBG ;
wire  jbh ;
wire  JBH ;
wire  jca ;
wire  JCA ;
wire  jcb ;
wire  JCB ;
wire  jcc ;
wire  JCC ;
wire  jcd ;
wire  JCD ;
wire  jce ;
wire  JCE ;
wire  jcf ;
wire  JCF ;
wire  jcg ;
wire  JCG ;
wire  jch ;
wire  JCH ;
wire  jda ;
wire  JDA ;
wire  jdb ;
wire  JDB ;
wire  jdc ;
wire  JDC ;
wire  jdd ;
wire  JDD ;
wire  jde ;
wire  JDE ;
wire  jdf ;
wire  JDF ;
wire  jdg ;
wire  JDG ;
wire  jdh ;
wire  JDH ;
wire  jea ;
wire  JEA ;
wire  jeb ;
wire  JEB ;
wire  jec ;
wire  JEC ;
wire  jed ;
wire  JED ;
wire  jee ;
wire  JEE ;
wire  jef ;
wire  JEF ;
wire  jeg ;
wire  JEG ;
wire  jeh ;
wire  JEH ;
wire  jfa ;
wire  JFA ;
wire  jfb ;
wire  JFB ;
wire  jfc ;
wire  JFC ;
wire  jfd ;
wire  JFD ;
wire  jfe ;
wire  JFE ;
wire  jff ;
wire  JFF ;
wire  jfg ;
wire  JFG ;
wire  jfh ;
wire  JFH ;
wire  jga ;
wire  JGA ;
wire  jgb ;
wire  JGB ;
wire  jgc ;
wire  JGC ;
wire  jgd ;
wire  JGD ;
wire  jge ;
wire  JGE ;
wire  jgf ;
wire  JGF ;
wire  jgg ;
wire  JGG ;
wire  jgh ;
wire  JGH ;
wire  jha ;
wire  JHA ;
wire  jhb ;
wire  JHB ;
wire  jhc ;
wire  JHC ;
wire  jhd ;
wire  JHD ;
wire  jhe ;
wire  JHE ;
wire  jhf ;
wire  JHF ;
wire  jhg ;
wire  JHG ;
wire  jhh ;
wire  JHH ;
wire  kac ;
wire  kad ;
wire  kae ;
wire  kaf ;
wire  kcc ;
wire  kcd ;
wire  kce ;
wire  kcf ;
wire  kec ;
wire  ked ;
wire  kee ;
wire  kef ;
wire  kgc ;
wire  kgd ;
wire  kge ;
wire  kgf ;
wire  laa ;
wire  lab ;
wire  lac ;
wire  lad ;
wire  lae ;
wire  laf ;
wire  lba ;
wire  lbb ;
wire  lbc ;
wire  lbd ;
wire  lbe ;
wire  lca ;
wire  lcb ;
wire  lcc ;
wire  lcd ;
wire  lce ;
wire  lcf ;
wire  lda ;
wire  ldb ;
wire  ldc ;
wire  ldd ;
wire  lde ;
wire  lea ;
wire  leb ;
wire  lec ;
wire  led ;
wire  lee ;
wire  lef ;
wire  lfa ;
wire  lfb ;
wire  lfc ;
wire  lfd ;
wire  lfe ;
wire  lga ;
wire  lgb ;
wire  lgc ;
wire  lgd ;
wire  lge ;
wire  lgf ;
wire  lha ;
wire  lhb ;
wire  lhc ;
wire  lhd ;
wire  lhe ;
wire  oaa ;
wire  oab ;
wire  oac ;
wire  oad ;
wire  oae ;
wire  oaf ;
wire  oag ;
wire  oah ;
wire  oai ;
wire  oaj ;
wire  oak ;
wire  oal ;
wire  oam ;
wire  oan ;
wire  oao ;
wire  oap ;
wire  oba ;
wire  obb ;
wire  obc ;
wire  obd ;
wire  obe ;
wire  obf ;
wire  obg ;
wire  obh ;
wire  obi ;
wire  obj ;
wire  obk ;
wire  obl ;
wire  obm ;
wire  obn ;
wire  obo ;
wire  obp ;
wire  oca ;
wire  ocb ;
wire  occ ;
wire  ocd ;
wire  oce ;
wire  ocf ;
wire  ocg ;
wire  och ;
wire  oci ;
wire  ocj ;
wire  ock ;
wire  ocl ;
wire  ocm ;
wire  ocn ;
wire  oco ;
wire  ocp ;
wire  oda ;
wire  odb ;
wire  odc ;
wire  odd ;
wire  ode ;
wire  odf ;
wire  odg ;
wire  odh ;
wire  odi ;
wire  odj ;
wire  odk ;
wire  odl ;
wire  odm ;
wire  odn ;
wire  odo ;
wire  odp ;
wire  oea ;
wire  oeb ;
wire  oec ;
wire  oed ;
wire  oee ;
wire  oef ;
wire  oeg ;
wire  oeh ;
wire  oei ;
wire  oej ;
wire  oek ;
wire  oel ;
wire  oem ;
wire  oen ;
wire  oeo ;
wire  oep ;
wire  ofa ;
wire  ofb ;
wire  ofc ;
wire  ofd ;
wire  ofe ;
wire  off ;
wire  ofg ;
wire  ofh ;
wire  ofi ;
wire  ofj ;
wire  ofk ;
wire  ofl ;
wire  ofm ;
wire  ofn ;
wire  ofo ;
wire  ofp ;
wire  oga ;
wire  ogb ;
wire  ogc ;
wire  ogd ;
wire  oge ;
wire  ogf ;
wire  ogg ;
wire  ogh ;
wire  ogi ;
wire  ogj ;
wire  ogk ;
wire  ogl ;
wire  ogm ;
wire  ogn ;
wire  ogo ;
wire  ogp ;
wire  oha ;
wire  ohb ;
wire  ohc ;
wire  ohd ;
wire  ohe ;
wire  ohf ;
wire  ohg ;
wire  ohh ;
wire  ohi ;
wire  ohj ;
wire  ohk ;
wire  ohl ;
wire  ohm ;
wire  ohn ;
wire  oho ;
wire  ohp ;
wire  oia ;
wire  oib ;
wire  oic ;
wire  oid ;
wire  oie ;
wire  oif ;
wire  oig ;
wire  oih ;
wire  oii ;
wire  oij ;
wire  oik ;
wire  oil ;
wire  oim ;
wire  oin ;
wire  oio ;
wire  oip ;
wire  oja ;
wire  ojb ;
wire  ojc ;
wire  ojd ;
wire  oje ;
wire  ojf ;
wire  ojg ;
wire  ojh ;
wire  oji ;
wire  ojj ;
wire  ojk ;
wire  ojl ;
wire  ojm ;
wire  ojn ;
wire  ojo ;
wire  ojp ;
wire  oka ;
wire  okb ;
wire  okc ;
wire  okd ;
wire  oke ;
wire  okf ;
wire  okg ;
wire  okh ;
wire  oki ;
wire  okj ;
wire  okk ;
wire  okl ;
wire  okm ;
wire  okn ;
wire  oko ;
wire  okp ;
wire  ola ;
wire  olb ;
wire  olc ;
wire  old ;
wire  ole ;
wire  olf ;
wire  olg ;
wire  olh ;
wire  oli ;
wire  olj ;
wire  olk ;
wire  oll ;
wire  olm ;
wire  oln ;
wire  olo ;
wire  olp ;
wire  oma ;
wire  omb ;
wire  omc ;
wire  omd ;
wire  ome ;
wire  omf ;
wire  omg ;
wire  omh ;
wire  omi ;
wire  omj ;
wire  omk ;
wire  oml ;
wire  omm ;
wire  omn ;
wire  omo ;
wire  omp ;
wire  ona ;
wire  onb ;
wire  onc ;
wire  ond ;
wire  one ;
wire  onf ;
wire  ong ;
wire  onh ;
wire  oni ;
wire  onj ;
wire  onk ;
wire  onl ;
wire  onm ;
wire  onn ;
wire  ono ;
wire  onp ;
wire  ooa ;
wire  oob ;
wire  ooc ;
wire  ood ;
wire  ooe ;
wire  oof ;
wire  oog ;
wire  ooh ;
wire  ooi ;
wire  ooj ;
wire  ook ;
wire  ool ;
wire  oom ;
wire  oon ;
wire  ooo ;
wire  oop ;
wire  opa ;
wire  opb ;
wire  opc ;
wire  opd ;
wire  ope ;
wire  opf ;
wire  opg ;
wire  oph ;
wire  opi ;
wire  opj ;
wire  opk ;
wire  opl ;
wire  opm ;
wire  opn ;
wire  opo ;
wire  opp ;
wire  oqa ;
wire  oqb ;
wire  oqc ;
wire  oqd ;
wire  paa ;
wire  pab ;
wire  pac ;
wire  pad ;
wire  pba ;
wire  pbb ;
wire  pbc ;
wire  pbd ;
wire  pca ;
wire  pcb ;
wire  pcc ;
wire  pcd ;
wire  pda ;
wire  pdb ;
wire  pdc ;
wire  pdd ;
wire  pea ;
wire  peb ;
wire  pec ;
wire  ped ;
wire  pfa ;
wire  pfb ;
wire  pfc ;
wire  pfd ;
wire  pga ;
wire  pgb ;
wire  pgc ;
wire  pgd ;
wire  pha ;
wire  phb ;
wire  phc ;
wire  phd ;
wire  QAA ;
wire  qab ;
wire  qac ;
wire  qad ;
wire  QAE ;
wire  QAF ;
wire  QAG ;
wire  QAH ;
wire  qai ;
wire  qaj ;
wire  qak ;
wire  qal ;
wire  qam ;
wire  QAN ;
wire  qap ;
wire  QBA ;
wire  qbb ;
wire  QCA ;
wire  qcb ;
wire  qcc ;
wire  qcd ;
wire  QCE ;
wire  QCF ;
wire  QCG ;
wire  QCH ;
wire  qci ;
wire  qcj ;
wire  qck ;
wire  qcl ;
wire  qcm ;
wire  QCN ;
wire  qcp ;
wire  QDA ;
wire  qdb ;
wire  QEA ;
wire  qeb ;
wire  qec ;
wire  qed ;
wire  QEE ;
wire  QEF ;
wire  QEG ;
wire  QEH ;
wire  qei ;
wire  qej ;
wire  qek ;
wire  qel ;
wire  qem ;
wire  QEN ;
wire  qep ;
wire  QFA ;
wire  qfb ;
wire  QGA ;
wire  qgb ;
wire  qgc ;
wire  qgd ;
wire  QGE ;
wire  QGF ;
wire  QGG ;
wire  QGH ;
wire  qgi ;
wire  qgj ;
wire  qgk ;
wire  qgl ;
wire  qgm ;
wire  QGN ;
wire  qgp ;
wire  QHA ;
wire  qhb ;
wire  qia ;
wire  QJA ;
wire  qka ;
wire  QKB ;
wire  QLA ;
wire  QLB ;
wire  qna ;
wire  qnb ;
wire  taa ;
wire  TAA ;
wire  tab ;
wire  TAB ;
wire  tac ;
wire  TAC ;
wire  tad ;
wire  TAD ;
wire  tae ;
wire  TAE ;
wire  tai ;
wire  TAI ;
wire  taj ;
wire  TAJ ;
wire  tak ;
wire  TAK ;
wire  tam ;
wire  TAM ;
wire  tan ;
wire  TAN ;
wire  tao ;
wire  TAO ;
wire  tap ;
wire  TAP ;
wire  tca ;
wire  TCA ;
wire  tcb ;
wire  TCB ;
wire  tcc ;
wire  TCC ;
wire  tcd ;
wire  TCD ;
wire  tce ;
wire  TCE ;
wire  tci ;
wire  TCI ;
wire  tcj ;
wire  TCJ ;
wire  tck ;
wire  TCK ;
wire  tcm ;
wire  TCM ;
wire  tcn ;
wire  TCN ;
wire  tco ;
wire  TCO ;
wire  tcp ;
wire  TCP ;
wire  tea ;
wire  TEA ;
wire  teb ;
wire  TEB ;
wire  tec ;
wire  TEC ;
wire  ted ;
wire  TED ;
wire  tee ;
wire  TEE ;
wire  tei ;
wire  TEI ;
wire  tej ;
wire  TEJ ;
wire  tek ;
wire  TEK ;
wire  tem ;
wire  TEM ;
wire  ten ;
wire  TEN ;
wire  teo ;
wire  TEO ;
wire  tep ;
wire  TEP ;
wire  tga ;
wire  TGA ;
wire  tgb ;
wire  TGB ;
wire  tgc ;
wire  TGC ;
wire  tgd ;
wire  TGD ;
wire  tge ;
wire  TGE ;
wire  tgi ;
wire  TGI ;
wire  tgj ;
wire  TGJ ;
wire  tgk ;
wire  TGK ;
wire  tgm ;
wire  TGM ;
wire  tgn ;
wire  TGN ;
wire  tgo ;
wire  TGO ;
wire  tgp ;
wire  TGP ;
wire  ZZI ;
wire  ZZO ;
assign ZZI = 1'b1;
assign ZZO = 1'b0;
assign HAA = ~haa;  //complement 
assign HBA = ~hba;  //complement 
assign GAA =  QAE  ; 
assign gaa = ~GAA;  //complement  
assign GAE =  QAF  ; 
assign gae = ~GAE;  //complement 
assign HAB = ~hab;  //complement 
assign HBB = ~hbb;  //complement 
assign GAB =  QAE & HAA  ; 
assign gab = ~GAB;  //complement  
assign GAF =  QAF & HAE  ; 
assign gaf = ~GAF;  //complement 
assign HAC = ~hac;  //complement 
assign HBC = ~hbc;  //complement 
assign GAC =  QAE & HAA & HAB  ; 
assign gac = ~GAC;  //complement  
assign GAG =  QAF & HAE & HAF  ; 
assign gag = ~GAG;  //complement 
assign HAD = ~had;  //complement 
assign HBD = ~hbd;  //complement 
assign GAD =  QAE & HAA & HAB & HAC  ; 
assign gad = ~GAD;  //complement  
assign GAH =  QAF & HAE & HAF & HAG  ; 
assign gah = ~GAH;  //complement 
assign QAE = ~qae;  //complement 
assign QAF = ~qaf;  //complement 
assign HAE = ~hae;  //complement 
assign HBE = ~hbe;  //complement 
assign paa = ~PAA;  //complement 
assign pba = ~PBA;  //complement 
assign EAA = PBA; 
assign eaa = ~EAA; //complement 
assign EAB = PBA; 
assign eab = ~EAB;  //complement 
assign EAC = PBA; 
assign eac = ~EAC;  //complement 
assign EAD = PBA; 
assign ead = ~EAD;  //complement 
assign HAF = ~haf;  //complement 
assign HBF = ~hbf;  //complement 
assign pab = ~PAB;  //complement 
assign pbb = ~PBB;  //complement 
assign EAE = PBB; 
assign eae = ~EAE; //complement 
assign EAF = PBB; 
assign eaf = ~EAF;  //complement 
assign EAG = PBB; 
assign eag = ~EAG;  //complement 
assign EAH = PBB; 
assign eah = ~EAH;  //complement 
assign HAG = ~hag;  //complement 
assign HBG = ~hbg;  //complement 
assign eaq = pbd & pbb ; 
assign EAQ = ~eaq ; //complement 
assign ear = pbd & pbc ; 
assign EAR = ~ear ;  //complement 
assign pac = ~PAC;  //complement 
assign pbc = ~PBC;  //complement 
assign EAI = PBC; 
assign eai = ~EAI; //complement 
assign EAJ = PBC; 
assign eaj = ~EAJ;  //complement 
assign EAK = PBC; 
assign eak = ~EAK;  //complement 
assign EAL = PBC; 
assign eal = ~EAL;  //complement 
assign HAH = ~hah;  //complement 
assign HBH = ~hbh;  //complement 
assign jba = qai & gaa ; 
assign JBA = ~jba ; //complement 
assign JBB = qai & PAB ; 
assign jbb = ~JBB ;  //complement 
assign JBC = qai & PAC ; 
assign jbc = ~JBC ;  //complement 
assign JBD = qai & PAD; 
assign jbd = ~JBD; 
assign pad = ~PAD;  //complement 
assign pbd = ~PBD;  //complement 
assign EAM = PBD; 
assign eam = ~EAM; //complement 
assign EAN = PBD; 
assign ean = ~EAN;  //complement 
assign EAO = PBD; 
assign eao = ~EAO;  //complement 
assign EAP = PBD; 
assign eap = ~EAP;  //complement 
assign TAM = QAI; 
assign tam = ~TAM; //complement 
assign TAN = QAI; 
assign tan = ~TAN;  //complement 
assign TAO = QAI; 
assign tao = ~TAO;  //complement 
assign TAP = QAI; 
assign tap = ~TAP;  //complement 
assign JBE = qam & PAD ; 
assign jbe = ~JBE ; //complement 
assign JBF = qam & PAA ; 
assign jbf = ~JBF ;  //complement 
assign JBG = qam & PAB ; 
assign jbg = ~JBG ;  //complement 
assign JBH = qam & PAC; 
assign jbh = ~JBH; 
assign TAA =  QBA & QLA  |  QBB & QAC  |  QAL & QAP  |  QAM  ; 
assign taa = ~TAA;  //complement 
assign TAB =  QBA & QLA  |  QBB & QAC  |  QAL & QAP  |  QAM  ; 
assign tab = ~TAB; //complement 
assign TAC =  QBA & QLA  |  QBB & QAC  |  QAL & QAP  |  QAM  ; 
assign tac = ~TAC;  //complement 
assign kac = ~KAC;  //complement 
assign kad = ~KAD;  //complement 
assign kae = ~KAE;  //complement 
assign kaf = ~KAF;  //complement 
assign oba = ~OBA;  //complement 
assign obb = ~OBB;  //complement 
assign obi = ~OBI;  //complement 
assign obj = ~OBJ;  //complement 
assign obc = ~OBC;  //complement 
assign obd = ~OBD;  //complement 
assign obk = ~OBK;  //complement 
assign obl = ~OBL;  //complement 
assign oaa = ~OAA;  //complement 
assign oab = ~OAB;  //complement 
assign oac = ~OAC;  //complement 
assign oad = ~OAD;  //complement 
assign obe = ~OBE;  //complement 
assign obf = ~OBF;  //complement 
assign obm = ~OBM;  //complement 
assign obn = ~OBN;  //complement 
assign TAK =  AAA  ; 
assign tak = ~TAK;  //complement 
assign qam = ~QAM;  //complement 
assign obg = ~OBG;  //complement 
assign obh = ~OBH;  //complement 
assign obo = ~OBO;  //complement 
assign obp = ~OBP;  //complement 
assign AAC = ~aac;  //complement 
assign AAD = ~aad;  //complement 
assign AAA = ~aaa;  //complement 
assign AAB = ~aab;  //complement 
assign JAG =  LAA & lab & lac & lad & lae & laf  ; 
assign jag = ~JAG;  //complement  
assign JAA =  laa  ; 
assign jaa = ~JAA;  //complement 
assign laa = ~LAA;  //complement 
assign lba = ~LBA;  //complement 
assign oqa = ~OQA;  //complement 
assign qai = ~QAI;  //complement 
assign JAB =  LAB & LAA  |  lab & laa  ; 
assign jab = ~JAB; //complement 
assign lab = ~LAB;  //complement 
assign lbb = ~LBB;  //complement 
assign oai = ~OAI;  //complement 
assign oaj = ~OAJ;  //complement 
assign oak = ~OAK;  //complement 
assign oal = ~OAL;  //complement 
assign JAC =  LAC & LAA  |  LAC & KAC  |  lac & kac & laa  ; 
assign jac = ~JAC; //complement 
assign lac = ~LAC;  //complement 
assign lbc = ~LBC;  //complement 
assign oae = ~OAE;  //complement 
assign oaf = ~OAF;  //complement 
assign oag = ~OAG;  //complement 
assign oah = ~OAH;  //complement 
assign oam = ~OAM;  //complement 
assign oan = ~OAN;  //complement 
assign oao = ~OAO;  //complement 
assign oap = ~OAP;  //complement 
assign HAI = ~hai;  //complement 
assign HBI = ~hbi;  //complement 
assign GAI =  QAG  ; 
assign gai = ~GAI;  //complement  
assign GAM =  QAH  ; 
assign gam = ~GAM;  //complement 
assign HAJ = ~haj;  //complement 
assign HBJ = ~hbj;  //complement 
assign GAJ =  QAG & HAI  ; 
assign gaj = ~GAJ;  //complement  
assign GAN =  QAH & HAM  ; 
assign gan = ~GAN;  //complement 
assign HAK = ~hak;  //complement 
assign HBK = ~hbk;  //complement 
assign GAK =  QAG & HAI & HAJ  ; 
assign gak = ~GAK;  //complement  
assign GAO =  QAH & HAM & HAN  ; 
assign gao = ~GAO;  //complement 
assign HAL = ~hal;  //complement 
assign HBL = ~hbl;  //complement 
assign GAL =  QAG & HAI & HAJ & HAK  ; 
assign gal = ~GAL;  //complement  
assign GAP =  QAH & HAM & HAN & HAO  ; 
assign gap = ~GAP;  //complement 
assign QAG = ~qag;  //complement 
assign QAH = ~qah;  //complement 
assign HAM = ~ham;  //complement 
assign HBM = ~hbm;  //complement 
assign HAN = ~han;  //complement 
assign HBN = ~hbn;  //complement 
assign ofc = ~OFC;  //complement 
assign HAO = ~hao;  //complement 
assign HBO = ~hbo;  //complement 
assign HAP = ~hap;  //complement 
assign HBP = ~hbp;  //complement 
assign qap = ~QAP;  //complement 
assign TAD =  QBA & QLA  |  QBB & QAC  |  QAL & QAP  |  QAM  ; 
assign tad = ~TAD;  //complement 
assign TAE =  QBA & QLA  |  QBB & QAC  |  QAL & QAP  |  QAM  ; 
assign tae = ~TAE; //complement 
assign oem = ~OEM;  //complement 
assign oeo = ~OEO;  //complement 
assign oca = ~OCA;  //complement 
assign ocb = ~OCB;  //complement 
assign oci = ~OCI;  //complement 
assign ocj = ~OCJ;  //complement 
assign taj =  qaa & qab & qak  ; 
assign TAJ = ~taj;  //complement 
assign jah =  qal  |  QAJ  ; 
assign JAH = ~jah; //complement 
assign occ = ~OCC;  //complement 
assign ocd = ~OCD;  //complement 
assign ock = ~OCK;  //complement 
assign ocl = ~OCL;  //complement 
assign tai =  qaa & qab & qak  ; 
assign TAI = ~tai;  //complement 
assign oda = ~ODA;  //complement 
assign odb = ~ODB;  //complement 
assign odc = ~ODC;  //complement 
assign odd = ~ODD;  //complement 
assign oce = ~OCE;  //complement 
assign ocf = ~OCF;  //complement 
assign ocm = ~OCM;  //complement 
assign ocn = ~OCN;  //complement 
assign qaj = ~QAJ;  //complement 
assign qal = ~QAL;  //complement 
assign ocg = ~OCG;  //complement 
assign och = ~OCH;  //complement 
assign oco = ~OCO;  //complement 
assign ocp = ~OCP;  //complement 
assign qab = ~QAB;  //complement 
assign qbb = ~QBB;  //complement 
assign QAA = ~qaa;  //complement 
assign QBA = ~qba;  //complement 
assign QAN = ~qan;  //complement 
assign qac = ~QAC;  //complement 
assign JAD =  LAD & LBA  |  LAD & KAD  |  lad & kad & lba  ; 
assign jad = ~JAD; //complement 
assign lad = ~LAD;  //complement 
assign lbd = ~LBD;  //complement 
assign qad = ~QAD;  //complement 
assign qak = ~QAK;  //complement 
assign JAE =  LAE & LBA  |  LAE & KAE  |  lae & kae & lba  ; 
assign jae = ~JAE; //complement 
assign lae = ~LAE;  //complement 
assign lbe = ~LBE;  //complement 
assign odi = ~ODI;  //complement 
assign odj = ~ODJ;  //complement 
assign odk = ~ODK;  //complement 
assign odl = ~ODL;  //complement 
assign JAF =  LAF & LBA  |  LAF & KAF  |  laf & kaf & lba  ; 
assign jaf = ~JAF; //complement 
assign laf = ~LAF;  //complement 
assign ode = ~ODE;  //complement 
assign odf = ~ODF;  //complement 
assign odg = ~ODG;  //complement 
assign odh = ~ODH;  //complement 
assign odm = ~ODM;  //complement 
assign odn = ~ODN;  //complement 
assign odo = ~ODO;  //complement 
assign odp = ~ODP;  //complement 
assign HCA = ~hca;  //complement 
assign HDA = ~hda;  //complement 
assign GCA =  QCE  ; 
assign gca = ~GCA;  //complement  
assign GCE =  QCF  ; 
assign gce = ~GCE;  //complement 
assign HCB = ~hcb;  //complement 
assign HDB = ~hdb;  //complement 
assign GCB =  QCE & HCA  ; 
assign gcb = ~GCB;  //complement  
assign GCF =  QCF & HCE  ; 
assign gcf = ~GCF;  //complement 
assign HCC = ~hcc;  //complement 
assign HDC = ~hdc;  //complement 
assign GCC =  QCE & HCA & HCB  ; 
assign gcc = ~GCC;  //complement  
assign GCG =  QCF & HCE & HCF  ; 
assign gcg = ~GCG;  //complement 
assign HCD = ~hcd;  //complement 
assign HDD = ~hdd;  //complement 
assign GCD =  QCE & HCA & HCB & HCC  ; 
assign gcd = ~GCD;  //complement  
assign GCH =  QCF & HCE & HCF & HCG  ; 
assign gch = ~GCH;  //complement 
assign QCE = ~qce;  //complement 
assign QCF = ~qcf;  //complement 
assign HCE = ~hce;  //complement 
assign HDE = ~hde;  //complement 
assign HDG = ~hdg;  //complement 
assign pca = ~PCA;  //complement 
assign pda = ~PDA;  //complement 
assign ECA = PDA; 
assign eca = ~ECA; //complement 
assign ECB = PDA; 
assign ecb = ~ECB;  //complement 
assign ECC = PDA; 
assign ecc = ~ECC;  //complement 
assign ECD = PDA; 
assign ecd = ~ECD;  //complement 
assign HCF = ~hcf;  //complement 
assign HDF = ~hdf;  //complement 
assign HHM = ~hhm;  //complement 
assign pcb = ~PCB;  //complement 
assign pdb = ~PDB;  //complement 
assign ECE = PDB; 
assign ece = ~ECE; //complement 
assign ECF = PDB; 
assign ecf = ~ECF;  //complement 
assign ECG = PDB; 
assign ecg = ~ECG;  //complement 
assign ECH = PDB; 
assign ech = ~ECH;  //complement 
assign HCG = ~hcg;  //complement 
assign ecq = pdd & pdb ; 
assign ECQ = ~ecq ; //complement 
assign ecr = pdd & pdc ; 
assign ECR = ~ecr ;  //complement 
assign pcc = ~PCC;  //complement 
assign pdc = ~PDC;  //complement 
assign ECI = PDC; 
assign eci = ~ECI; //complement 
assign ECJ = PDC; 
assign ecj = ~ECJ;  //complement 
assign ECK = PDC; 
assign eck = ~ECK;  //complement 
assign ECL = PDC; 
assign ecl = ~ECL;  //complement 
assign HCH = ~hch;  //complement 
assign HDH = ~hdh;  //complement 
assign jda = qci & gca ; 
assign JDA = ~jda ; //complement 
assign JDB = qci & PCB ; 
assign jdb = ~JDB ;  //complement 
assign JDC = qci & PCC ; 
assign jdc = ~JDC ;  //complement 
assign JDD = qci & PCD; 
assign jdd = ~JDD; 
assign pcd = ~PCD;  //complement 
assign pdd = ~PDD;  //complement 
assign ECM = PDD; 
assign ecm = ~ECM; //complement 
assign ECN = PDD; 
assign ecn = ~ECN;  //complement 
assign ECO = PDD; 
assign eco = ~ECO;  //complement 
assign ECP = PDD; 
assign ecp = ~ECP;  //complement 
assign TCM = QCI; 
assign tcm = ~TCM; //complement 
assign TCN = QCI; 
assign tcn = ~TCN;  //complement 
assign TCO = QCI; 
assign tco = ~TCO;  //complement 
assign TCP = QCI; 
assign tcp = ~TCP;  //complement 
assign JDE = qcm & PCD ; 
assign jde = ~JDE ; //complement 
assign JDF = qcm & PCA ; 
assign jdf = ~JDF ;  //complement 
assign JDG = qcm & PCB ; 
assign jdg = ~JDG ;  //complement 
assign JDH = qcm & PCC; 
assign jdh = ~JDH; 
assign TCA =  QDA & QLA  |  QDB & QCC  |  QCL & QCP  |  QCM  ; 
assign tca = ~TCA;  //complement 
assign TCB =  QDA & QLA  |  QDB & QCC  |  QCL & QCP  |  QCM  ; 
assign tcb = ~TCB; //complement 
assign TCC =  QDA & QLA  |  QDB & QCC  |  QCL & QCP  |  QCM  ; 
assign tcc = ~TCC;  //complement 
assign kcc = ~KCC;  //complement 
assign kcd = ~KCD;  //complement 
assign kce = ~KCE;  //complement 
assign kcf = ~KCF;  //complement 
assign ofa = ~OFA;  //complement 
assign ofb = ~OFB;  //complement 
assign ofi = ~OFI;  //complement 
assign ofj = ~OFJ;  //complement 
assign ofd = ~OFD;  //complement 
assign ofk = ~OFK;  //complement 
assign ofl = ~OFL;  //complement 
assign oea = ~OEA;  //complement 
assign oeb = ~OEB;  //complement 
assign oec = ~OEC;  //complement 
assign oed = ~OED;  //complement 
assign ofe = ~OFE;  //complement 
assign off = ~OFF;  //complement 
assign ofm = ~OFM;  //complement 
assign ofn = ~OFN;  //complement 
assign TCK =  AAB  ; 
assign tck = ~TCK;  //complement 
assign qcm = ~QCM;  //complement 
assign ofg = ~OFG;  //complement 
assign ofh = ~OFH;  //complement 
assign ofo = ~OFO;  //complement 
assign ofp = ~OFP;  //complement 
assign QLA = ~qla;  //complement 
assign QLB = ~qlb;  //complement 
assign QJA = ~qja;  //complement 
assign QKB = ~qkb;  //complement 
assign JCG =  LCA & lcb & lcc & lcd & lce & lcf  ; 
assign jcg = ~JCG;  //complement  
assign JCA =  lca  ; 
assign jca = ~JCA;  //complement 
assign lca = ~LCA;  //complement 
assign lda = ~LDA;  //complement 
assign oqb = ~OQB;  //complement 
assign qci = ~QCI;  //complement 
assign JCB =  LCB & LCA  |  lcb & lca  ; 
assign jcb = ~JCB; //complement 
assign lcb = ~LCB;  //complement 
assign ldb = ~LDB;  //complement 
assign oei = ~OEI;  //complement 
assign oej = ~OEJ;  //complement 
assign oek = ~OEK;  //complement 
assign oel = ~OEL;  //complement 
assign JCC =  LCC & LCA  |  LCC & KCC  |  lcc & kcc & lca  ; 
assign jcc = ~JCC; //complement 
assign lcc = ~LCC;  //complement 
assign ldc = ~LDC;  //complement 
assign oee = ~OEE;  //complement 
assign oef = ~OEF;  //complement 
assign oeg = ~OEG;  //complement 
assign oeh = ~OEH;  //complement 
assign oen = ~OEN;  //complement 
assign oep = ~OEP;  //complement 
assign HCI = ~hci;  //complement 
assign HDI = ~hdi;  //complement 
assign GCI =  QCG  ; 
assign gci = ~GCI;  //complement  
assign GCM =  QCH  ; 
assign gcm = ~GCM;  //complement 
assign HCJ = ~hcj;  //complement 
assign HDJ = ~hdj;  //complement 
assign GCJ =  QCG & HCI  ; 
assign gcj = ~GCJ;  //complement  
assign GCN =  QCH & HCM  ; 
assign gcn = ~GCN;  //complement 
assign HCK = ~hck;  //complement 
assign HDK = ~hdk;  //complement 
assign GCK =  QCG & HCI & HCJ  ; 
assign gck = ~GCK;  //complement  
assign GCO =  QCH & HCM & HCN  ; 
assign gco = ~GCO;  //complement 
assign HCL = ~hcl;  //complement 
assign HDL = ~hdl;  //complement 
assign GCL =  QCG & HCI & HCJ & HCK  ; 
assign gcl = ~GCL;  //complement  
assign GCP =  QCH & HCM & HCN & HCO  ; 
assign gcp = ~GCP;  //complement 
assign QCG = ~qcg;  //complement 
assign QCH = ~qch;  //complement 
assign HCM = ~hcm;  //complement 
assign HDM = ~hdm;  //complement 
assign HCN = ~hcn;  //complement 
assign HDN = ~hdn;  //complement 
assign HCO = ~hco;  //complement 
assign HDO = ~hdo;  //complement 
assign HCP = ~hcp;  //complement 
assign HDP = ~hdp;  //complement 
assign qcp = ~QCP;  //complement 
assign TCD =  QDA & QLA  |  QDB & QCC  |  QCL & QCP  |  QCM  ; 
assign tcd = ~TCD;  //complement 
assign TCE =  QDA & QLA  |  QDB & QCC  |  QCL & QCP  |  QCM  ; 
assign tce = ~TCE; //complement 
assign oga = ~OGA;  //complement 
assign ogb = ~OGB;  //complement 
assign ogi = ~OGI;  //complement 
assign ogj = ~OGJ;  //complement 
assign jch =  qcl  |  QCJ  ; 
assign JCH = ~jch; //complement 
assign qck = ~QCK;  //complement 
assign ogc = ~OGC;  //complement 
assign ogd = ~OGD;  //complement 
assign ogk = ~OGK;  //complement 
assign ogl = ~OGL;  //complement 
assign tci =  qca & qcb & qck  ; 
assign TCI = ~tci;  //complement 
assign tcj =  qca & qcb & qck  ; 
assign TCJ = ~tcj;  //complement 
assign oha = ~OHA;  //complement 
assign ohb = ~OHB;  //complement 
assign ohc = ~OHC;  //complement 
assign ohd = ~OHD;  //complement 
assign oge = ~OGE;  //complement 
assign ogf = ~OGF;  //complement 
assign ogm = ~OGM;  //complement 
assign ogn = ~OGN;  //complement 
assign qcj = ~QCJ;  //complement 
assign qcl = ~QCL;  //complement 
assign ogg = ~OGG;  //complement 
assign ogh = ~OGH;  //complement 
assign ogo = ~OGO;  //complement 
assign ogp = ~OGP;  //complement 
assign qcb = ~QCB;  //complement 
assign qdb = ~QDB;  //complement 
assign QCA = ~qca;  //complement 
assign QDA = ~qda;  //complement 
assign QCN = ~qcn;  //complement 
assign qcc = ~QCC;  //complement 
assign JCD =  LCD & LDA  |  LCD & KCD  |  lcd & kcd & lda  ; 
assign jcd = ~JCD; //complement 
assign lcd = ~LCD;  //complement 
assign ldd = ~LDD;  //complement 
assign qcd = ~QCD;  //complement 
assign JCE =  LCE & LDA  |  LCE & KCE  |  lce & kce & lda  ; 
assign jce = ~JCE; //complement 
assign lce = ~LCE;  //complement 
assign lde = ~LDE;  //complement 
assign ohi = ~OHI;  //complement 
assign ohj = ~OHJ;  //complement 
assign ohk = ~OHK;  //complement 
assign ohl = ~OHL;  //complement 
assign JCF =  LCF & LDA  |  LCF & KCF  |  lcf & kcf & lda  ; 
assign jcf = ~JCF; //complement 
assign lcf = ~LCF;  //complement 
assign ohe = ~OHE;  //complement 
assign ohf = ~OHF;  //complement 
assign ohg = ~OHG;  //complement 
assign ohh = ~OHH;  //complement 
assign ohm = ~OHM;  //complement 
assign ohn = ~OHN;  //complement 
assign oho = ~OHO;  //complement 
assign ohp = ~OHP;  //complement 
assign HEA = ~hea;  //complement 
assign HFA = ~hfa;  //complement 
assign GEA =  QEE  ; 
assign gea = ~GEA;  //complement  
assign GEE =  QEF  ; 
assign gee = ~GEE;  //complement 
assign HEB = ~heb;  //complement 
assign HFB = ~hfb;  //complement 
assign GEB =  QEE & HEA  ; 
assign geb = ~GEB;  //complement  
assign GEF =  QEF & HEE  ; 
assign gef = ~GEF;  //complement 
assign HHO = ~hho;  //complement 
assign HEC = ~hec;  //complement 
assign HFC = ~hfc;  //complement 
assign GEC =  QEE & HEA & HEB  ; 
assign gec = ~GEC;  //complement  
assign GEG =  QEF & HEE & HEF  ; 
assign geg = ~GEG;  //complement 
assign HED = ~hed;  //complement 
assign HFD = ~hfd;  //complement 
assign GED =  QEE & HEA & HEB & HEC  ; 
assign ged = ~GED;  //complement  
assign GEH =  QEF & HEE & HEF & HEG  ; 
assign geh = ~GEH;  //complement 
assign QEE = ~qee;  //complement 
assign QEF = ~qef;  //complement 
assign HEE = ~hee;  //complement 
assign HFE = ~hfe;  //complement 
assign pea = ~PEA;  //complement 
assign pfa = ~PFA;  //complement 
assign EEA = PFA; 
assign eea = ~EEA; //complement 
assign EEB = PFA; 
assign eeb = ~EEB;  //complement 
assign EEC = PFA; 
assign eec = ~EEC;  //complement 
assign EED = PFA; 
assign eed = ~EED;  //complement 
assign HEF = ~hef;  //complement 
assign HFF = ~hff;  //complement 
assign eeq = pfd & pfb ; 
assign EEQ = ~eeq ; //complement 
assign eer = pfd & pfc ; 
assign EER = ~eer ;  //complement 
assign peb = ~PEB;  //complement 
assign pfb = ~PFB;  //complement 
assign EEE = PFB; 
assign eee = ~EEE; //complement 
assign EEF = PFB; 
assign eef = ~EEF;  //complement 
assign EEG = PFB; 
assign eeg = ~EEG;  //complement 
assign EEH = PFB; 
assign eeh = ~EEH;  //complement 
assign HEG = ~heg;  //complement 
assign HFG = ~hfg;  //complement 
assign pec = ~PEC;  //complement 
assign pfc = ~PFC;  //complement 
assign EEI = PFC; 
assign eei = ~EEI; //complement 
assign EEJ = PFC; 
assign eej = ~EEJ;  //complement 
assign EEK = PFC; 
assign eek = ~EEK;  //complement 
assign EEL = PFC; 
assign eel = ~EEL;  //complement 
assign HEH = ~heh;  //complement 
assign HFH = ~hfh;  //complement 
assign jfa = qei & gea ; 
assign JFA = ~jfa ; //complement 
assign JFB = qei & PEB ; 
assign jfb = ~JFB ;  //complement 
assign JFC = qei & PEC ; 
assign jfc = ~JFC ;  //complement 
assign JFD = qei & PED; 
assign jfd = ~JFD; 
assign ped = ~PED;  //complement 
assign pfd = ~PFD;  //complement 
assign EEM = PFD; 
assign eem = ~EEM; //complement 
assign EEN = PFD; 
assign een = ~EEN;  //complement 
assign EEO = PFD; 
assign eeo = ~EEO;  //complement 
assign EEP = PFD; 
assign eep = ~EEP;  //complement 
assign TEM = QEI; 
assign tem = ~TEM; //complement 
assign TEN = QEI; 
assign ten = ~TEN;  //complement 
assign TEO = QEI; 
assign teo = ~TEO;  //complement 
assign TEP = QEI; 
assign tep = ~TEP;  //complement 
assign JFE = qem & PED ; 
assign jfe = ~JFE ; //complement 
assign JFF = qem & PEA ; 
assign jff = ~JFF ;  //complement 
assign JFG = qem & PEB ; 
assign jfg = ~JFG ;  //complement 
assign JFH = qem & PEC; 
assign jfh = ~JFH; 
assign TEA =  QFA & QLB  |  QFB & QEC  |  QEL & QEP  |  QEM  ; 
assign tea = ~TEA;  //complement 
assign TEB =  QFA & QLB  |  QFB & QEC  |  QEL & QEP  |  QEM  ; 
assign teb = ~TEB; //complement 
assign TEC =  QFA & QLB  |  QFB & QEC  |  QEL & QEP  |  QEM  ; 
assign tec = ~TEC;  //complement 
assign kec = ~KEC;  //complement 
assign ked = ~KED;  //complement 
assign kee = ~KEE;  //complement 
assign kef = ~KEF;  //complement 
assign oja = ~OJA;  //complement 
assign ojb = ~OJB;  //complement 
assign oji = ~OJI;  //complement 
assign ojj = ~OJJ;  //complement 
assign ojc = ~OJC;  //complement 
assign ojd = ~OJD;  //complement 
assign ojk = ~OJK;  //complement 
assign ojl = ~OJL;  //complement 
assign oia = ~OIA;  //complement 
assign oib = ~OIB;  //complement 
assign oic = ~OIC;  //complement 
assign oid = ~OID;  //complement 
assign ojf = ~OJF;  //complement 
assign oje = ~OJE;  //complement 
assign ojm = ~OJM;  //complement 
assign ojn = ~OJN;  //complement 
assign TEK =  AAC  ; 
assign tek = ~TEK;  //complement 
assign qem = ~QEM;  //complement 
assign ojg = ~OJG;  //complement 
assign ojh = ~OJH;  //complement 
assign ojo = ~OJO;  //complement 
assign ojp = ~OJP;  //complement 
assign ABA = ~aba;  //complement 
assign ABB = ~abb;  //complement 
assign ABC = ~abc;  //complement 
assign ABD = ~abd;  //complement 
assign JEG =  LEA & leb & lec & led & lee & lef  ; 
assign jeg = ~JEG;  //complement  
assign JEA =  lea  ; 
assign jea = ~JEA;  //complement 
assign lea = ~LEA;  //complement 
assign lfa = ~LFA;  //complement 
assign oqc = ~OQC;  //complement 
assign qei = ~QEI;  //complement 
assign JEB =  LEB & LEA  |  leb & lea  ; 
assign jeb = ~JEB; //complement 
assign leb = ~LEB;  //complement 
assign lfb = ~LFB;  //complement 
assign oii = ~OII;  //complement 
assign oij = ~OIJ;  //complement 
assign oik = ~OIK;  //complement 
assign oil = ~OIL;  //complement 
assign JEC =  LEC & LEA  |  LEC & KEC  |  lec & kec & lea  ; 
assign jec = ~JEC; //complement 
assign lec = ~LEC;  //complement 
assign lfc = ~LFC;  //complement 
assign oie = ~OIE;  //complement 
assign oif = ~OIF;  //complement 
assign oig = ~OIG;  //complement 
assign oih = ~OIH;  //complement 
assign oim = ~OIM;  //complement 
assign oin = ~OIN;  //complement 
assign oio = ~OIO;  //complement 
assign oip = ~OIP;  //complement 
assign HEI = ~hei;  //complement 
assign HFI = ~hfi;  //complement 
assign GEI =  QEG  ; 
assign gei = ~GEI;  //complement  
assign GEM =  QEH  ; 
assign gem = ~GEM;  //complement 
assign HEJ = ~hej;  //complement 
assign HFJ = ~hfj;  //complement 
assign GEJ =  QEG & HEI  ; 
assign gej = ~GEJ;  //complement  
assign GEN =  QEH & HEM  ; 
assign gen = ~GEN;  //complement 
assign HEK = ~hek;  //complement 
assign HFK = ~hfk;  //complement 
assign GEK =  QEG & HEI & HEJ  ; 
assign gek = ~GEK;  //complement  
assign GEO =  QEH & HEM & HEN  ; 
assign geo = ~GEO;  //complement 
assign HEL = ~hel;  //complement 
assign HFL = ~hfl;  //complement 
assign GEL =  QEG & HEI & HEJ & HEK  ; 
assign gel = ~GEL;  //complement  
assign GEP =  QEH & HEM & HEN & HEO  ; 
assign gep = ~GEP;  //complement 
assign QEG = ~qeg;  //complement 
assign QEH = ~qeh;  //complement 
assign HEM = ~hem;  //complement 
assign HFM = ~hfm;  //complement 
assign HEN = ~hen;  //complement 
assign HFN = ~hfn;  //complement 
assign HEO = ~heo;  //complement 
assign HFO = ~hfo;  //complement 
assign HEP = ~hep;  //complement 
assign HFP = ~hfp;  //complement 
assign qep = ~QEP;  //complement 
assign TED =  QFA & QLB  |  QFB & QEC  |  QEL & QEP  |  QEM  ; 
assign ted = ~TED;  //complement 
assign TEE =  QFA & QLB  |  QFB & QEC  |  QEL & QEP  |  QEM  ; 
assign tee = ~TEE; //complement 
assign oka = ~OKA;  //complement 
assign okb = ~OKB;  //complement 
assign oki = ~OKI;  //complement 
assign okj = ~OKJ;  //complement 
assign okc = ~OKC;  //complement 
assign okd = ~OKD;  //complement 
assign okk = ~OKK;  //complement 
assign okl = ~OKL;  //complement 
assign tei =  qea & qeb & qek  ; 
assign TEI = ~tei;  //complement 
assign tej =  qea & qeb & qek  ; 
assign TEJ = ~tej;  //complement 
assign jeh =  qel  |  QEJ  ; 
assign JEH = ~jeh; //complement 
assign oke = ~OKE;  //complement 
assign okf = ~OKF;  //complement 
assign okm = ~OKM;  //complement 
assign okn = ~OKN;  //complement 
assign qej = ~QEJ;  //complement 
assign qek = ~QEK;  //complement 
assign qel = ~QEL;  //complement 
assign okg = ~OKG;  //complement 
assign okh = ~OKH;  //complement 
assign oko = ~OKO;  //complement 
assign okp = ~OKP;  //complement 
assign qeb = ~QEB;  //complement 
assign qfb = ~QFB;  //complement 
assign QEA = ~qea;  //complement 
assign QFA = ~qfa;  //complement 
assign QEN = ~qen;  //complement 
assign qna = ~QNA;  //complement 
assign qec = ~QEC;  //complement 
assign JED =  LED & LFA  |  LED & KED  |  led & ked & lfa  ; 
assign jed = ~JED; //complement 
assign led = ~LED;  //complement 
assign lfd = ~LFD;  //complement 
assign qed = ~QED;  //complement 
assign JEE =  LEE & LFA  |  LEE & KEE  |  lee & kee & lfa  ; 
assign jee = ~JEE; //complement 
assign lee = ~LEE;  //complement 
assign lfe = ~LFE;  //complement 
assign ola = ~OLA;  //complement 
assign olb = ~OLB;  //complement 
assign olc = ~OLC;  //complement 
assign old = ~OLD;  //complement 
assign oli = ~OLI;  //complement 
assign olj = ~OLJ;  //complement 
assign olk = ~OLK;  //complement 
assign oll = ~OLL;  //complement 
assign JEF =  LEF & LFA  |  LEF & KEF  |  lef & kef & lfa  ; 
assign jef = ~JEF; //complement 
assign lef = ~LEF;  //complement 
assign ole = ~OLE;  //complement 
assign olf = ~OLF;  //complement 
assign olg = ~OLG;  //complement 
assign olh = ~OLH;  //complement 
assign olm = ~OLM;  //complement 
assign oln = ~OLN;  //complement 
assign olo = ~OLO;  //complement 
assign olp = ~OLP;  //complement 
assign HGA = ~hga;  //complement 
assign HHA = ~hha;  //complement 
assign GGA =  QGE  ; 
assign gga = ~GGA;  //complement  
assign GGE =  QGF  ; 
assign gge = ~GGE;  //complement 
assign HGB = ~hgb;  //complement 
assign HHB = ~hhb;  //complement 
assign GGB =  QGE & HGA  ; 
assign ggb = ~GGB;  //complement  
assign GGF =  QGF & HGE  ; 
assign ggf = ~GGF;  //complement 
assign HGC = ~hgc;  //complement 
assign HHC = ~hhc;  //complement 
assign GGC =  QGE & HGA & HGB  ; 
assign ggc = ~GGC;  //complement  
assign GGG =  QGF & HGE & HGF  ; 
assign ggg = ~GGG;  //complement 
assign HGD = ~hgd;  //complement 
assign HHD = ~hhd;  //complement 
assign GGD =  QGE & HGA & HGB & HGC  ; 
assign ggd = ~GGD;  //complement  
assign GGH =  QGF & HGE & HGF & HGG  ; 
assign ggh = ~GGH;  //complement 
assign QGE = ~qge;  //complement 
assign QGF = ~qgf;  //complement 
assign HGE = ~hge;  //complement 
assign HHE = ~hhe;  //complement 
assign pga = ~PGA;  //complement 
assign pha = ~PHA;  //complement 
assign EGA = PHA; 
assign ega = ~EGA; //complement 
assign EGB = PHA; 
assign egb = ~EGB;  //complement 
assign EGC = PHA; 
assign egc = ~EGC;  //complement 
assign EGD = PHA; 
assign egd = ~EGD;  //complement 
assign HGF = ~hgf;  //complement 
assign HHF = ~hhf;  //complement 
assign pgb = ~PGB;  //complement 
assign phb = ~PHB;  //complement 
assign EGE = PHB; 
assign ege = ~EGE; //complement 
assign EGF = PHB; 
assign egf = ~EGF;  //complement 
assign EGG = PHB; 
assign egg = ~EGG;  //complement 
assign EGH = PHB; 
assign egh = ~EGH;  //complement 
assign HGG = ~hgg;  //complement 
assign HHG = ~hhg;  //complement 
assign egq = phd & phb ; 
assign EGQ = ~egq ; //complement 
assign egr = phd & phc ; 
assign EGR = ~egr ;  //complement 
assign pgc = ~PGC;  //complement 
assign phc = ~PHC;  //complement 
assign EGI = PHC; 
assign egi = ~EGI; //complement 
assign EGJ = PHC; 
assign egj = ~EGJ;  //complement 
assign EGK = PHC; 
assign egk = ~EGK;  //complement 
assign EGL = PHC; 
assign egl = ~EGL;  //complement 
assign HGH = ~hgh;  //complement 
assign HHH = ~hhh;  //complement 
assign jha = qgi & gga ; 
assign JHA = ~jha ; //complement 
assign JHB = qgi & PGB ; 
assign jhb = ~JHB ;  //complement 
assign JHC = qgi & PGC ; 
assign jhc = ~JHC ;  //complement 
assign JHD = qgi & PGD; 
assign jhd = ~JHD; 
assign pgd = ~PGD;  //complement 
assign phd = ~PHD;  //complement 
assign EGM = PHD; 
assign egm = ~EGM; //complement 
assign EGN = PHD; 
assign egn = ~EGN;  //complement 
assign EGO = PHD; 
assign ego = ~EGO;  //complement 
assign EGP = PHD; 
assign egp = ~EGP;  //complement 
assign TGM = QGI; 
assign tgm = ~TGM; //complement 
assign TGN = QGI; 
assign tgn = ~TGN;  //complement 
assign TGO = QGI; 
assign tgo = ~TGO;  //complement 
assign TGP = QGI; 
assign tgp = ~TGP;  //complement 
assign JHE = qgm & PGD ; 
assign jhe = ~JHE ; //complement 
assign JHF = qgm & PGA ; 
assign jhf = ~JHF ;  //complement 
assign JHG = qgm & PGB ; 
assign jhg = ~JHG ;  //complement 
assign JHH = qgm & PGC; 
assign jhh = ~JHH; 
assign TGA =  QHA & QLB  |  QHB & QGC  |  QGL & QGP  |  QGM  ; 
assign tga = ~TGA;  //complement 
assign TGB =  QHA & QLB  |  QHB & QGC  |  QGL & QGP  |  QGM  ; 
assign tgb = ~TGB; //complement 
assign TGC =  QHA & QLB  |  QHB & QGC  |  QGL & QGP  |  QGM  ; 
assign tgc = ~TGC;  //complement 
assign kgc = ~KGC;  //complement 
assign kge = ~KGE;  //complement 
assign kgd = ~KGD;  //complement 
assign kgf = ~KGF;  //complement 
assign ona = ~ONA;  //complement 
assign onb = ~ONB;  //complement 
assign oni = ~ONI;  //complement 
assign onj = ~ONJ;  //complement 
assign onc = ~ONC;  //complement 
assign ond = ~OND;  //complement 
assign onk = ~ONK;  //complement 
assign onl = ~ONL;  //complement 
assign one = ~ONE;  //complement 
assign onf = ~ONF;  //complement 
assign onm = ~ONM;  //complement 
assign onn = ~ONN;  //complement 
assign TGK =  AAD  ; 
assign tgk = ~TGK;  //complement 
assign qgm = ~QGM;  //complement 
assign ong = ~ONG;  //complement 
assign onh = ~ONH;  //complement 
assign ono = ~ONO;  //complement 
assign onp = ~ONP;  //complement 
assign qka = ~QKA;  //complement 
assign JGG =  LGA & lgb & lgc & lgd & lge & lgf  ; 
assign jgg = ~JGG;  //complement  
assign JGA =  lga  ; 
assign jga = ~JGA;  //complement 
assign lga = ~LGA;  //complement 
assign lha = ~LHA;  //complement 
assign qia = ~QIA;  //complement 
assign oqd = ~OQD;  //complement 
assign qgi = ~QGI;  //complement 
assign JGB =  LGB & LGA  |  lgb & lga  ; 
assign jgb = ~JGB; //complement 
assign lgb = ~LGB;  //complement 
assign lhb = ~LHB;  //complement 
assign oma = ~OMA;  //complement 
assign omb = ~OMB;  //complement 
assign omc = ~OMC;  //complement 
assign omd = ~OMD;  //complement 
assign omi = ~OMI;  //complement 
assign omj = ~OMJ;  //complement 
assign omk = ~OMK;  //complement 
assign oml = ~OML;  //complement 
assign JGC =  LGC & LGA  |  LGC & KGC  |  lgc & kgc & lga  ; 
assign jgc = ~JGC; //complement 
assign lgc = ~LGC;  //complement 
assign lhc = ~LHC;  //complement 
assign ome = ~OME;  //complement 
assign omf = ~OMF;  //complement 
assign omg = ~OMG;  //complement 
assign omh = ~OMH;  //complement 
assign omm = ~OMM;  //complement 
assign omn = ~OMN;  //complement 
assign omo = ~OMO;  //complement 
assign omp = ~OMP;  //complement 
assign HGI = ~hgi;  //complement 
assign HHI = ~hhi;  //complement 
assign GGI =  QGG  ; 
assign ggi = ~GGI;  //complement  
assign GGM =  QGH  ; 
assign ggm = ~GGM;  //complement 
assign HHN = ~hhn;  //complement 
assign HGJ = ~hgj;  //complement 
assign HHJ = ~hhj;  //complement 
assign GGJ =  QGG & HGI  ; 
assign ggj = ~GGJ;  //complement  
assign GGN =  QGH & HGM  ; 
assign ggn = ~GGN;  //complement 
assign HGK = ~hgk;  //complement 
assign HHK = ~hhk;  //complement 
assign GGK =  QGG & HGI & HGJ  ; 
assign ggk = ~GGK;  //complement  
assign GGO =  QGH & HGM & HGN  ; 
assign ggo = ~GGO;  //complement 
assign HGL = ~hgl;  //complement 
assign HHL = ~hhl;  //complement 
assign GGL =  QGG & HGI & HGJ & HGK  ; 
assign ggl = ~GGL;  //complement  
assign GGP =  QGH & HGM & HGN & HGO  ; 
assign ggp = ~GGP;  //complement 
assign QGG = ~qgg;  //complement 
assign QGH = ~qgh;  //complement 
assign HGM = ~hgm;  //complement 
assign HGN = ~hgn;  //complement 
assign HGO = ~hgo;  //complement 
assign HGP = ~hgp;  //complement 
assign HHP = ~hhp;  //complement 
assign qgp = ~QGP;  //complement 
assign TGD =  QHA & QLB  |  QHB & QGC  |  QGL & QGP  |  QGM  ; 
assign tgd = ~TGD;  //complement 
assign TGE =  QHA & QLB  |  QHB & QGC  |  QGL & QGP  |  QGM  ; 
assign tge = ~TGE; //complement 
assign ooa = ~OOA;  //complement 
assign oob = ~OOB;  //complement 
assign ooi = ~OOI;  //complement 
assign ooj = ~OOJ;  //complement 
assign tgi =  qga & qgb & qgk  ; 
assign TGI = ~tgi;  //complement 
assign tgj =  qga & qgb & qgk  ; 
assign TGJ = ~tgj;  //complement 
assign qgk = ~QGK;  //complement 
assign ooc = ~OOC;  //complement 
assign ood = ~OOD;  //complement 
assign ook = ~OOK;  //complement 
assign ool = ~OOL;  //complement 
assign jgh =  qgl  |  QGJ  ; 
assign JGH = ~jgh; //complement 
assign opa = ~OPA;  //complement 
assign opb = ~OPB;  //complement 
assign opc = ~OPC;  //complement 
assign opd = ~OPD;  //complement 
assign ooe = ~OOE;  //complement 
assign oof = ~OOF;  //complement 
assign oom = ~OOM;  //complement 
assign oon = ~OON;  //complement 
assign qgj = ~QGJ;  //complement 
assign qgl = ~QGL;  //complement 
assign oog = ~OOG;  //complement 
assign ooh = ~OOH;  //complement 
assign ooo = ~OOO;  //complement 
assign oop = ~OOP;  //complement 
assign qgb = ~QGB;  //complement 
assign qhb = ~QHB;  //complement 
assign QGA = ~qga;  //complement 
assign QHA = ~qha;  //complement 
assign QGN = ~qgn;  //complement 
assign qgc = ~QGC;  //complement 
assign JGD =  LGD & LHA  |  LGD & KGD  |  lgd & kgd & lha  ; 
assign jgd = ~JGD; //complement 
assign lgd = ~LGD;  //complement 
assign lhd = ~LHD;  //complement 
assign qgd = ~QGD;  //complement 
assign qnb = ~QNB;  //complement 
assign JGE =  LGE & LHA  |  LGE & KGE  |  lge & kge & lha  ; 
assign jge = ~JGE; //complement 
assign lge = ~LGE;  //complement 
assign lhe = ~LHE;  //complement 
assign opi = ~OPI;  //complement 
assign opj = ~OPJ;  //complement 
assign opk = ~OPK;  //complement 
assign opl = ~OPL;  //complement 
assign JGF =  LGF & LHA  |  LGF & KGF  |  lgf & kgf & lha  ; 
assign jgf = ~JGF; //complement 
assign lgf = ~LGF;  //complement 
assign ope = ~OPE;  //complement 
assign opf = ~OPF;  //complement 
assign opg = ~OPG;  //complement 
assign oph = ~OPH;  //complement 
assign opm = ~OPM;  //complement 
assign opn = ~OPN;  //complement 
assign opo = ~OPO;  //complement 
assign opp = ~OPP;  //complement 
assign iaa = ~IAA; //complement 
assign iab = ~IAB; //complement 
assign iba = ~IBA; //complement 
assign ibb = ~IBB; //complement 
assign ibc = ~IBC; //complement 
assign ibd = ~IBD; //complement 
assign ibe = ~IBE; //complement 
assign ica = ~ICA; //complement 
assign icb = ~ICB; //complement 
assign ida = ~IDA; //complement 
assign idb = ~IDB; //complement 
assign idc = ~IDC; //complement 
assign idd = ~IDD; //complement 
assign iea = ~IEA; //complement 
assign ieb = ~IEB; //complement 
assign iec = ~IEC; //complement 
assign ied = ~IED; //complement 
assign iee = ~IEE; //complement 
assign ifa = ~IFA; //complement 
assign ifb = ~IFB; //complement 
assign ifc = ~IFC; //complement 
assign ifd = ~IFD; //complement 
assign ife = ~IFE; //complement 
assign ifff  = ~IFFF ; //complement 
assign iga = ~IGA; //complement 
assign iha = ~IHA; //complement 
assign ihb = ~IHB; //complement 
assign izz = ~IZZ; //complement 
always@(posedge IZZ )
   begin 
 haa <=  haa & gaa  |  HAA & GAA  |  TAM  ; 
 hba <=  haa & gaa  |  HAA & GAA  |  TAM  ; 
 hab <=  hab & gab  |  HAB & GAB  |  TAM  ; 
 hbb <=  hab & gab  |  HAB & GAB  |  TAM  ; 
 hac <=  hac & gac  |  HAC & GAC  |  TAM  ; 
 hbc <=  hac & gac  |  HAC & GAC  |  TAM  ; 
 had <=  had & gad  |  HAD & GAD  |  TAM  ; 
 hbd <=  had & gad  |  HAD & GAD  |  TAM  ; 
 qae <=  tac  |  paa  ; 
 qaf <=  tac  |  pab  ; 
 hae <=  hae & gae  |  HAE & GAE  |  TAN  ; 
 hbe <=  hae & gae  |  HAE & GAE  |  TAN  ; 
 PAA <=  JBA & tak & taa  |  ABA & TAK  |  JBE & TAA  ; 
 PBA <=  JBA & tak & taa  |  ABA & TAK  |  JBE & TAA  ; 
 haf <=  haf & gaf  |  HAF & GAF  |  TAN  ; 
 hbf <=  haf & gaf  |  HAF & GAF  |  TAN  ; 
 PAB <=  JBB & tak & taa  |  ABB & TAK  |  JBF & TAA  ; 
 PBB <=  JBB & tak & taa  |  ABB & TAK  |  JBF & TAA  ; 
 hag <=  hag & gag  |  HAG & GAG  |  TAN  ; 
 hbg <=  hag & gag  |  HAG & GAG  |  TAN  ; 
 PAC <=  JBC & tak & taa  |  ABC & TAK  |  JBG & TAA  ; 
 PBC <=  JBC & tak & taa  |  ABC & TAK  |  JBG & TAA  ; 
 hah <=  hah & gah  |  HAH & GAH  |  TAN  ; 
 hbh <=  hah & gah  |  HAH & GAH  |  TAN  ; 
 PAD <=  JBD & tak & taa  |  ABD & TAK  |  JBH & TAA  ; 
 PBD <=  JBD & tak & taa  |  ABD & TAK  |  JBH & TAA  ; 
 KAC <= LBB ; 
 KAD <=  LBB  |  LBC  ; 
 KAE <=  LBB  |  LBC  |  LBD  ; 
 KAF <=  LBB  |  LBC  |  LBD  |  LBE  ; 
 OBA <=  HBA & EAA  |  HBE & EAE  |  HBI & EAI  |  HBM & EAM  ; 
 OBB <=  HBA & EAA  |  HBE & EAE  |  HBI & EAI  |  HBM & EAM  ; 
 OBI <=  HBB & EAB  |  HBF & EAF  |  HBJ & EAJ  |  HBN & EAN  ; 
 OBJ <=  HBB & EAB  |  HBF & EAF  |  HBJ & EAJ  |  HBN & EAN  ; 
 OBC <=  HBA & EAA  |  HBE & EAE  |  HBI & EAI  |  HBM & EAM  ; 
 OBD <=  HBA & EAA  |  HBE & EAE  |  HBI & EAI  |  HBM & EAM  ; 
 OBK <=  HBB & EAB  |  HBF & EAF  |  HBJ & EAJ  |  HBN & EAN  ; 
 OBL <=  HBB & EAB  |  HBF & EAF  |  HBJ & EAJ  |  HBN & EAN  ; 
 OAA <= EAQ ; 
 OAB <= EAQ ; 
 OAC <= EAQ ; 
 OAD <= EAQ ; 
 OBE <=  HBA & EAA  |  HBE & EAE  |  HBI & EAI  |  HBM & EAM  ; 
 OBF <=  HBA & EAA  |  HBE & EAE  |  HBI & EAI  |  HBM & EAM  ; 
 OBM <=  HBB & EAB  |  HBF & EAF  |  HBJ & EAJ  |  HBN & EAN  ; 
 OBN <=  HBB & EAB  |  HBF & EAF  |  HBJ & EAJ  |  HBN & EAN  ; 
 QAM <= AAA ; 
 OBG <=  HBA & EAA  |  HBE & EAE  |  HBI & EAI  |  HBM & EAM  ; 
 OBH <=  HBA & EAA  |  HBE & EAE  |  HBI & EAI  |  HBM & EAM  ; 
 OBO <=  HBB & EAB  |  HBF & EAF  |  HBJ & EAJ  |  HBN & EAN  ; 
 OBP <=  HBB & EAB  |  HBF & EAF  |  HBJ & EAJ  |  HBN & EAN  ; 
 aac <=  iee  |  ied  |  IEC  ; 
 aad <=  iee  |  ied  |  iec  ; 
 aaa <=  iee  |  IED  |  IEC  ; 
 aab <=  iee  |  IED  |  iec  ; 
 LAA <=  LAA & TAI & tab  |  IFA & tai  |  JAA & TAB  ; 
 LBA <=  LAA & TAI & tab  |  IFA & tai  |  JAA & TAB  ; 
 OQA <=  TAC & JAG & jah  |  QIA  |  JAH & QNB  ; 
 QAI <=  TAC & JAG & jah  |  QIA  |  JAH & QNB  ; 
 LAB <=  LAB & TAI & tab  |  IFB & tai  |  JAB & TAB  ; 
 LBB <=  LAB & TAI & tab  |  IFB & tai  |  JAB & TAB  ; 
 OAI <= EAR ; 
 OAJ <= EAR ; 
 OAK <= EAR ; 
 OAL <= EAR ; 
 LAC <=  LAC & TAI & tab  |  IFC & tai  |  JAC & TAB  ; 
 LBC <=  LAC & TAI & tab  |  IFC & tai  |  JAC & TAB  ; 
 OAE <= EAQ ; 
 OAF <= EAQ ; 
 OAG <= EAQ ; 
 OAH <= EAQ ; 
 OAM <= EAR ; 
 OAN <= EAR ; 
 OAO <= EAR ; 
 OAP <= EAR ; 
 hai <=  hai & gai  |  HAI & GAI  |  TAO  ; 
 hbi <=  hai & gai  |  HAI & GAI  |  TAO  ; 
 haj <=  haj & gaj  |  HAJ & GAJ  |  TAO  ; 
 hbj <=  haj & gaj  |  HAJ & GAJ  |  TAO  ; 
 hak <=  hak & gak  |  HAK & GAK  |  TAO  ; 
 hbk <=  hak & gak  |  HAK & GAK  |  TAO  ; 
 hal <=  hal & gal  |  HAL & GAL  |  TAO  ; 
 hbl <=  hal & gal  |  HAL & GAL  |  TAO  ; 
 qag <=  tae  |  pac  ; 
 qah <=  tae  |  pad  ; 
 ham <=  ham & gam  |  HAM & GAM  |  TAP  ; 
 hbm <=  ham & gam  |  HAM & GAM  |  TAP  ; 
 han <=  han & gan  |  HAN & GAN  |  TAP  ; 
 hbn <=  han & gan  |  HAN & GAN  |  TAP  ; 
 OFC <=  HDA & ECA  |  HDE & ECE  |  HDI & ECI  |  HDM & ECM  ; 
 hao <=  hao & gao  |  HAO & GAO  |  TAP  ; 
 hbo <=  hao & gao  |  HAO & GAO  |  TAP  ; 
 hap <=  hap & gap  |  HAP & GAP  |  TAP  ; 
 hbp <=  hap & gap  |  HAP & GAP  |  TAP  ; 
 QAP <=  QAJ  |  QNA  ; 
 OEM <= ECR ; 
 OEO <= ECR ; 
 OCA <=  HBC & EAC  |  HBG & EAG  |  HBK & EAK  |  HBO & EAO  ; 
 OCB <=  HBC & EAC  |  HBG & EAG  |  HBK & EAK  |  HBO & EAO  ; 
 OCI <=  HBD & EAD  |  HBH & EAH  |  HBL & EAL  |  HBP & EAP  ; 
 OCJ <=  HBD & EAD  |  HBH & EAH  |  HBL & EAL  |  HBP & EAP  ; 
 OCC <=  HBC & EAC  |  HBG & EAG  |  HBK & EAK  |  HBO & EAO  ; 
 OCD <=  HBC & EAC  |  HBG & EAG  |  HBK & EAK  |  HBO & EAO  ; 
 OCK <=  HBD & EAD  |  HBH & EAH  |  HBL & EAL  |  HBP & EAP  ; 
 OCL <=  HBD & EAD  |  HBH & EAH  |  HBL & EAL  |  HBP & EAP  ; 
 ODA <= QAK ; 
 ODB <= QAK ; 
 ODC <= QAK ; 
 ODD <= QAK ; 
 OCE <=  HBC & EAC  |  HBG & EAG  |  HBK & EAK  |  HBO & EAO  ; 
 OCF <=  HBC & EAC  |  HBG & EAG  |  HBK & EAK  |  HBO & EAO  ; 
 OCM <=  HBD & EAD  |  HBH & EAH  |  HBL & EAL  |  HBP & EAP  ; 
 OCN <=  HBD & EAD  |  HBH & EAH  |  HBL & EAL  |  HBP & EAP  ; 
 QAJ <=  QAJ & qai  |  QAN & QKB  ; 
 QAL <=  QAL & jag & jah  |  JAH & qnb  |  IDA  ; 
 OCG <=  HBC & EAC  |  HBG & EAG  |  HBK & EAK  |  HBO & EAO  ; 
 OCH <=  HBC & EAC  |  HBG & EAG  |  HBK & EAK  |  HBO & EAO  ; 
 OCO <=  HBD & EAD  |  HBH & EAH  |  HBL & EAL  |  HBP & EAP  ; 
 OCP <=  HBD & EAD  |  HBH & EAH  |  HBL & EAL  |  HBP & EAP  ; 
 QAB <=  QAA & qla  |  QAA & jag  |  QAB & qac  |  QAB & jag  ; 
 QBB <=  QAA & qla  |  QAA & jag  |  QAB & qac  |  QAB & jag  ; 
 qaa <=  iaa  |  iab  |  iba  ; 
 qba <=  iaa  |  iab  |  iba  ; 
 qan <= iba ; 
 QAC <=  ica & icb  |  QAA & QJA  |  QAD  ; 
 LAD <=  LAD & TAJ & tad  |  IFD & taj  |  JAD & TAD  ; 
 LBD <=  LAD & TAJ & tad  |  IFD & taj  |  JAD & TAD  ; 
 QAD <=  QAA & QJA  |  QAB & QAD  ; 
 QAK <=  QKA & IBA  |  QAK & qai  ; 
 LAE <=  LAE & TAJ & tad  |  IFE & taj  |  JAE & TAD  ; 
 LBE <=  LAE & TAJ & tad  |  IFE & taj  |  JAE & TAD  ; 
 ODI <= TAE ; 
 ODJ <= TAE ; 
 ODK <= TAE ; 
 ODL <= TAE ; 
 LAF <=  LAF & TAJ & tad  |  IFFF  & taj  |  JAF & TAD  ; 
 ODE <= QAK ; 
 ODF <= QAK ; 
 ODG <= QAK ; 
 ODH <= QAK ; 
 ODM <= TAE ; 
 ODN <= TAE ; 
 ODO <= TAE ; 
 ODP <= TAE ; 
 hca <=  hca & gca  |  HCA & GCA  |  TCM  ; 
 hda <=  hca & gca  |  HCA & GCA  |  TCM  ; 
 hcb <=  hcb & gcb  |  HCB & GCB  |  TCM  ; 
 hdb <=  hcb & gcb  |  HCB & GCB  |  TCM  ; 
 hcc <=  hcc & gcc  |  HCC & GCC  |  TCM  ; 
 hdc <=  hcc & gcc  |  HCC & GCC  |  TCM  ; 
 hcd <=  hcd & gcd  |  HCD & GCD  |  TCM  ; 
 hdd <=  hcd & gcd  |  HCD & GCD  |  TCM  ; 
 qce <=  tcc  |  pca  ; 
 qcf <=  tcc  |  pcb  ; 
 hce <=  hce & gce  |  HCE & GCE  |  TCN  ; 
 hde <=  hce & gce  |  HCE & GCE  |  TCN  ; 
 hdg <=  hcg & gcg  |  HCG & GCG  |  TCN  ; 
 PCA <=  JDA & tck & tca  |  ABA & TCK  |  JDE & TCA  ; 
 PDA <=  JDA & tck & tca  |  ABA & TCK  |  JDE & TCA  ; 
 hcf <=  hcf & gcf  |  HCF & GCF  |  TCN  ; 
 hdf <=  hcf & gcf  |  HCF & GCF  |  TCN  ; 
 hhm <=  hgm & ggm  |  HGM & GGM  |  TGP  ; 
 PCB <=  JDB & tck & tca  |  ABB & TCK  |  JDF & TCA  ; 
 PDB <=  JDB & tck & tca  |  ABB & TCK  |  JDF & TCA  ; 
 hcg <=  hcg & gcg  |  HCG & GCG  |  TCN  ; 
 PCC <=  JDC & tck & tca  |  ABC & TCK  |  JDG & TCA  ; 
 PDC <=  JDC & tck & tca  |  ABC & TCK  |  JDG & TCA  ; 
 hch <=  hch & gch  |  HCH & GCH  |  TCN  ; 
 hdh <=  hch & gch  |  HCH & GCH  |  TCN  ; 
 PCD <=  JDD & tck & tca  |  ABD & TCK  |  JDH & TCA  ; 
 PDD <=  JDD & tck & tca  |  ABD & TCK  |  JDH & TCA  ; 
 KCC <= LDB ; 
 KCD <=  LDB  |  LDC  ; 
 KCE <=  LDB  |  LDC  |  LDD  ; 
 KCF <=  LDB  |  LDC  |  LDD  |  LDE  ; 
 OFA <=  HDA & ECA  |  HDE & ECE  |  HDI & ECI  |  HDM & ECM  ; 
 OFB <=  HDA & ECA  |  HDE & ECE  |  HDI & ECI  |  HDM & ECM  ; 
 OFI <=  HDB & ECB  |  HDF & ECF  |  HDJ & ECJ  |  HDN & ECN  ; 
 OFJ <=  HDB & ECB  |  HDF & ECF  |  HDJ & ECJ  |  HDN & ECN  ; 
 OFD <=  HDA & ECA  |  HDE & ECE  |  HDI & ECI  |  HDM & ECM  ; 
 OFK <=  HDB & ECB  |  HDF & ECF  |  HDJ & ECJ  |  HDN & ECN  ; 
 OFL <=  HDB & ECB  |  HDF & ECF  |  HDJ & ECJ  |  HDN & ECN  ; 
 OEA <= ECQ ; 
 OEB <= ECQ ; 
 OEC <= ECQ ; 
 OED <= ECQ ; 
 OFE <=  HDA & ECA  |  HDE & ECE  |  HDI & ECI  |  HDM & ECM  ; 
 OFF <=  HDA & ECA  |  HDE & ECE  |  HDI & ECI  |  HDM & ECM  ; 
 OFM <=  HDB & ECB  |  HDF & ECF  |  HDJ & ECJ  |  HDN & ECN  ; 
 OFN <=  HDB & ECB  |  HDF & ECF  |  HDJ & ECJ  |  HDN & ECN  ; 
 QCM <= AAB ; 
 OFG <=  HDA & ECA  |  HDE & ECE  |  HDI & ECI  |  HDM & ECM  ; 
 OFH <=  HDA & ECA  |  HDE & ECE  |  HDI & ECI  |  HDM & ECM  ; 
 OFO <=  HDB & ECB  |  HDF & ECF  |  HDJ & ECJ  |  HDN & ECN  ; 
 OFP <=  HDB & ECB  |  HDF & ECF  |  HDJ & ECJ  |  HDN & ECN  ; 
 qla <=  ICA & ibe  |  ICB & ibe  ; 
 qlb <=  ICA & ibe  |  ICB & ibe  ; 
 qja <=  ibe  ; 
 qkb <=  qka  |  ibe  ; 
 LCA <=  LCA & TCI & tcb  |  IFA & tci  |  JCA & TCB  ; 
 LDA <=  LCA & TCI & tcb  |  IFA & tci  |  JCA & TCB  ; 
 OQB <=  TCC & JCG & JCH  |  QIA  |  JCH & QNB  ; 
 QCI <=  TCC & JCG & JCH  |  QIA  |  JCH & QNB  ; 
 LCB <=  LCB & TCI & tcb  |  IFB & tci  |  JCB & TCB  ; 
 LDB <=  LCB & TCI & tcb  |  IFB & tci  |  JCB & TCB  ; 
 OEI <= ECR ; 
 OEJ <= ECR ; 
 OEK <= ECR ; 
 OEL <= ECR ; 
 LCC <=  LCC & TCI & tcb  |  IFC & tci  |  JCC & TCB  ; 
 LDC <=  LCC & TCI & tcb  |  IFC & tci  |  JCC & TCB  ; 
 OEE <= ECQ ; 
 OEF <= ECQ ; 
 OEG <= ECQ ; 
 OEH <= ECQ ; 
 OEN <= ECR ; 
 OEP <= ECR ; 
 hci <=  hci & gci  |  HCI & GCI  |  TCO  ; 
 hdi <=  hci & gci  |  HCI & GCI  |  TCO  ; 
 hcj <=  hcj & gcj  |  HCJ & GCJ  |  TCO  ; 
 hdj <=  hcj & gcj  |  HCJ & GCJ  |  TCO  ; 
 hck <=  hck & gck  |  HCK & GCK  |  TCO  ; 
 hdk <=  hck & gck  |  HCK & GCK  |  TCO  ; 
 hcl <=  hcl & gcl  |  HCL & GCL  |  TCO  ; 
 hdl <=  hcl & gcl  |  HCL & GCL  |  TCO  ; 
 qcg <=  tce  |  pcc  ; 
 qch <=  tce  |  pcd  ; 
 hcm <=  hcm & gcm  |  HCM & GCM  |  TCP  ; 
 hdm <=  hcm & gcm  |  HCM & GCM  |  TCP  ; 
 hcn <=  hcn & gcn  |  HCN & GCN  |  TCP  ; 
 hdn <=  hcn & gcn  |  HCN & GCN  |  TCP  ; 
 hco <=  hco & gco  |  HCO & GCO  |  TCP  ; 
 hdo <=  hco & gco  |  HCO & GCO  |  TCP  ; 
 hcp <=  hcp & gcp  |  HCP & GCP  |  TCP  ; 
 hdp <=  hcp & gcp  |  HCP & GCP  |  TCP  ; 
 QCP <=  QCJ  |  QNA  ; 
 OGA <=  HDC & ECC  |  HDG & ECG  |  HDK & ECK  |  HDO & ECO  ; 
 OGB <=  HDC & ECC  |  HDG & ECG  |  HDK & ECK  |  HDO & ECO  ; 
 OGI <=  HDD & ECD  |  HDH & ECH  |  HDL & ECL  |  HDP & ECP  ; 
 OGJ <=  HDD & ECD  |  HDH & ECH  |  HDL & ECL  |  HDP & ECP  ; 
 QCK <=  QKA & IBB  |  QCK & gci  ; 
 OGC <=  HDC & ECC  |  HDG & ECG  |  HDK & ECK  |  HDO & ECO  ; 
 OGD <=  HDC & ECC  |  HDG & ECG  |  HDK & ECK  |  HDO & ECO  ; 
 OGK <=  HDD & ECD  |  HDH & ECH  |  HDL & ECL  |  HDP & ECP  ; 
 OGL <=  HDD & ECD  |  HDH & ECH  |  HDL & ECL  |  HDP & ECP  ; 
 OHA <= QCK ; 
 OHB <= QCK ; 
 OHC <= QCK ; 
 OHD <= QCK ; 
 OGE <=  HDC & ECC  |  HDG & ECG  |  HDK & ECK  |  HDO & ECO  ; 
 OGF <=  HDC & ECC  |  HDG & ECG  |  HDK & ECK  |  HDO & ECO  ; 
 OGM <=  HDD & ECD  |  HDH & ECH  |  HDL & ECL  |  HDP & ECP  ; 
 OGN <=  HDD & ECD  |  HDH & ECH  |  HDL & ECL  |  HDP & ECP  ; 
 QCJ <=  QCJ & gci  |  QCN & QKB  ; 
 QCL <=  QCL & jcg & jch  |  JCH & qnb  |  IDB  ; 
 OGG <=  HDC & ECC  |  HDG & ECG  |  HDK & ECK  |  HDO & ECO  ; 
 OGH <=  HDC & ECC  |  HDG & ECG  |  HDK & ECK  |  HDO & ECO  ; 
 OGO <=  HDD & ECD  |  HDH & ECH  |  HDL & ECL  |  HDP & ECP  ; 
 OGP <=  HDD & ECD  |  HDH & ECH  |  HDL & ECL  |  HDP & ECP  ; 
 QCB <=  QCA & qla  |  QCA & jcg  |  QCB & qcc  |  QCB & jcg  ; 
 QDB <=  QCA & qla  |  QCA & jcg  |  QCB & qcc  |  QCB & jcg  ; 
 qca <=  iaa  |  iab  |  ibb  ; 
 qda <=  iaa  |  iab  |  ibb  ; 
 qcn <= ibb ; 
 QCC <=  ica & icb  |  QCA & QJA  |  QCD  ; 
 LCD <=  LCD & TCJ & tcd  |  IFD & tcj  |  JCD & TCD  ; 
 LDD <=  LCD & TCJ & tcd  |  IFD & tcj  |  JCD & TCD  ; 
 QCD <=  QCA & QJA  |  QCB & QCD  ; 
 LCE <=  LCE & TCJ & tcd  |  IFE & tcj  |  JCE & TCD  ; 
 LDE <=  LCE & TCJ & tcd  |  IFE & tcj  |  JCE & TCD  ; 
 OHI <= TCE ; 
 OHJ <= TCE ; 
 OHK <= TCE ; 
 OHL <= TCE ; 
 LCF <=  LCF & TCJ & tcd  |  IFFF  & tcj  |  JCF & TCD  ; 
 OHE <= QCK ; 
 OHF <= QCK ; 
 OHG <= QCK ; 
 OHH <= QCK ; 
 OHM <= TCE ; 
 OHN <= TCE ; 
 OHO <= TCE ; 
 OHP <= TCE ; 
 hea <=  hea & gea  |  HEA & GEA  |  TEM  ; 
 hfa <=  hea & gea  |  HEA & GEA  |  TEM  ; 
 heb <=  heb & geb  |  HEB & GEB  |  TEM  ; 
 hfb <=  heb & geb  |  HEB & GEB  |  TEM  ; 
 hho <=  hgo & ggo  |  HGO & GGO  |  TGP  ; 
 hec <=  hec & gec  |  HEC & GEC  |  TEM  ; 
 hfc <=  hec & gec  |  HEC & GEC  |  TEM  ; 
 hed <=  hed & ged  |  HED & GED  |  TEM  ; 
 hfd <=  hed & ged  |  HED & GED  |  TEM  ; 
 qee <=  tec  |  pea  ; 
 qef <=  tec  |  peb  ; 
 hee <=  hee & gee  |  HEE & GEE  |  TEN  ; 
 hfe <=  hee & gee  |  HEE & GEE  |  TEN  ; 
 PEA <=  JFA & tek & tea  |  ABA & TEK  |  JFE & TEA  ; 
 PFA <=  JFA & tek & tea  |  ABA & TEK  |  JFE & TEA  ; 
 hef <=  hef & gef  |  HEF & GEF  |  TEN  ; 
 hff <=  hef & gef  |  HEF & GEF  |  TEN  ; 
 PEB <=  JFB & tek & tea  |  ABB & TEK  |  JFF & TEA  ; 
 PFB <=  JFB & tek & tea  |  ABB & TEK  |  JFF & TEA  ; 
 heg <=  heg & geg  |  HEG & GEG  |  TEN  ; 
 hfg <=  heg & geg  |  HEG & GEG  |  TEN  ; 
 PEC <=  JFC & tek & tea  |  ABC & TEK  |  JFG & TEA  ; 
 PFC <=  JFC & tek & tea  |  ABC & TEK  |  JFG & TEA  ; 
 heh <=  heh & geh  |  HEH & GEH  |  TEN  ; 
 hfh <=  heh & geh  |  HEH & GEH  |  TEN  ; 
 PED <=  JFD & tek & tea  |  ABD & TEK  |  JFH & TEA  ; 
 PFD <=  JFD & tek & tea  |  ABD & TEK  |  JFH & TEA  ; 
 KEC <= LFB ; 
 KED <=  LFB  |  LFC  ; 
 KEE <=  LFB  |  LFC  |  LFD  ; 
 KEF <=  LFB  |  LFC  |  LFD  |  LFE  ; 
 OJA <=  HFA & EEA  |  HFE & EEE  |  HFI & EEI  |  HFM & EEM  ; 
 OJB <=  HFA & EEA  |  HFE & EEE  |  HFI & EEI  |  HFM & EEM  ; 
 OJI <=  HFB & EEB  |  HFF & EEF  |  HFJ & EEJ  |  HFN & EEN  ; 
 OJJ <=  HFB & EEB  |  HFF & EEF  |  HFJ & EEJ  |  HFN & EEN  ; 
 OJC <=  HFA & EEA  |  HFE & EEE  |  HFI & EEI  |  HFM & EEM  ; 
 OJD <=  HFA & EEA  |  HFE & EEE  |  HFI & EEI  |  HFM & EEM  ; 
 OJK <=  HFB & EEB  |  HFF & EEF  |  HFJ & EEJ  |  HFN & EEN  ; 
 OJL <=  HFB & EEB  |  HFF & EEF  |  HFJ & EEJ  |  HFN & EEN  ; 
 OIA <= EEQ ; 
 OIB <= EEQ ; 
 OIC <= EEQ ; 
 OID <= EEQ ; 
 OJF <=  HFA & EEA  |  HFE & EEE  |  HFI & EEI  |  HFM & EEM  ; 
 OJE <=  HFA & EEA  |  HFE & EEE  |  HFI & EEI  |  HFM & EEM  ; 
 OJM <=  HFB & EEB  |  HFF & EEF  |  HFJ & EEJ  |  HFN & EEN  ; 
 OJN <=  HFB & EEB  |  HFF & EEF  |  HFJ & EEJ  |  HFN & EEN  ; 
 QEM <= AAC ; 
 OJG <=  HFA & EEA  |  HFE & EEE  |  HFI & EEI  |  HFM & EEM  ; 
 OJH <=  HFA & EEA  |  HFE & EEE  |  HFI & EEI  |  HFM & EEM  ; 
 OJO <=  HFB & EEB  |  HFF & EEF  |  HFJ & EEJ  |  HFN & EEN  ; 
 OJP <=  HFB & EEB  |  HFF & EEF  |  HFJ & EEJ  |  HFN & EEN  ; 
 aba <=  IEB  |  IEA  ; 
 abb <=  IEB  |  iea  ; 
 abc <=  ieb  |  EEA  ; 
 abd <=  ieb  |  iea  ; 
 LEA <=  LEA & TEI & teb  |  IFA & tei  |  JEA & TEB  ; 
 LFA <=  LEA & TEI & teb  |  IFA & tei  |  JEA & TEB  ; 
 OQC <=  TEC & JEG & jeh  |  QIA  |  JEH & QNB  ; 
 QEI <=  TEC & JEG & jeh  |  QIA  |  JEH & QNB  ; 
 LEB <=  LEB & TEI & teb  |  IFB & tei  |  JEB & TEB  ; 
 LFB <=  LEB & TEI & teb  |  IFB & tei  |  JEB & TEB  ; 
 OII <= EER ; 
 OIJ <= EER ; 
 OIK <= EER ; 
 OIL <= EER ; 
 LEC <=  LEC & TEI & teb  |  IFC & tei  |  JEC & TEB  ; 
 LFC <=  LEC & TEI & teb  |  IFC & tei  |  JEC & TEB  ; 
 OIE <= EEQ ; 
 OIF <= EEQ ; 
 OIG <= EEQ ; 
 OIH <= EEQ ; 
 OIM <= EER ; 
 OIN <= EER ; 
 OIO <= EER ; 
 OIP <= EER ; 
 hei <=  hei & gei  |  HEI & GEI  |  TEO  ; 
 hfi <=  hei & gei  |  HEI & GEI  |  TEO  ; 
 hej <=  hej & gej  |  HEJ & GEJ  |  TEO  ; 
 hfj <=  hej & gej  |  HEJ & GEJ  |  TEO  ; 
 hek <=  hek & gek  |  HEK & GEK  |  TEO  ; 
 hfk <=  hek & gek  |  HEK & GEK  |  TEO  ; 
 hel <=  hel & gel  |  HEL & GEL  |  TEO  ; 
 hfl <=  hel & gel  |  HEL & GEL  |  TEO  ; 
 qeg <=  tee  |  pec  ; 
 qeh <=  tee  |  ped  ; 
 hem <=  hem & gem  |  HEM & GEM  |  TEP  ; 
 hfm <=  hem & gem  |  HEM & GEM  |  TEP  ; 
 hen <=  hen & gen  |  HEN & GEN  |  TEP  ; 
 hfn <=  hen & gen  |  HEN & GEN  |  TEP  ; 
 heo <=  heo & geo  |  HEO & GEO  |  TEP  ; 
 hfo <=  heo & geo  |  HEO & GEO  |  TEP  ; 
 hep <=  hep & gep  |  HEP & GEP  |  TEP  ; 
 hfp <=  hep & gep  |  HEP & GEP  |  TEP  ; 
 QEP <=  QEJ  |  QNA  ; 
 OKA <=  HFC & EEC  |  HFG & EEG  |  HFK & EEK  |  HFO & EEO  ; 
 OKB <=  HFC & EEC  |  HFG & EEG  |  HFK & EEK  |  HFO & EEO  ; 
 OKI <=  HFD & EED  |  HFH & EEH  |  HFL & EEL  |  HFP & EEP  ; 
 OKJ <=  HFD & EED  |  HFH & EEH  |  HFL & EEL  |  HFP & EEP  ; 
 OKC <=  HFC & EEC  |  HFG & EEG  |  HFK & EEK  |  HFO & EEO  ; 
 OKD <=  HFC & EEC  |  HFG & EEG  |  HFK & EEK  |  HFO & EEO  ; 
 OKK <=  HFD & EED  |  HFH & EEH  |  HFL & EEL  |  HFP & EEP  ; 
 OKL <=  HFD & EED  |  HFH & EEH  |  HFL & EEL  |  HFP & EEP  ; 
 OKE <=  HFC & EEC  |  HFG & EEG  |  HFK & EEK  |  HFO & EEO  ; 
 OKF <=  HFC & EEC  |  HFG & EEG  |  HFK & EEK  |  HFO & EEO  ; 
 OKM <=  HFD & EED  |  HFH & EEH  |  HFL & EEL  |  HFP & EEP  ; 
 OKN <=  HFD & EED  |  HFH & EEH  |  HFL & EEL  |  HFP & EEP  ; 
 QEJ <=  QEJ & qei  |  QEN & QKB  ; 
 QEK <=  QEK & qei  |  ZZI & QKB  |  QKA & IBC  ; 
 QEL <=  QEL & jeg & jeh  |  JEH & qnb  |  IDC  ; 
 OKG <=  HFC & EEC  |  HFG & EEG  |  HFK & EEK  |  HFO & EEO  ; 
 OKH <=  HFC & EEC  |  HFG & EEG  |  HFK & EEK  |  HFO & EEO  ; 
 OKO <=  HFD & EED  |  HFH & EEH  |  HFL & EEL  |  HFP & EEP  ; 
 OKP <=  HFD & EED  |  HFH & EEH  |  HFL & EEL  |  HFP & EEP  ; 
 QEB <=  QEA & qla  |  QEA & jeg  |  QEB & qec  |  QEB & jeg  ; 
 QFB <=  QEA & qla  |  QEA & jeg  |  QEB & qec  |  QEB & jeg  ; 
 qea <=  iaa  |  iab  |  ibc  ; 
 qfa <=  iaa  |  iab  |  ibc  ; 
 qen <= ibc ; 
 QNA <= IHA ; 
 QEC <=  ica & icb  |  QEA & QJA  |  QED  ; 
 LED <=  LED & TEJ & ted  |  IFD & tej  |  JED & TED  ; 
 LFD <=  LED & TEJ & ted  |  IFD & tej  |  JED & TED  ; 
 QED <=  QEA & QJA  |  QEB & QED  ; 
 LEE <=  LEE & TEJ & ted  |  IFE & tej  |  JEE & TED  ; 
 LFE <=  LEE & TEJ & ted  |  IFE & tej  |  JEE & TED  ; 
 OLA <= QEK ; 
 OLB <= QEK ; 
 OLC <= QEK ; 
 OLD <= QEK ; 
 OLI <= TEE ; 
 OLJ <= TEE ; 
 OLK <= TEE ; 
 OLL <= TEE ; 
 LEF <=  LEF & TEJ & ted  |  IFFF  & tej  |  JEF & TED  ; 
 OLE <= QEK ; 
 OLF <= QEK ; 
 OLG <= QEK ; 
 OLH <= QEK ; 
 OLM <= TEE ; 
 OLN <= TEE ; 
 OLO <= TEE ; 
 OLP <= TEE ; 
 hga <=  hga & gga  |  HGA & GGA  |  TGM  ; 
 hha <=  hga & gga  |  HGA & GGA  |  TGM  ; 
 hgb <=  hgb & ggb  |  HGB & GGB  |  TGM  ; 
 hhb <=  hgb & ggb  |  HGB & GGB  |  TGM  ; 
 hgc <=  hgc & ggc  |  HGC & GGC  |  TGM  ; 
 hhc <=  hgc & ggc  |  HGC & GGC  |  TGM  ; 
 hgd <=  hgd & ggd  |  HGD & GGD  |  TGM  ; 
 hhd <=  hgd & ggd  |  HGD & GGD  |  TGM  ; 
 qge <=  tgc  |  pga  ; 
 qgf <=  tgc  |  pgb  ; 
 hge <=  hge & gge  |  HGE & GGE  |  TGN  ; 
 hhe <=  hge & gge  |  HGE & GGE  |  TGN  ; 
 PGA <=  JHA & tgk & tga  |  ABA & TGK  |  JHE & TGA  ; 
 PHA <=  JHA & tgk & tga  |  ABA & TGK  |  JHE & TGA  ; 
 hgf <=  hgf & ggf  |  HGF & GGF  |  TGN  ; 
 hhf <=  hgf & ggf  |  HGF & GGF  |  TGN  ; 
 PGB <=  JHB & tgk & tga  |  ABB & TGK  |  JHF & TGA  ; 
 PHB <=  JHB & tgk & tga  |  ABB & TGK  |  JHF & TGA  ; 
 hgg <=  hgg & ggg  |  HGG & GGG  |  TGN  ; 
 hhg <=  hgg & ggg  |  HGG & GGG  |  TGN  ; 
 PGC <=  JHC & tgk & tga  |  ABC & TGK  |  JHG & TGA  ; 
 PHC <=  JHC & tgk & tga  |  ABC & TGK  |  JHG & TGA  ; 
 hgh <=  hgh & ggh  |  HGH & GGH  |  TGN  ; 
 hhh <=  hgh & ggh  |  HGH & GGH  |  TGN  ; 
 PGD <=  JHD & tgk & tga  |  ABD & TGK  |  JHH & TGA  ; 
 PHD <=  JHD & tgk & tga  |  ABD & TGK  |  JHH & TGA  ; 
 KGC <= LHB ; 
 KGE <=  LHB  |  LHC  |  LHD  ; 
 KGD <=  LHB  |  LHC  ; 
 KGF <=  LHB  |  LHC  |  LHD  |  LHE  ; 
 ONA <=  HHA & EGA  |  HHE & EGE  |  HHI & EGI  |  HHM & EGM  ; 
 ONB <=  HHA & EGA  |  HHE & EGE  |  HHI & EGI  |  HHM & EGM  ; 
 ONI <=  HHB & EGB  |  HHF & EGF  |  HHJ & EGJ  |  HHN & EGN  ; 
 ONJ <=  HHB & EGB  |  HHF & EGF  |  HHJ & EGJ  |  HHN & EGN  ; 
 ONC <=  HHA & EGA  |  HHE & EGE  |  HHI & EGI  |  HHM & EGM  ; 
 OND <=  HHA & EGA  |  HHE & EGE  |  HHI & EGI  |  HHM & EGM  ; 
 ONK <=  HHB & EGB  |  HHF & EGF  |  HHJ & EGJ  |  HHN & EGN  ; 
 ONL <=  HHB & EGB  |  HHF & EGF  |  HHJ & EGJ  |  HHN & EGN  ; 
 ONE <=  HHA & EGA  |  HHE & EGE  |  HHI & EGI  |  HHM & EGM  ; 
 ONF <=  HHA & EGA  |  HHE & EGE  |  HHI & EGI  |  HHM & EGM  ; 
 ONM <=  HHB & EGB  |  HHF & EGF  |  HHJ & EGJ  |  HHN & EGN  ; 
 ONN <=  HHB & EGB  |  HHF & EGF  |  HHJ & EGJ  |  HHN & EGN  ; 
 QGM <= AAD ; 
 ONG <=  HHA & EGA  |  HHE & EGE  |  HHI & EGI  |  HHM & EGM  ; 
 ONH <=  HHA & EGA  |  HHE & EGE  |  HHI & EGI  |  HHM & EGM  ; 
 ONO <=  HHB & EGB  |  HHF & EGF  |  HHJ & EGJ  |  HHN & EGN  ; 
 ONP <=  HHB & EGB  |  HHF & EGF  |  HHJ & EGJ  |  HHN & EGN  ; 
 QKA <=  IAA & IAB  ; 
 LGA <=  LGA & TGI & tgb  |  IFA & tgi  |  JGA & TGB  ; 
 LHA <=  LGA & TGI & tgb  |  IFA & tgi  |  JGA & TGB  ; 
 QIA <= IGA ; 
 OQD <=  TGC & JGG & jgh  |  QIA  |  JGH & QNB  ; 
 QGI <=  TGC & JGG & jgh  |  QIA  |  JGH & QNB  ; 
 LGB <=  LGB & TGI & tgb  |  IFB & tgi  |  JGB & TGB  ; 
 LHB <=  LGB & TGI & tgb  |  IFB & tgi  |  JGB & TGB  ; 
 OMA <= EGQ ; 
 OMB <= EGQ ; 
 OMC <= EGQ ; 
 OMD <= EGQ ; 
 OMI <= EGR ; 
 OMJ <= EGR ; 
 OMK <= EGR ; 
 OML <= EGR ; 
 LGC <=  LGC & TGI & tgb  |  IFC & tgi  |  JGC & TGB  ; 
 LHC <=  LGC & TGI & tgb  |  IFC & tgi  |  JGC & TGB  ; 
 OME <= EGQ ; 
 OMF <= EGQ ; 
 OMG <= EGQ ; 
 OMH <= EGQ ; 
 OMM <= EGR ; 
 OMN <= EGR ; 
 OMO <= EGR ; 
 OMP <= EGR ; 
 hgi <=  hgi & ggi  |  HGI & GGI  |  TGO  ; 
 hhi <=  hgi & ggi  |  HGI & GGI  |  TGO  ; 
 hhn <=  hgn & ggn  |  HGN & GGN  |  TGP  ; 
 hgj <=  hgj & ggj  |  HGJ & GGJ  |  TGO  ; 
 hhj <=  hgj & ggj  |  HGJ & GGJ  |  TGO  ; 
 hgk <=  hgk & ggk  |  HGK & GGK  |  TGO  ; 
 hhk <=  hgk & ggk  |  HGK & GGK  |  TGO  ; 
 hgl <=  hgl & ggl  |  HGL & GGL  |  TGO  ; 
 hhl <=  hgl & ggl  |  HGL & GGL  |  TGO  ; 
 qgg <=  tge  |  pgc  ; 
 qgh <=  tge  |  pgd  ; 
 hgm <=  hgm & ggm  |  HGM & GGM  |  TGP  ; 
 hgn <=  hgn & ggn  |  HGN & GGN  |  TGP  ; 
 hgo <=  hgo & ggo  |  HGO & GGO  |  TGP  ; 
 hgp <=  hgp & ggp  |  HGP & GGP  |  TGP  ; 
 hhp <=  hgp & ggp  |  HGP & GGP  |  TGP  ; 
 QGP <=  QGJ  |  QNA  ; 
 OOA <=  HHC & EGC  |  HHG & EGG  |  HHK & EGK  |  HHO & EGO  ; 
 OOB <=  HHC & EGC  |  HHG & EGG  |  HHK & EGK  |  HHO & EGO  ; 
 OOI <=  HHD & EGD  |  HHH & EGH  |  HHL & EGL  |  HHP & EGP  ; 
 OOJ <=  HHD & EGD  |  HHH & EGH  |  HHL & EGL  |  HHP & EGP  ; 
 QGK <=  QKA & IBD  |  QGK & qgi  ; 
 OOC <=  HHC & EGC  |  HHG & EGG  |  HHK & EGK  |  HHO & EGO  ; 
 OOD <=  HHC & EGC  |  HHG & EGG  |  HHK & EGK  |  HHO & EGO  ; 
 OOK <=  HHD & EGD  |  HHH & EGH  |  HHL & EGL  |  HHP & EGP  ; 
 OOL <=  HHD & EGD  |  HHH & EGH  |  HHL & EGL  |  HHP & EGP  ; 
 OPA <= QGK ; 
 OPB <= QGK ; 
 OPC <= QGK ; 
 OPD <= QGK ; 
 OOE <=  HHC & EGC  |  HHG & EGG  |  HHK & EGK  |  HHO & EGO  ; 
 OOF <=  HHC & EGC  |  HHG & EGG  |  HHK & EGK  |  HHO & EGO  ; 
 OOM <=  HHD & EGD  |  HHH & EGH  |  HHL & EGL  |  HHP & EGP  ; 
 OON <=  HHD & EGD  |  HHH & EGH  |  HHL & EGL  |  HHP & EGP  ; 
 QGJ <=  QGJ & qgi  |  QGN & QKB  ; 
 QGL <=  QGL & jgg & jgh  |  JGH & qnb  |  IDD  ; 
 OOG <=  HHC & EGC  |  HHG & EGG  |  HHK & EGK  |  HHO & EGO  ; 
 OOH <=  HHC & EGC  |  HHG & EGG  |  HHK & EGK  |  HHO & EGO  ; 
 OOO <=  HHD & EGD  |  HHH & EGH  |  HHL & EGL  |  HHP & EGP  ; 
 OOP <=  HHD & EGD  |  HHH & EGH  |  HHL & EGL  |  HHP & EGP  ; 
 QGB <=  QGA & qla  |  QGA & jgg  |  QGB & qgc  |  QGB & jgg  ; 
 QHB <=  QGA & qla  |  QGA & jgg  |  QGB & qgc  |  QGB & jgg  ; 
 qga <=  iaa  |  iab  |  ibd  ; 
 qha <=  iaa  |  iab  |  ibd  ; 
 qgn <= ibd ; 
 QGC <=  ica & icb  |  QGA & QJA  |  QGD  ; 
 LGD <=  LGD & TGJ & tgd  |  IFD & tgj  |  JGD & TGD  ; 
 LHD <=  LGD & TGJ & tgd  |  IFD & tgj  |  JGD & TGD  ; 
 QGD <=  QGA & QJA  |  QGB & QGD  ; 
 QNB <=  IHB  |  QIA  ; 
 LGE <=  LGE & TGJ & tgd  |  IFE & tgj  |  JGE & TGD  ; 
 LHE <=  LGE & TGJ & tgd  |  IFE & tgj  |  JGE & TGD  ; 
 OPI <= TGE ; 
 OPJ <= TGE ; 
 OPK <= TGE ; 
 OPL <= TGE ; 
 LGF <=  LGF & TGJ & tgd  |  IFFF  & tgj  |  JGF & TGD  ; 
 OPE <= QGK ; 
 OPF <= QGK ; 
 OPG <= QGK ; 
 OPH <= QGK ; 
 OPM <= TGE ; 
 OPN <= TGE ; 
 OPO <= TGE ; 
 OPP <= TGE ; 
end 
endmodule;
