module ie( IZZ,
 IAA, 
 IAB, 
 IAC, 
 IAD, 
 IAE, 
 IAF, 
 IAG, 
 IAH, 
 IAI, 
 IAJ, 
 IAK, 
 IAL, 
 IAM, 
 IAN, 
 IAO, 
 IAP, 
 IBA, 
 IBB, 
 IBC, 
 IBD, 
 IBE, 
 IBF, 
 IBG, 
 IBH, 
 IBI, 
 IBJ, 
 IBK, 
 IBL, 
 IBM, 
 IBN, 
 IBO, 
 IBP, 
 ICA, 
 ICB, 
 ICC, 
 ICD, 
 ICE, 
 ICF, 
 ICG, 
 ICH, 
 ICI, 
 ICJ, 
 ICK, 
 ICL, 
 ICM, 
 ICN, 
 ICO, 
 ICP, 
 IDA, 
 IDB, 
 IDC, 
 IDD, 
 IDE, 
 IDF, 
 IDG, 
 IDH, 
 IDI, 
 IDJ, 
 IDK, 
 IDL, 
 IDM, 
 IDN, 
 IDO, 
 IDP, 
 IEA, 
 IEB, 
 IEC, 
 IED, 
 IEE, 
 IEF, 
 IEG, 
 IEH, 
 IEI, 
 IEJ, 
 IFA, 
 IFB, 
 IFC, 
 IFD, 
 IFE, 
 IGA, 
 IGB, 
 IGC, 
 IHA, 
 IHB, 
 IJA, 
 IJB, 
 IJD, 
 IJE, 
 IJF, 
 IJG, 
 OAA, 
 OAB, 
 OAC, 
 OAD, 
 OAE, 
 OAF, 
 OAG, 
 OAH, 
 OAI, 
 OAJ, 
 OAK, 
 OAL, 
 OAM, 
 OAN, 
 OAO, 
 OAP, 
 OBA, 
 OBB, 
 OBC, 
 OBD, 
 OBE, 
 OBF, 
 OBG, 
 OBH, 
 OBI, 
 OBJ, 
 OBK, 
 OBL, 
 OBM, 
 OBN, 
 OBO, 
 OBP, 
 OCA, 
 OCB, 
 OCC, 
 OCD, 
 OCE, 
 OCF, 
 OCG, 
 OCH, 
 OCI, 
 OCJ, 
 OCK, 
 OCL, 
 OCM, 
 OCN, 
 OCO, 
 OCP, 
 ODA, 
 ODB, 
 ODC, 
 ODD, 
 ODE, 
 ODF, 
 ODG, 
 ODH, 
 ODI, 
 ODJ, 
 ODK, 
 ODL, 
 ODM, 
 ODN, 
 ODO, 
 ODP, 
 OEA, 
 OEB, 
 OEC, 
 OED, 
 OEE, 
 OEF, 
 OEG, 
 OEH, 
 OEI, 
 OEJ, 
 OEK, 
 OEL, 
 OEM, 
 OEN, 
 OEO, 
 OEP, 
 OFA, 
 OFB, 
 OFC, 
 OFD, 
 OFE, 
 OFF, 
 OFG, 
 OFH, 
 OFI, 
 OFJ, 
 OFK, 
 OFL, 
 OFM, 
 OFN, 
 OFO, 
 OFP, 
 OGA, 
 OGB, 
 OGC, 
 OGD, 
 OGE, 
 OGF, 
 OGG, 
 OGH, 
 OGI, 
 OGJ, 
 OGK, 
 OGL, 
 OGM, 
 OGN, 
 OGO, 
 OGP, 
 OHA, 
 OHB, 
 OHC, 
 OHD, 
 OHE, 
 OHF, 
 OHG, 
 OHH, 
 OHI, 
 OHJ, 
 OHK, 
 OHL, 
 OHM, 
 OHN, 
 OHO, 
 OHP, 
 OJA, 
 OJB, 
 OJD, 
 OJF, 
 OKA, 
 OKB, 
 OKC, 
 OKG, 
 OKH, 
 OKI, 
 OKJ, 
 OKK, 
 OKL, 
 OKM, 
 OKN, 
 OKO, 
 OKP, 
 OKQ, 
 OKR, 
 OKS, 
 OKT, 
 OKU, 
 OKV, 
 OKW, 
OKX ); 
    
 input IZZ; 
 input IAA; 
 input IAB; 
 input IAC; 
 input IAD; 
 input IAE; 
 input IAF; 
 input IAG; 
 input IAH; 
 input IAI; 
 input IAJ; 
 input IAK; 
 input IAL; 
 input IAM; 
 input IAN; 
 input IAO; 
 input IAP; 
 input IBA; 
 input IBB; 
 input IBC; 
 input IBD; 
 input IBE; 
 input IBF; 
 input IBG; 
 input IBH; 
 input IBI; 
 input IBJ; 
 input IBK; 
 input IBL; 
 input IBM; 
 input IBN; 
 input IBO; 
 input IBP; 
 input ICA; 
 input ICB; 
 input ICC; 
 input ICD; 
 input ICE; 
 input ICF; 
 input ICG; 
 input ICH; 
 input ICI; 
 input ICJ; 
 input ICK; 
 input ICL; 
 input ICM; 
 input ICN; 
 input ICO; 
 input ICP; 
 input IDA; 
 input IDB; 
 input IDC; 
 input IDD; 
 input IDE; 
 input IDF; 
 input IDG; 
 input IDH; 
 input IDI; 
 input IDJ; 
 input IDK; 
 input IDL; 
 input IDM; 
 input IDN; 
 input IDO; 
 input IDP; 
 input IEA; 
 input IEB; 
 input IEC; 
 input IED; 
 input IEE; 
 input IEF; 
 input IEG; 
 input IEH; 
 input IEI; 
 input IEJ; 
 input IFA; 
 input IFB; 
 input IFC; 
 input IFD; 
 input IFE; 
 input IGA; 
 input IGB; 
 input IGC; 
 input IHA; 
 input IHB; 
 input IJA; 
 input IJB; 
 input IJD; 
 input IJE; 
 input IJF; 
 input IJG; 
 output OAA; 
 output OAB; 
 output OAC; 
 output OAD; 
 output OAE; 
 output OAF; 
 output OAG; 
 output OAH; 
 output OAI; 
 output OAJ; 
 output OAK; 
 output OAL; 
 output OAM; 
 output OAN; 
 output OAO; 
 output OAP; 
 output OBA; 
 output OBB; 
 output OBC; 
 output OBD; 
 output OBE; 
 output OBF; 
 output OBG; 
 output OBH; 
 output OBI; 
 output OBJ; 
 output OBK; 
 output OBL; 
 output OBM; 
 output OBN; 
 output OBO; 
 output OBP; 
 output OCA; 
 output OCB; 
 output OCC; 
 output OCD; 
 output OCE; 
 output OCF; 
 output OCG; 
 output OCH; 
 output OCI; 
 output OCJ; 
 output OCK; 
 output OCL; 
 output OCM; 
 output OCN; 
 output OCO; 
 output OCP; 
 output ODA; 
 output ODB; 
 output ODC; 
 output ODD; 
 output ODE; 
 output ODF; 
 output ODG; 
 output ODH; 
 output ODI; 
 output ODJ; 
 output ODK; 
 output ODL; 
 output ODM; 
 output ODN; 
 output ODO; 
 output ODP; 
 output OEA; 
 output OEB; 
 output OEC; 
 output OED; 
 output OEE; 
 output OEF; 
 output OEG; 
 output OEH; 
 output OEI; 
 output OEJ; 
 output OEK; 
 output OEL; 
 output OEM; 
 output OEN; 
 output OEO; 
 output OEP; 
 output OFA; 
 output OFB; 
 output OFC; 
 output OFD; 
 output OFE; 
 output OFF; 
 output OFG; 
 output OFH; 
 output OFI; 
 output OFJ; 
 output OFK; 
 output OFL; 
 output OFM; 
 output OFN; 
 output OFO; 
 output OFP; 
 output OGA; 
 output OGB; 
 output OGC; 
 output OGD; 
 output OGE; 
 output OGF; 
 output OGG; 
 output OGH; 
 output OGI; 
 output OGJ; 
 output OGK; 
 output OGL; 
 output OGM; 
 output OGN; 
 output OGO; 
 output OGP; 
 output OHA; 
 output OHB; 
 output OHC; 
 output OHD; 
 output OHE; 
 output OHF; 
 output OHG; 
 output OHH; 
 output OHI; 
 output OHJ; 
 output OHK; 
 output OHL; 
 output OHM; 
 output OHN; 
 output OHO; 
 output OHP; 
 output OJA; 
 output OJB; 
 output OJD; 
 output OJF; 
 output OKA; 
 output OKB; 
 output OKC; 
 output OKG; 
 output OKH; 
 output OKI; 
 output OKJ; 
 output OKK; 
 output OKL; 
 output OKM; 
 output OKN; 
 output OKO; 
 output OKP; 
 output OKQ; 
 output OKR; 
 output OKS; 
 output OKT; 
 output OKU; 
 output OKV; 
 output OKW; 
 output OKX; 
  
  
reg  DAA ;
reg  DAB ;
reg  DAC ;
reg  DAD ;
reg  DAE ;
reg  DAF ;
reg  DAG ;
reg  DAH ;
reg  DAI ;
reg  DAJ ;
reg  DAK ;
reg  DAL ;
reg  DAM ;
reg  DAN ;
reg  DAO ;
reg  DBA ;
reg  DBB ;
reg  DBC ;
reg  DBE ;
reg  DBF ;
reg  DBG ;
reg  DBI ;
reg  DBJ ;
reg  DBK ;
reg  DBM ;
reg  DBN ;
reg  DBO ;
reg  EAA ;
reg  EAB ;
reg  EAC ;
reg  EAD ;
reg  EAE ;
reg  eba ;
reg  ebb ;
reg  ebc ;
reg  ECA ;
reg  ECB ;
reg  ECC ;
reg  EDA ;
reg  EDB ;
reg  EDC ;
reg  EEA ;
reg  EEB ;
reg  EEC ;
reg  EFA ;
reg  EFB ;
reg  FAA ;
reg  FAB ;
reg  FAC ;
reg  FAD ;
reg  FAE ;
reg  FBA ;
reg  FBB ;
reg  FBC ;
reg  FBD ;
reg  FBE ;
reg  OAA ;
reg  OAB ;
reg  OAC ;
reg  OAD ;
reg  OAE ;
reg  OAF ;
reg  OAG ;
reg  OAH ;
reg  OAI ;
reg  OAJ ;
reg  OAK ;
reg  OAL ;
reg  OAM ;
reg  OAN ;
reg  OAO ;
reg  OAP ;
reg  OBA ;
reg  OBB ;
reg  OBC ;
reg  OBD ;
reg  OBE ;
reg  OBF ;
reg  OBG ;
reg  OBH ;
reg  OBI ;
reg  OBJ ;
reg  OBK ;
reg  OBL ;
reg  OBM ;
reg  OBN ;
reg  OBO ;
reg  OBP ;
reg  OCA ;
reg  OCB ;
reg  OCC ;
reg  OCD ;
reg  OCE ;
reg  OCF ;
reg  OCG ;
reg  OCH ;
reg  OCI ;
reg  OCJ ;
reg  OCK ;
reg  OCL ;
reg  OCM ;
reg  OCN ;
reg  OCO ;
reg  OCP ;
reg  ODA ;
reg  ODB ;
reg  ODC ;
reg  ODD ;
reg  ODE ;
reg  ODF ;
reg  ODG ;
reg  ODH ;
reg  ODI ;
reg  ODJ ;
reg  ODK ;
reg  ODL ;
reg  ODM ;
reg  ODN ;
reg  ODO ;
reg  ODP ;
reg  oea ;
reg  oeb ;
reg  oec ;
reg  oed ;
reg  oee ;
reg  oef ;
reg  oeg ;
reg  oeh ;
reg  oei ;
reg  oej ;
reg  oek ;
reg  oel ;
reg  oem ;
reg  oen ;
reg  oeo ;
reg  oep ;
reg  ofa ;
reg  ofb ;
reg  ofc ;
reg  ofd ;
reg  ofe ;
reg  off ;
reg  ofg ;
reg  ofh ;
reg  ofi ;
reg  ofj ;
reg  ofk ;
reg  ofl ;
reg  ofm ;
reg  ofn ;
reg  ofo ;
reg  ofp ;
reg  oga ;
reg  ogb ;
reg  ogc ;
reg  ogd ;
reg  oge ;
reg  ogf ;
reg  ogg ;
reg  ogh ;
reg  ogi ;
reg  ogj ;
reg  ogk ;
reg  ogl ;
reg  ogm ;
reg  ogn ;
reg  ogo ;
reg  ogp ;
reg  oha ;
reg  ohb ;
reg  ohc ;
reg  ohd ;
reg  ohe ;
reg  ohf ;
reg  ohg ;
reg  ohh ;
reg  ohi ;
reg  ohj ;
reg  ohk ;
reg  ohl ;
reg  ohm ;
reg  ohn ;
reg  oho ;
reg  ohp ;
reg  OJA ;
reg  OJB ;
reg  OJD ;
reg  OJF ;
reg  OKA ;
reg  OKB ;
reg  OKC ;
reg  OKG ;
reg  OKH ;
reg  oki ;
reg  okj ;
reg  okk ;
reg  okl ;
reg  okm ;
reg  okn ;
reg  oko ;
reg  okp ;
reg  okq ;
reg  okr ;
reg  oks ;
reg  OKT ;
reg  oku ;
reg  okv ;
reg  okw ;
reg  okx ;
reg  PAA ;
reg  PAB ;
reg  PAC ;
reg  PAD ;
reg  PAE ;
reg  PAF ;
reg  PAG ;
reg  PAH ;
reg  PAI ;
reg  PBA ;
reg  PBB ;
reg  PBC ;
reg  PBD ;
reg  PBE ;
reg  PBF ;
reg  PBG ;
reg  PBH ;
reg  PBI ;
reg  PCA ;
reg  PCB ;
reg  PCC ;
reg  PCD ;
reg  PCE ;
reg  PCF ;
reg  PCG ;
reg  PCH ;
reg  PCI ;
reg  PDA ;
reg  PDB ;
reg  PDC ;
reg  PDD ;
reg  PDE ;
reg  PDF ;
reg  PDG ;
reg  PDH ;
reg  PDI ;
reg  PEA ;
reg  PEB ;
reg  PEC ;
reg  PFA ;
reg  PFB ;
reg  PFC ;
reg  PGA ;
reg  PGB ;
reg  PGC ;
reg  PXA ;
reg  PXB ;
reg  PXC ;
reg  qaa ;
reg  qab ;
reg  qac ;
reg  qad ;
reg  QAE ;
reg  QBA ;
reg  QBB ;
reg  QBC ;
reg  QBD ;
reg  QBE ;
reg  QCA ;
reg  QCB ;
reg  QCC ;
reg  QCD ;
reg  QCE ;
reg  QCI ;
reg  QCJ ;
reg  QCK ;
reg  QCL ;
reg  QDA ;
reg  qdb ;
reg  QDC ;
reg  QDD ;
reg  QDE ;
reg  QEB ;
reg  qec ;
reg  qed ;
reg  qee ;
reg  QEF ;
reg  qha ;
reg  qhb ;
reg  qhc ;
reg  qhd ;
reg  qja ;
reg  QJB ;
reg  QJC ;
reg  QJD ;
reg  QJE ;
reg  QJF ;
reg  QJG ;
reg  QJH ;
reg  QJI ;
reg  qjj ;
reg  QJK ;
reg  QJL ;
reg  QJM ;
reg  QJN ;
reg  QJO ;
reg  QJP ;
reg  QJQ ;
reg  QJR ;
reg  QJS ;
reg  QJT ;
reg  QJU ;
reg  QJV ;
reg  QJW ;
reg  QJX ;
reg  QJY ;
reg  qjz ;
reg  QKA ;
reg  QKB ;
reg  qla ;
reg  qlb ;
reg  qld ;
reg  QLF ;
reg  QLG ;
reg  QLH ;
reg  qlj ;
reg  QPA ;
reg  QPB ;
reg  QPC ;
reg  QPD ;
reg  QQA ;
reg  QQB ;
reg  QQC ;
reg  QQD ;
reg  QQE ;
reg  QQF ;
reg  QQG ;
reg  QQH ;
reg  QQI ;
reg  QQJ ;
reg  QQK ;
reg  QQL ;
reg  QQM ;
reg  QQN ;
reg  QQO ;
reg  TAA ;
reg  TAB ;
reg  TAC ;
reg  TAD ;
reg  TAE ;
reg  TAF ;
reg  TAG ;
reg  TAH ;
reg  TBA ;
reg  TBB ;
reg  TBC ;
reg  TBD ;
reg  TBE ;
reg  TBF ;
reg  TBG ;
reg  TBH ;
reg  TCA ;
reg  TCB ;
reg  TCC ;
reg  TCD ;
reg  TCE ;
reg  TCF ;
reg  TCG ;
reg  TCH ;
reg  TDA ;
reg  TDB ;
reg  TDC ;
reg  TDD ;
reg  TDE ;
reg  TDF ;
reg  TDG ;
reg  TDH ;
reg  TEA ;
reg  TEB ;
reg  TEC ;
reg  TED ;
reg  TEE ;
reg  TEF ;
reg  TEG ;
reg  TEH ;
reg  tfa ;
reg  tfb ;
reg  tfc ;
reg  tfd ;
reg  tfe ;
reg  tff ;
reg  tfg ;
reg  tfh ;
reg  TGA ;
reg  TGB ;
reg  TGC ;
reg  TGD ;
reg  TGE ;
reg  TGF ;
reg  TGG ;
reg  TGH ;
reg  TJA ;
reg  TJB ;
reg  TJC ;
reg  TJD ;
reg  TMA ;
reg  UAA ;
reg  UAB ;
reg  UAC ;
reg  UAD ;
reg  UAE ;
reg  UAF ;
reg  UAG ;
reg  UAH ;
reg  UAI ;
reg  UAJ ;
reg  UAK ;
reg  UAL ;
reg  UAM ;
reg  UAN ;
reg  UAO ;
reg  UAP ;
reg  uba ;
reg  ubb ;
reg  ubc ;
reg  ubd ;
reg  ube ;
reg  ubf ;
reg  UBG ;
reg  UBH ;
reg  ubi ;
reg  ubj ;
reg  ubk ;
reg  ubl ;
reg  ubm ;
reg  ubn ;
reg  UBO ;
reg  UBP ;
reg  UCA ;
reg  UCB ;
reg  UCC ;
reg  UCD ;
reg  UCE ;
reg  UCF ;
reg  UCG ;
reg  UCH ;
reg  UCI ;
reg  UCJ ;
reg  UCK ;
reg  UCL ;
reg  UCM ;
reg  UCN ;
reg  UCO ;
reg  UCP ;
reg  uda ;
reg  udb ;
reg  udc ;
reg  udd ;
reg  ude ;
reg  udf ;
reg  UDG ;
reg  UDH ;
reg  udi ;
reg  udj ;
reg  udk ;
reg  udl ;
reg  udm ;
reg  udn ;
reg  UDO ;
reg  UDP ;
reg  UEA ;
reg  UEB ;
reg  UEC ;
reg  UED ;
reg  UEE ;
reg  UEF ;
reg  UEG ;
reg  UEH ;
reg  UEI ;
reg  UEJ ;
reg  UEK ;
reg  UEL ;
reg  UEM ;
reg  UEN ;
reg  UEO ;
reg  UEP ;
reg  ufa ;
reg  ufb ;
reg  ufc ;
reg  ufd ;
reg  ufe ;
reg  uff ;
reg  UFG ;
reg  UFH ;
reg  ufi ;
reg  ufj ;
reg  ufk ;
reg  ufl ;
reg  ufm ;
reg  ufn ;
reg  UFO ;
reg  UFP ;
reg  UGA ;
reg  UGB ;
reg  UGC ;
reg  UGD ;
reg  UGE ;
reg  UGF ;
reg  UGG ;
reg  UGH ;
reg  UGI ;
reg  UGJ ;
reg  UGK ;
reg  UGL ;
reg  UGM ;
reg  UGN ;
reg  UGO ;
reg  UGP ;
reg  uha ;
reg  uhb ;
reg  uhc ;
reg  uhd ;
reg  uhe ;
reg  uhf ;
reg  UHG ;
reg  UHH ;
reg  uhi ;
reg  uhj ;
reg  uhk ;
reg  uhl ;
reg  uhm ;
reg  uhn ;
reg  UHO ;
reg  UHP ;
reg  UIA ;
reg  UIB ;
reg  UIC ;
reg  UID ;
reg  UIE ;
reg  UIF ;
reg  UIG ;
reg  UIH ;
reg  UII ;
reg  UIJ ;
reg  UIK ;
reg  UIL ;
reg  UIM ;
reg  UIN ;
reg  UIO ;
reg  UIP ;
reg  uja ;
reg  ujb ;
reg  ujc ;
reg  ujd ;
reg  uje ;
reg  ujf ;
reg  UJG ;
reg  UJH ;
reg  uji ;
reg  ujj ;
reg  ujk ;
reg  ujl ;
reg  ujm ;
reg  ujn ;
reg  UJO ;
reg  UJP ;
reg  UKA ;
reg  UKB ;
reg  UKC ;
reg  UKD ;
reg  UKE ;
reg  UKF ;
reg  UKG ;
reg  UKH ;
reg  UKI ;
reg  UKJ ;
reg  UKK ;
reg  UKL ;
reg  UKM ;
reg  UKN ;
reg  UKO ;
reg  UKP ;
reg  ula ;
reg  ulb ;
reg  ulc ;
reg  uld ;
reg  ule ;
reg  ulf ;
reg  ULG ;
reg  ULH ;
reg  uli ;
reg  ulj ;
reg  ulk ;
reg  ull ;
reg  ulm ;
reg  uln ;
reg  ULO ;
reg  ULP ;
reg  UMA ;
reg  UMB ;
reg  UMC ;
reg  UMD ;
reg  UME ;
reg  UMF ;
reg  UMG ;
reg  UMH ;
reg  UMI ;
reg  UMJ ;
reg  UMK ;
reg  UML ;
reg  UMM ;
reg  UMN ;
reg  UMO ;
reg  UMP ;
reg  una ;
reg  unb ;
reg  unc ;
reg  und ;
reg  une ;
reg  unf ;
reg  UNG ;
reg  UNH ;
reg  uni ;
reg  unj ;
reg  unk ;
reg  unl ;
reg  unm ;
reg  unn ;
reg  UNO ;
reg  UNP ;
reg  UOA ;
reg  UOB ;
reg  UOC ;
reg  UOD ;
reg  UOE ;
reg  UOF ;
reg  UOG ;
reg  UOH ;
reg  UOI ;
reg  UOJ ;
reg  UOK ;
reg  UOL ;
reg  UOM ;
reg  UON ;
reg  UOO ;
reg  UOP ;
reg  upa ;
reg  upb ;
reg  upc ;
reg  upd ;
reg  upe ;
reg  upf ;
reg  UPG ;
reg  UPH ;
reg  upi ;
reg  upj ;
reg  upk ;
reg  upl ;
reg  upm ;
reg  upn ;
reg  UPO ;
reg  UPP ;
reg  VAA ;
reg  VAB ;
reg  VAC ;
reg  VAD ;
reg  VAE ;
reg  VAF ;
reg  VAG ;
reg  VAH ;
reg  VAI ;
reg  VAJ ;
reg  VAK ;
reg  VAL ;
reg  VAM ;
reg  VAN ;
reg  VAO ;
reg  VAP ;
reg  VBA ;
reg  VBB ;
reg  VBC ;
reg  VBD ;
reg  VBE ;
reg  VBF ;
reg  VBG ;
reg  VBH ;
reg  VBI ;
reg  VBJ ;
reg  VBK ;
reg  VBL ;
reg  VBM ;
reg  VBN ;
reg  VBO ;
reg  VBP ;
reg  VCA ;
reg  VCB ;
reg  VCC ;
reg  VCD ;
reg  VCE ;
reg  VCF ;
reg  VCG ;
reg  VCH ;
reg  VCI ;
reg  VCJ ;
reg  VCK ;
reg  VCL ;
reg  VCM ;
reg  VCN ;
reg  VCO ;
reg  VCP ;
reg  VDA ;
reg  VDB ;
reg  VDC ;
reg  VDD ;
reg  VDE ;
reg  VDF ;
reg  VDG ;
reg  VDH ;
reg  VDI ;
reg  VDJ ;
reg  VDK ;
reg  VDL ;
reg  VDM ;
reg  VDN ;
reg  VDO ;
reg  VDP ;
reg  WAA ;
reg  WAB ;
reg  WAC ;
reg  WAD ;
reg  WAE ;
reg  WAF ;
reg  WAG ;
reg  WAH ;
reg  WAI ;
reg  WAJ ;
reg  WAK ;
reg  WAL ;
reg  WAM ;
reg  WAN ;
reg  WAO ;
reg  WAP ;
reg  WBA ;
reg  WBB ;
reg  WBC ;
reg  WBD ;
reg  WBE ;
reg  WBF ;
reg  WBG ;
reg  WBH ;
reg  WBI ;
reg  WBJ ;
reg  WBK ;
reg  WBL ;
reg  WBM ;
reg  WBN ;
reg  WBO ;
reg  WBP ;
reg  WCA ;
reg  WCB ;
reg  WCC ;
reg  WCD ;
reg  WCE ;
reg  WCF ;
reg  WCG ;
reg  WCH ;
reg  WCI ;
reg  WCJ ;
reg  WCK ;
reg  WCL ;
reg  WCM ;
reg  WCN ;
reg  WCO ;
reg  WCP ;
reg  WDA ;
reg  WDB ;
reg  WDC ;
reg  WDD ;
reg  WDE ;
reg  WDF ;
reg  WDG ;
reg  WDH ;
reg  WDI ;
reg  WDJ ;
reg  WDK ;
reg  WDL ;
reg  WDM ;
reg  WDN ;
reg  WDO ;
reg  WDP ;
reg  WEA ;
reg  WEB ;
reg  WEC ;
reg  WED ;
reg  WEE ;
reg  WEF ;
reg  WEG ;
reg  WEH ;
reg  WEI ;
reg  WEJ ;
reg  WEK ;
reg  WEL ;
reg  WEM ;
reg  WEN ;
reg  WEO ;
reg  WEP ;
reg  WFA ;
reg  WFB ;
reg  WFC ;
reg  WFD ;
reg  WFE ;
reg  WFF ;
reg  WFG ;
reg  WFH ;
reg  WFI ;
reg  WFJ ;
reg  WFK ;
reg  WFL ;
reg  WFM ;
reg  WFN ;
reg  WFO ;
reg  WFP ;
reg  WGA ;
reg  WGB ;
reg  WGC ;
reg  WGD ;
reg  WGE ;
reg  WGF ;
reg  WGG ;
reg  WGH ;
reg  WGI ;
reg  WGJ ;
reg  WGK ;
reg  WGL ;
reg  WGM ;
reg  WGN ;
reg  WGO ;
reg  WGP ;
reg  WHA ;
reg  WHB ;
reg  WHC ;
reg  WHD ;
reg  WHE ;
reg  WHF ;
reg  WHG ;
reg  WHH ;
reg  WHI ;
reg  WHJ ;
reg  WHK ;
reg  WHL ;
reg  WHM ;
reg  WHN ;
reg  WHO ;
reg  WHP ;
reg  WIA ;
reg  WIB ;
reg  WIC ;
reg  WID ;
reg  WIE ;
reg  WIF ;
reg  WIG ;
reg  WIH ;
reg  WII ;
reg  WIJ ;
reg  WIK ;
reg  WIL ;
reg  WIM ;
reg  WIN ;
reg  WIO ;
reg  WIP ;
reg  WJA ;
reg  WJB ;
reg  WJC ;
reg  WJD ;
reg  WJE ;
reg  WJF ;
reg  WJG ;
reg  WJH ;
reg  WJI ;
reg  WJJ ;
reg  WJK ;
reg  WJL ;
reg  WJM ;
reg  WJN ;
reg  WJO ;
reg  WJP ;
reg  WKA ;
reg  WKB ;
reg  WKC ;
reg  WKD ;
reg  WKE ;
reg  WKF ;
reg  WKG ;
reg  WKH ;
reg  WKI ;
reg  WKJ ;
reg  WKK ;
reg  WKL ;
reg  WKM ;
reg  WKN ;
reg  WKO ;
reg  WKP ;
reg  WLA ;
reg  WLB ;
reg  WLC ;
reg  WLD ;
reg  WLE ;
reg  WLF ;
reg  WLG ;
reg  WLH ;
reg  WLI ;
reg  WLJ ;
reg  WLK ;
reg  WLL ;
reg  WLM ;
reg  WLN ;
reg  WLO ;
reg  WLP ;
reg  WMA ;
reg  WMB ;
reg  WMC ;
reg  WMD ;
reg  WME ;
reg  WMF ;
reg  WMG ;
reg  WMH ;
reg  WMI ;
reg  WMJ ;
reg  WMK ;
reg  WML ;
reg  WMM ;
reg  WMN ;
reg  WMO ;
reg  WMP ;
reg  WNA ;
reg  WNB ;
reg  WNC ;
reg  WND ;
reg  WNE ;
reg  WNF ;
reg  WNG ;
reg  WNH ;
reg  WNI ;
reg  WNJ ;
reg  WNK ;
reg  WNL ;
reg  WNM ;
reg  WNN ;
reg  WNO ;
reg  WNP ;
reg  WOA ;
reg  WOB ;
reg  WOC ;
reg  WOD ;
reg  WOE ;
reg  WOF ;
reg  WOG ;
reg  WOH ;
reg  WOI ;
reg  WOJ ;
reg  WOK ;
reg  WOL ;
reg  WOM ;
reg  WON ;
reg  WOO ;
reg  WOP ;
reg  WPA ;
reg  WPB ;
reg  WPC ;
reg  WPD ;
reg  WPE ;
reg  WPF ;
reg  WPG ;
reg  WPH ;
reg  WPI ;
reg  WPJ ;
reg  WPK ;
reg  WPL ;
reg  WPM ;
reg  WPN ;
reg  WPO ;
reg  WPP ;
wire  daa ;
wire  dab ;
wire  dac ;
wire  dad ;
wire  dae ;
wire  daf ;
wire  dag ;
wire  dah ;
wire  dai ;
wire  daj ;
wire  dak ;
wire  dal ;
wire  dam ;
wire  dan ;
wire  dao ;
wire  dba ;
wire  dbb ;
wire  dbc ;
wire  dbe ;
wire  dbf ;
wire  dbg ;
wire  dbi ;
wire  dbj ;
wire  dbk ;
wire  dbm ;
wire  dbn ;
wire  dbo ;
wire  eaa ;
wire  eab ;
wire  eac ;
wire  ead ;
wire  eae ;
wire  EBA ;
wire  EBB ;
wire  EBC ;
wire  eca ;
wire  ecb ;
wire  ecc ;
wire  eda ;
wire  edb ;
wire  edc ;
wire  eea ;
wire  eeb ;
wire  eec ;
wire  efa ;
wire  efb ;
wire  faa ;
wire  fab ;
wire  fac ;
wire  fad ;
wire  fae ;
wire  fba ;
wire  fbb ;
wire  fbc ;
wire  fbd ;
wire  fbe ;
wire  gaa ;
wire  GAA ;
wire  gab ;
wire  GAB ;
wire  gac ;
wire  GAC ;
wire  gad ;
wire  GAD ;
wire  gae ;
wire  GAE ;
wire  gaf ;
wire  GAF ;
wire  gag ;
wire  GAG ;
wire  gah ;
wire  GAH ;
wire  gba ;
wire  GBA ;
wire  gbb ;
wire  GBB ;
wire  gbc ;
wire  GBC ;
wire  gbd ;
wire  GBD ;
wire  gbe ;
wire  GBE ;
wire  gbf ;
wire  GBF ;
wire  gbg ;
wire  GBG ;
wire  gbh ;
wire  GBH ;
wire  gca ;
wire  GCA ;
wire  gcb ;
wire  GCB ;
wire  gcc ;
wire  GCC ;
wire  gcd ;
wire  GCD ;
wire  gce ;
wire  GCE ;
wire  gcf ;
wire  GCF ;
wire  gcg ;
wire  GCG ;
wire  gch ;
wire  GCH ;
wire  gda ;
wire  GDA ;
wire  gdb ;
wire  GDB ;
wire  gdc ;
wire  GDC ;
wire  gdd ;
wire  GDD ;
wire  gde ;
wire  GDE ;
wire  gdf ;
wire  GDF ;
wire  gdg ;
wire  GDG ;
wire  gdh ;
wire  GDH ;
wire  gea ;
wire  GEA ;
wire  geb ;
wire  GEB ;
wire  gec ;
wire  GEC ;
wire  ged ;
wire  GED ;
wire  gee ;
wire  GEE ;
wire  gef ;
wire  GEF ;
wire  geg ;
wire  GEG ;
wire  geh ;
wire  GEH ;
wire  gfa ;
wire  GFA ;
wire  gfb ;
wire  GFB ;
wire  gfc ;
wire  GFC ;
wire  gfd ;
wire  GFD ;
wire  gfe ;
wire  GFE ;
wire  gff ;
wire  GFF ;
wire  gfg ;
wire  GFG ;
wire  gfh ;
wire  GFH ;
wire  gga ;
wire  GGA ;
wire  ggb ;
wire  GGB ;
wire  ggc ;
wire  GGC ;
wire  ggd ;
wire  GGD ;
wire  gge ;
wire  GGE ;
wire  ggf ;
wire  GGF ;
wire  ggg ;
wire  GGG ;
wire  ggh ;
wire  GGH ;
wire  gha ;
wire  GHA ;
wire  ghb ;
wire  GHB ;
wire  ghc ;
wire  GHC ;
wire  ghd ;
wire  GHD ;
wire  ghe ;
wire  GHE ;
wire  ghf ;
wire  GHF ;
wire  ghg ;
wire  GHG ;
wire  ghh ;
wire  GHH ;
wire  gia ;
wire  GIA ;
wire  gib ;
wire  GIB ;
wire  gic ;
wire  GIC ;
wire  gid ;
wire  GID ;
wire  gie ;
wire  GIE ;
wire  gif ;
wire  GIF ;
wire  gig ;
wire  GIG ;
wire  gih ;
wire  GIH ;
wire  gja ;
wire  GJA ;
wire  gjb ;
wire  GJB ;
wire  gjc ;
wire  GJC ;
wire  gjd ;
wire  GJD ;
wire  gje ;
wire  GJE ;
wire  gjf ;
wire  GJF ;
wire  gjg ;
wire  GJG ;
wire  gjh ;
wire  GJH ;
wire  gka ;
wire  GKA ;
wire  gkb ;
wire  GKB ;
wire  gkc ;
wire  GKC ;
wire  gkd ;
wire  GKD ;
wire  gke ;
wire  GKE ;
wire  gkf ;
wire  GKF ;
wire  gkg ;
wire  GKG ;
wire  gkh ;
wire  GKH ;
wire  gla ;
wire  GLA ;
wire  glb ;
wire  GLB ;
wire  glc ;
wire  GLC ;
wire  gld ;
wire  GLD ;
wire  gle ;
wire  GLE ;
wire  glf ;
wire  GLF ;
wire  glg ;
wire  GLG ;
wire  glh ;
wire  GLH ;
wire  gma ;
wire  GMA ;
wire  gmb ;
wire  GMB ;
wire  gmc ;
wire  GMC ;
wire  gmd ;
wire  GMD ;
wire  gme ;
wire  GME ;
wire  gmf ;
wire  GMF ;
wire  gmg ;
wire  GMG ;
wire  gmh ;
wire  GMH ;
wire  gna ;
wire  GNA ;
wire  gnb ;
wire  GNB ;
wire  gnc ;
wire  GNC ;
wire  gnd ;
wire  GND ;
wire  gne ;
wire  GNE ;
wire  gnf ;
wire  GNF ;
wire  gng ;
wire  GNG ;
wire  gnh ;
wire  GNH ;
wire  goa ;
wire  GOA ;
wire  gob ;
wire  GOB ;
wire  goc ;
wire  GOC ;
wire  god ;
wire  GOD ;
wire  goe ;
wire  GOE ;
wire  gof ;
wire  GOF ;
wire  gog ;
wire  GOG ;
wire  goh ;
wire  GOH ;
wire  gpa ;
wire  GPA ;
wire  gpb ;
wire  GPB ;
wire  gpc ;
wire  GPC ;
wire  gpd ;
wire  GPD ;
wire  gpe ;
wire  GPE ;
wire  gpf ;
wire  GPF ;
wire  gpg ;
wire  GPG ;
wire  gph ;
wire  GPH ;
wire  iaa ;
wire  iab ;
wire  iac ;
wire  iad ;
wire  iae ;
wire  iaf ;
wire  iag ;
wire  iah ;
wire  iai ;
wire  iaj ;
wire  iak ;
wire  ial ;
wire  iam ;
wire  ian ;
wire  iao ;
wire  iap ;
wire  iba ;
wire  ibb ;
wire  ibc ;
wire  ibd ;
wire  ibe ;
wire  ibf ;
wire  ibg ;
wire  ibh ;
wire  ibi ;
wire  ibj ;
wire  ibk ;
wire  ibl ;
wire  ibm ;
wire  ibn ;
wire  ibo ;
wire  ibp ;
wire  ica ;
wire  icb ;
wire  icc ;
wire  icd ;
wire  ice ;
wire  icf ;
wire  icg ;
wire  ich ;
wire  ici ;
wire  icj ;
wire  ick ;
wire  icl ;
wire  icm ;
wire  icn ;
wire  ico ;
wire  icp ;
wire  ida ;
wire  idb ;
wire  idc ;
wire  idd ;
wire  ide ;
wire  idf ;
wire  idg ;
wire  idh ;
wire  idi ;
wire  idj ;
wire  idk ;
wire  idl ;
wire  idm ;
wire  idn ;
wire  ido ;
wire  idp ;
wire  iea ;
wire  ieb ;
wire  iec ;
wire  ied ;
wire  iee ;
wire  ief ;
wire  ieg ;
wire  ieh ;
wire  iei ;
wire  iej ;
wire  ifa ;
wire  ifb ;
wire  ifc ;
wire  ifd ;
wire  ife ;
wire  iga ;
wire  igb ;
wire  igc ;
wire  iha ;
wire  ihb ;
wire  ija ;
wire  ijb ;
wire  ijd ;
wire  ije ;
wire  ijf ;
wire  ijg ;
wire  izz ;
wire  jaa ;
wire  JAA ;
wire  jab ;
wire  JAB ;
wire  jac ;
wire  JAC ;
wire  jad ;
wire  JAD ;
wire  jba ;
wire  JBA ;
wire  jbb ;
wire  JBB ;
wire  jbc ;
wire  JBC ;
wire  jbd ;
wire  JBD ;
wire  jca ;
wire  JCA ;
wire  jcb ;
wire  JCB ;
wire  jcc ;
wire  JCC ;
wire  jcd ;
wire  JCD ;
wire  jda ;
wire  JDA ;
wire  jdb ;
wire  JDB ;
wire  jdc ;
wire  JDC ;
wire  jdd ;
wire  JDD ;
wire  jea ;
wire  JEA ;
wire  jeb ;
wire  JEB ;
wire  jec ;
wire  JEC ;
wire  jed ;
wire  JED ;
wire  jee ;
wire  JEE ;
wire  jef ;
wire  JEF ;
wire  jfa ;
wire  JFA ;
wire  jfb ;
wire  JFB ;
wire  jfc ;
wire  JFC ;
wire  jga ;
wire  JGA ;
wire  jgb ;
wire  JGB ;
wire  jgc ;
wire  JGC ;
wire  jge ;
wire  JGE ;
wire  jgf ;
wire  JGF ;
wire  jgg ;
wire  JGG ;
wire  jha ;
wire  JHA ;
wire  jhb ;
wire  JHB ;
wire  jhc ;
wire  JHC ;
wire  jia ;
wire  JIA ;
wire  jib ;
wire  JIB ;
wire  jic ;
wire  JIC ;
wire  jid ;
wire  JID ;
wire  jja ;
wire  JJA ;
wire  jjb ;
wire  JJB ;
wire  jjc ;
wire  JJC ;
wire  jjd ;
wire  JJD ;
wire  jje ;
wire  JJE ;
wire  jjf ;
wire  JJF ;
wire  jjg ;
wire  JJG ;
wire  jjh ;
wire  JJH ;
wire  jji ;
wire  JJI ;
wire  jjj ;
wire  JJJ ;
wire  jjs ;
wire  JJS ;
wire  jjt ;
wire  JJT ;
wire  jju ;
wire  JJU ;
wire  jjv ;
wire  JJV ;
wire  jjw ;
wire  JJW ;
wire  jjx ;
wire  JJX ;
wire  jjy ;
wire  JJY ;
wire  jjz ;
wire  JJZ ;
wire  jla ;
wire  JLA ;
wire  jlb ;
wire  JLB ;
wire  jlc ;
wire  JLC ;
wire  jld ;
wire  JLD ;
wire  jle ;
wire  JLE ;
wire  jlf ;
wire  JLF ;
wire  jlx ;
wire  JLX ;
wire  jma ;
wire  JMA ;
wire  jmb ;
wire  JMB ;
wire  jmc ;
wire  JMC ;
wire  jna ;
wire  JNA ;
wire  jnb ;
wire  JNB ;
wire  jnc ;
wire  JNC ;
wire  jnd ;
wire  JND ;
wire  jpc ;
wire  JPC ;
wire  jpd ;
wire  JPD ;
wire  jpe ;
wire  JPE ;
wire  jpf ;
wire  JPF ;
wire  jpg ;
wire  JPG ;
wire  jxa ;
wire  JXA ;
wire  jxb ;
wire  JXB ;
wire  kaa ;
wire  KAA ;
wire  kab ;
wire  KAB ;
wire  kac ;
wire  KAC ;
wire  kad ;
wire  KAD ;
wire  kae ;
wire  KAE ;
wire  kaf ;
wire  KAF ;
wire  kag ;
wire  KAG ;
wire  kah ;
wire  KAH ;
wire  kai ;
wire  KAI ;
wire  kaj ;
wire  KAJ ;
wire  kak ;
wire  KAK ;
wire  kal ;
wire  KAL ;
wire  kam ;
wire  KAM ;
wire  kan ;
wire  KAN ;
wire  kao ;
wire  KAO ;
wire  kap ;
wire  KAP ;
wire  kba ;
wire  KBA ;
wire  kbb ;
wire  KBB ;
wire  kbc ;
wire  KBC ;
wire  kbd ;
wire  KBD ;
wire  kbe ;
wire  KBE ;
wire  kbf ;
wire  KBF ;
wire  kbg ;
wire  KBG ;
wire  kbh ;
wire  KBH ;
wire  kbi ;
wire  KBI ;
wire  kbj ;
wire  KBJ ;
wire  kbk ;
wire  KBK ;
wire  kbl ;
wire  KBL ;
wire  kbm ;
wire  KBM ;
wire  kbn ;
wire  KBN ;
wire  kbo ;
wire  KBO ;
wire  kbp ;
wire  KBP ;
wire  kca ;
wire  KCA ;
wire  kcb ;
wire  KCB ;
wire  kcc ;
wire  KCC ;
wire  kcd ;
wire  KCD ;
wire  kce ;
wire  KCE ;
wire  kcf ;
wire  KCF ;
wire  kcg ;
wire  KCG ;
wire  kch ;
wire  KCH ;
wire  kci ;
wire  KCI ;
wire  kcj ;
wire  KCJ ;
wire  kck ;
wire  KCK ;
wire  kcl ;
wire  KCL ;
wire  kcm ;
wire  KCM ;
wire  kcn ;
wire  KCN ;
wire  kco ;
wire  KCO ;
wire  kcp ;
wire  KCP ;
wire  kda ;
wire  KDA ;
wire  kdb ;
wire  KDB ;
wire  kdc ;
wire  KDC ;
wire  kdd ;
wire  KDD ;
wire  kde ;
wire  KDE ;
wire  kdf ;
wire  KDF ;
wire  kdg ;
wire  KDG ;
wire  kdh ;
wire  KDH ;
wire  kdi ;
wire  KDI ;
wire  kdj ;
wire  KDJ ;
wire  kdk ;
wire  KDK ;
wire  kdl ;
wire  KDL ;
wire  kdm ;
wire  KDM ;
wire  kdn ;
wire  KDN ;
wire  kdo ;
wire  KDO ;
wire  kdp ;
wire  KDP ;
wire  oaa ;
wire  oab ;
wire  oac ;
wire  oad ;
wire  oae ;
wire  oaf ;
wire  oag ;
wire  oah ;
wire  oai ;
wire  oaj ;
wire  oak ;
wire  oal ;
wire  oam ;
wire  oan ;
wire  oao ;
wire  oap ;
wire  oba ;
wire  obb ;
wire  obc ;
wire  obd ;
wire  obe ;
wire  obf ;
wire  obg ;
wire  obh ;
wire  obi ;
wire  obj ;
wire  obk ;
wire  obl ;
wire  obm ;
wire  obn ;
wire  obo ;
wire  obp ;
wire  oca ;
wire  ocb ;
wire  occ ;
wire  ocd ;
wire  oce ;
wire  ocf ;
wire  ocg ;
wire  och ;
wire  oci ;
wire  ocj ;
wire  ock ;
wire  ocl ;
wire  ocm ;
wire  ocn ;
wire  oco ;
wire  ocp ;
wire  oda ;
wire  odb ;
wire  odc ;
wire  odd ;
wire  ode ;
wire  odf ;
wire  odg ;
wire  odh ;
wire  odi ;
wire  odj ;
wire  odk ;
wire  odl ;
wire  odm ;
wire  odn ;
wire  odo ;
wire  odp ;
wire  OEA ;
wire  OEB ;
wire  OEC ;
wire  OED ;
wire  OEE ;
wire  OEF ;
wire  OEG ;
wire  OEH ;
wire  OEI ;
wire  OEJ ;
wire  OEK ;
wire  OEL ;
wire  OEM ;
wire  OEN ;
wire  OEO ;
wire  OEP ;
wire  OFA ;
wire  OFB ;
wire  OFC ;
wire  OFD ;
wire  OFE ;
wire  OFF ;
wire  OFG ;
wire  OFH ;
wire  OFI ;
wire  OFJ ;
wire  OFK ;
wire  OFL ;
wire  OFM ;
wire  OFN ;
wire  OFO ;
wire  OFP ;
wire  OGA ;
wire  OGB ;
wire  OGC ;
wire  OGD ;
wire  OGE ;
wire  OGF ;
wire  OGG ;
wire  OGH ;
wire  OGI ;
wire  OGJ ;
wire  OGK ;
wire  OGL ;
wire  OGM ;
wire  OGN ;
wire  OGO ;
wire  OGP ;
wire  OHA ;
wire  OHB ;
wire  OHC ;
wire  OHD ;
wire  OHE ;
wire  OHF ;
wire  OHG ;
wire  OHH ;
wire  OHI ;
wire  OHJ ;
wire  OHK ;
wire  OHL ;
wire  OHM ;
wire  OHN ;
wire  OHO ;
wire  OHP ;
wire  oja ;
wire  ojb ;
wire  ojd ;
wire  ojf ;
wire  oka ;
wire  okb ;
wire  okc ;
wire  okg ;
wire  okh ;
wire  OKI ;
wire  OKJ ;
wire  OKK ;
wire  OKL ;
wire  OKM ;
wire  OKN ;
wire  OKO ;
wire  OKP ;
wire  OKQ ;
wire  OKR ;
wire  OKS ;
wire  okt ;
wire  OKU ;
wire  OKV ;
wire  OKW ;
wire  OKX ;
wire  paa ;
wire  pab ;
wire  pac ;
wire  pad ;
wire  pae ;
wire  paf ;
wire  pag ;
wire  pah ;
wire  pai ;
wire  pba ;
wire  pbb ;
wire  pbc ;
wire  pbd ;
wire  pbe ;
wire  pbf ;
wire  pbg ;
wire  pbh ;
wire  pbi ;
wire  pca ;
wire  pcb ;
wire  pcc ;
wire  pcd ;
wire  pce ;
wire  pcf ;
wire  pcg ;
wire  pch ;
wire  pci ;
wire  pda ;
wire  pdb ;
wire  pdc ;
wire  pdd ;
wire  pde ;
wire  pdf ;
wire  pdg ;
wire  pdh ;
wire  pdi ;
wire  pea ;
wire  peb ;
wire  pec ;
wire  pfa ;
wire  pfb ;
wire  pfc ;
wire  pga ;
wire  pgb ;
wire  pgc ;
wire  pxa ;
wire  pxb ;
wire  pxc ;
wire  QAA ;
wire  QAB ;
wire  QAC ;
wire  QAD ;
wire  qae ;
wire  qba ;
wire  qbb ;
wire  qbc ;
wire  qbd ;
wire  qbe ;
wire  qca ;
wire  qcb ;
wire  qcc ;
wire  qcd ;
wire  qce ;
wire  qci ;
wire  qcj ;
wire  qck ;
wire  qcl ;
wire  qda ;
wire  QDB ;
wire  qdc ;
wire  qdd ;
wire  qde ;
wire  qeb ;
wire  QEC ;
wire  QED ;
wire  QEE ;
wire  qef ;
wire  QHA ;
wire  QHB ;
wire  QHC ;
wire  QHD ;
wire  QJA ;
wire  qjb ;
wire  qjc ;
wire  qjd ;
wire  qje ;
wire  qjf ;
wire  qjg ;
wire  qjh ;
wire  qji ;
wire  QJJ ;
wire  qjk ;
wire  qjl ;
wire  qjm ;
wire  qjn ;
wire  qjo ;
wire  qjp ;
wire  qjq ;
wire  qjr ;
wire  qjs ;
wire  qjt ;
wire  qju ;
wire  qjv ;
wire  qjw ;
wire  qjx ;
wire  qjy ;
wire  QJZ ;
wire  qka ;
wire  qkb ;
wire  QLA ;
wire  QLB ;
wire  QLD ;
wire  qlf ;
wire  qlg ;
wire  qlh ;
wire  QLJ ;
wire  qpa ;
wire  qpb ;
wire  qpc ;
wire  qpd ;
wire  qqa ;
wire  qqb ;
wire  qqc ;
wire  qqd ;
wire  qqe ;
wire  qqf ;
wire  qqg ;
wire  qqh ;
wire  qqi ;
wire  qqj ;
wire  qqk ;
wire  qql ;
wire  qqm ;
wire  qqn ;
wire  qqo ;
wire  taa ;
wire  tab ;
wire  tac ;
wire  tad ;
wire  tae ;
wire  taf ;
wire  tag ;
wire  tah ;
wire  tba ;
wire  tbb ;
wire  tbc ;
wire  tbd ;
wire  tbe ;
wire  tbf ;
wire  tbg ;
wire  tbh ;
wire  tca ;
wire  tcb ;
wire  tcc ;
wire  tcd ;
wire  tce ;
wire  tcf ;
wire  tcg ;
wire  tch ;
wire  tda ;
wire  tdb ;
wire  tdc ;
wire  tdd ;
wire  tde ;
wire  tdf ;
wire  tdg ;
wire  tdh ;
wire  tea ;
wire  teb ;
wire  tec ;
wire  ted ;
wire  tee ;
wire  tef ;
wire  teg ;
wire  teh ;
wire  TFA ;
wire  TFB ;
wire  TFC ;
wire  TFD ;
wire  TFE ;
wire  TFF ;
wire  TFG ;
wire  TFH ;
wire  tga ;
wire  tgb ;
wire  tgc ;
wire  tgd ;
wire  tge ;
wire  tgf ;
wire  tgg ;
wire  tgh ;
wire  tja ;
wire  tjb ;
wire  tjc ;
wire  tjd ;
wire  tma ;
wire  uaa ;
wire  uab ;
wire  uac ;
wire  uad ;
wire  uae ;
wire  uaf ;
wire  uag ;
wire  uah ;
wire  uai ;
wire  uaj ;
wire  uak ;
wire  ual ;
wire  uam ;
wire  uan ;
wire  uao ;
wire  uap ;
wire  UBA ;
wire  UBB ;
wire  UBC ;
wire  UBD ;
wire  UBE ;
wire  UBF ;
wire  ubg ;
wire  ubh ;
wire  UBI ;
wire  UBJ ;
wire  UBK ;
wire  UBL ;
wire  UBM ;
wire  UBN ;
wire  ubo ;
wire  ubp ;
wire  uca ;
wire  ucb ;
wire  ucc ;
wire  ucd ;
wire  uce ;
wire  ucf ;
wire  ucg ;
wire  uch ;
wire  uci ;
wire  ucj ;
wire  uck ;
wire  ucl ;
wire  ucm ;
wire  ucn ;
wire  uco ;
wire  ucp ;
wire  UDA ;
wire  UDB ;
wire  UDC ;
wire  UDD ;
wire  UDE ;
wire  UDF ;
wire  udg ;
wire  udh ;
wire  UDI ;
wire  UDJ ;
wire  UDK ;
wire  UDL ;
wire  UDM ;
wire  UDN ;
wire  udo ;
wire  udp ;
wire  uea ;
wire  ueb ;
wire  uec ;
wire  ued ;
wire  uee ;
wire  uef ;
wire  ueg ;
wire  ueh ;
wire  uei ;
wire  uej ;
wire  uek ;
wire  uel ;
wire  uem ;
wire  uen ;
wire  ueo ;
wire  uep ;
wire  UFA ;
wire  UFB ;
wire  UFC ;
wire  UFD ;
wire  UFE ;
wire  UFF ;
wire  ufg ;
wire  ufh ;
wire  UFI ;
wire  UFJ ;
wire  UFK ;
wire  UFL ;
wire  UFM ;
wire  UFN ;
wire  ufo ;
wire  ufp ;
wire  uga ;
wire  ugb ;
wire  ugc ;
wire  ugd ;
wire  uge ;
wire  ugf ;
wire  ugg ;
wire  ugh ;
wire  ugi ;
wire  ugj ;
wire  ugk ;
wire  ugl ;
wire  ugm ;
wire  ugn ;
wire  ugo ;
wire  ugp ;
wire  UHA ;
wire  UHB ;
wire  UHC ;
wire  UHD ;
wire  UHE ;
wire  UHF ;
wire  uhg ;
wire  uhh ;
wire  UHI ;
wire  UHJ ;
wire  UHK ;
wire  UHL ;
wire  UHM ;
wire  UHN ;
wire  uho ;
wire  uhp ;
wire  uia ;
wire  uib ;
wire  uic ;
wire  uid ;
wire  uie ;
wire  uif ;
wire  uig ;
wire  uih ;
wire  uii ;
wire  uij ;
wire  uik ;
wire  uil ;
wire  uim ;
wire  uin ;
wire  uio ;
wire  uip ;
wire  UJA ;
wire  UJB ;
wire  UJC ;
wire  UJD ;
wire  UJE ;
wire  UJF ;
wire  ujg ;
wire  ujh ;
wire  UJI ;
wire  UJJ ;
wire  UJK ;
wire  UJL ;
wire  UJM ;
wire  UJN ;
wire  ujo ;
wire  ujp ;
wire  uka ;
wire  ukb ;
wire  ukc ;
wire  ukd ;
wire  uke ;
wire  ukf ;
wire  ukg ;
wire  ukh ;
wire  uki ;
wire  ukj ;
wire  ukk ;
wire  ukl ;
wire  ukm ;
wire  ukn ;
wire  uko ;
wire  ukp ;
wire  ULA ;
wire  ULB ;
wire  ULC ;
wire  ULD ;
wire  ULE ;
wire  ULF ;
wire  ulg ;
wire  ulh ;
wire  ULI ;
wire  ULJ ;
wire  ULK ;
wire  ULL ;
wire  ULM ;
wire  ULN ;
wire  ulo ;
wire  ulp ;
wire  uma ;
wire  umb ;
wire  umc ;
wire  umd ;
wire  ume ;
wire  umf ;
wire  umg ;
wire  umh ;
wire  umi ;
wire  umj ;
wire  umk ;
wire  uml ;
wire  umm ;
wire  umn ;
wire  umo ;
wire  ump ;
wire  UNA ;
wire  UNB ;
wire  UNC ;
wire  UND ;
wire  UNE ;
wire  UNF ;
wire  ung ;
wire  unh ;
wire  UNI ;
wire  UNJ ;
wire  UNK ;
wire  UNL ;
wire  UNM ;
wire  UNN ;
wire  uno ;
wire  unp ;
wire  uoa ;
wire  uob ;
wire  uoc ;
wire  uod ;
wire  uoe ;
wire  uof ;
wire  uog ;
wire  uoh ;
wire  uoi ;
wire  uoj ;
wire  uok ;
wire  uol ;
wire  uom ;
wire  uon ;
wire  uoo ;
wire  uop ;
wire  UPA ;
wire  UPB ;
wire  UPC ;
wire  UPD ;
wire  UPE ;
wire  UPF ;
wire  upg ;
wire  uph ;
wire  UPI ;
wire  UPJ ;
wire  UPK ;
wire  UPL ;
wire  UPM ;
wire  UPN ;
wire  upo ;
wire  upp ;
wire  vaa ;
wire  vab ;
wire  vac ;
wire  vad ;
wire  vae ;
wire  vaf ;
wire  vag ;
wire  vah ;
wire  vai ;
wire  vaj ;
wire  vak ;
wire  val ;
wire  vam ;
wire  van ;
wire  vao ;
wire  vap ;
wire  vba ;
wire  vbb ;
wire  vbc ;
wire  vbd ;
wire  vbe ;
wire  vbf ;
wire  vbg ;
wire  vbh ;
wire  vbi ;
wire  vbj ;
wire  vbk ;
wire  vbl ;
wire  vbm ;
wire  vbn ;
wire  vbo ;
wire  vbp ;
wire  vca ;
wire  vcb ;
wire  vcc ;
wire  vcd ;
wire  vce ;
wire  vcf ;
wire  vcg ;
wire  vch ;
wire  vci ;
wire  vcj ;
wire  vck ;
wire  vcl ;
wire  vcm ;
wire  vcn ;
wire  vco ;
wire  vcp ;
wire  vda ;
wire  vdb ;
wire  vdc ;
wire  vdd ;
wire  vde ;
wire  vdf ;
wire  vdg ;
wire  vdh ;
wire  vdi ;
wire  vdj ;
wire  vdk ;
wire  vdl ;
wire  vdm ;
wire  vdn ;
wire  vdo ;
wire  vdp ;
wire  waa ;
wire  wab ;
wire  wac ;
wire  wad ;
wire  wae ;
wire  waf ;
wire  wag ;
wire  wah ;
wire  wai ;
wire  waj ;
wire  wak ;
wire  wal ;
wire  wam ;
wire  wan ;
wire  wao ;
wire  wap ;
wire  wba ;
wire  wbb ;
wire  wbc ;
wire  wbd ;
wire  wbe ;
wire  wbf ;
wire  wbg ;
wire  wbh ;
wire  wbi ;
wire  wbj ;
wire  wbk ;
wire  wbl ;
wire  wbm ;
wire  wbn ;
wire  wbo ;
wire  wbp ;
wire  wca ;
wire  wcb ;
wire  wcc ;
wire  wcd ;
wire  wce ;
wire  wcf ;
wire  wcg ;
wire  wch ;
wire  wci ;
wire  wcj ;
wire  wck ;
wire  wcl ;
wire  wcm ;
wire  wcn ;
wire  wco ;
wire  wcp ;
wire  wda ;
wire  wdb ;
wire  wdc ;
wire  wdd ;
wire  wde ;
wire  wdf ;
wire  wdg ;
wire  wdh ;
wire  wdi ;
wire  wdj ;
wire  wdk ;
wire  wdl ;
wire  wdm ;
wire  wdn ;
wire  wdo ;
wire  wdp ;
wire  wea ;
wire  web ;
wire  wec ;
wire  wed ;
wire  wee ;
wire  wef ;
wire  weg ;
wire  weh ;
wire  wei ;
wire  wej ;
wire  wek ;
wire  wel ;
wire  wem ;
wire  wen ;
wire  weo ;
wire  wep ;
wire  wfa ;
wire  wfb ;
wire  wfc ;
wire  wfd ;
wire  wfe ;
wire  wff ;
wire  wfg ;
wire  wfh ;
wire  wfi ;
wire  wfj ;
wire  wfk ;
wire  wfl ;
wire  wfm ;
wire  wfn ;
wire  wfo ;
wire  wfp ;
wire  wga ;
wire  wgb ;
wire  wgc ;
wire  wgd ;
wire  wge ;
wire  wgf ;
wire  wgg ;
wire  wgh ;
wire  wgi ;
wire  wgj ;
wire  wgk ;
wire  wgl ;
wire  wgm ;
wire  wgn ;
wire  wgo ;
wire  wgp ;
wire  wha ;
wire  whb ;
wire  whc ;
wire  whd ;
wire  whe ;
wire  whf ;
wire  whg ;
wire  whh ;
wire  whi ;
wire  whj ;
wire  whk ;
wire  whl ;
wire  whm ;
wire  whn ;
wire  who ;
wire  whp ;
wire  wia ;
wire  wib ;
wire  wic ;
wire  wid ;
wire  wie ;
wire  wif ;
wire  wig ;
wire  wih ;
wire  wii ;
wire  wij ;
wire  wik ;
wire  wil ;
wire  wim ;
wire  win ;
wire  wio ;
wire  wip ;
wire  wja ;
wire  wjb ;
wire  wjc ;
wire  wjd ;
wire  wje ;
wire  wjf ;
wire  wjg ;
wire  wjh ;
wire  wji ;
wire  wjj ;
wire  wjk ;
wire  wjl ;
wire  wjm ;
wire  wjn ;
wire  wjo ;
wire  wjp ;
wire  wka ;
wire  wkb ;
wire  wkc ;
wire  wkd ;
wire  wke ;
wire  wkf ;
wire  wkg ;
wire  wkh ;
wire  wki ;
wire  wkj ;
wire  wkk ;
wire  wkl ;
wire  wkm ;
wire  wkn ;
wire  wko ;
wire  wkp ;
wire  wla ;
wire  wlb ;
wire  wlc ;
wire  wld ;
wire  wle ;
wire  wlf ;
wire  wlg ;
wire  wlh ;
wire  wli ;
wire  wlj ;
wire  wlk ;
wire  wll ;
wire  wlm ;
wire  wln ;
wire  wlo ;
wire  wlp ;
wire  wma ;
wire  wmb ;
wire  wmc ;
wire  wmd ;
wire  wme ;
wire  wmf ;
wire  wmg ;
wire  wmh ;
wire  wmi ;
wire  wmj ;
wire  wmk ;
wire  wml ;
wire  wmm ;
wire  wmn ;
wire  wmo ;
wire  wmp ;
wire  wna ;
wire  wnb ;
wire  wnc ;
wire  wnd ;
wire  wne ;
wire  wnf ;
wire  wng ;
wire  wnh ;
wire  wni ;
wire  wnj ;
wire  wnk ;
wire  wnl ;
wire  wnm ;
wire  wnn ;
wire  wno ;
wire  wnp ;
wire  woa ;
wire  wob ;
wire  woc ;
wire  wod ;
wire  woe ;
wire  wof ;
wire  wog ;
wire  woh ;
wire  woi ;
wire  woj ;
wire  wok ;
wire  wol ;
wire  wom ;
wire  won ;
wire  woo ;
wire  wop ;
wire  wpa ;
wire  wpb ;
wire  wpc ;
wire  wpd ;
wire  wpe ;
wire  wpf ;
wire  wpg ;
wire  wph ;
wire  wpi ;
wire  wpj ;
wire  wpk ;
wire  wpl ;
wire  wpm ;
wire  wpn ;
wire  wpo ;
wire  wpp ;
wire  ZZI ;
wire  ZZO ;

wire NAA ;
wire NAB ;
wire NAC ;
wire NAD ;
wire NAE ;
wire NAF ;
wire NAG ;
wire NAH ;
wire NAI ;
wire NAJ ;
wire NAK ;
wire NAL ;
wire NAM ;
wire NAN ;
wire NAO ;
wire NAP ;
wire NBA ;
wire NBB ;
wire NBC ;
wire NBD ;
wire NBE ;
wire NBF ;
wire NBG ;
wire NBH ;
wire NBI ;
wire NBJ ;
wire NBK ;
wire NBL ;
wire NBM ;
wire NBN ;
wire NBO ;
wire NBP ;
wire NCA ;
wire NCB ;
wire NCC ;
wire NCD ;
wire NCE ;
wire NCF ;
wire NCG ;
wire NCH ;
wire NCI ;
wire NCJ ;
wire NCK ;
wire NCL ;
wire NCM ;
wire NCN ;
wire NCO ;
wire NCP ;
wire NDA ;
wire NDB ;
wire NDC ;
wire NDD ;
wire NDE ;
wire NDF ;
wire NDG ;
wire NDH ;
wire NDI ;
wire NDJ ;
wire NDK ;
wire NDL ;
wire NDM ;
wire NDN ;
wire NDO ;
wire NDP ;
wire NEA ;
wire NEB ;
wire NEC ;
wire NED ;
wire NEE ;
wire NEF ;
wire NEG ;
wire NEH ;
wire NEI ;
wire NEJ ;
wire NEK ;
wire NEL ;
wire NEM ;
wire NEN ;
wire NEO ;
wire NEP ;
wire NFA ;
wire NFB ;
wire NFC ;
wire NFD ;
wire NFE ;
wire NFF ;
wire NFG ;
wire NFH ;
wire NFI ;
wire NFJ ;
wire NFK ;
wire NFL ;
wire NFM ;
wire NFN ;
wire NFO ;
wire NFP ;
wire NGA ;
wire NGB ;
wire NGC ;
wire NGD ;
wire NGE ;
wire NGF ;
wire NGG ;
wire NGH ;
wire NGI ;
wire NGJ ;
wire NGK ;
wire NGL ;
wire NGM ;
wire NGN ;
wire NGO ;
wire NGP ;
wire NHA ;
wire NHB ;
wire NHC ;
wire NHD ;
wire NHE ;
wire NHF ;
wire NHG ;
wire NHH ;
wire NHI ;
wire NHJ ;
wire NHK ;
wire NHL ;
wire NHM ;
wire NHN ;
wire NHO ;
wire NHP ;
wire NIA ;
wire NIB ;
wire NIC ;
wire NID ;
wire NIE ;
wire NIF ;
wire NIG ;
wire NIH ;
wire NII ;
wire NIJ ;
wire NIK ;
wire NIL ;
wire NIM ;
wire NIN ;
wire NIO ;
wire NIP ;
wire NJA ;
wire NJB ;
wire NJC ;
wire NJD ;
wire NJE ;
wire NJF ;
wire NJG ;
wire NJH ;
wire NJI ;
wire NJJ ;
wire NJK ;
wire NJL ;
wire NJM ;
wire NJN ;
wire NJO ;
wire NJP ;
wire NKA ;
wire NKB ;
wire NKC ;
wire NKD ;
wire NKE ;
wire NKF ;
wire NKG ;
wire NKH ;
wire NKI ;
wire NKJ ;
wire NKK ;
wire NKL ;
wire NKM ;
wire NKN ;
wire NKO ;
wire NKP ;
wire NKA ;
wire NKB ;
wire NKC ;
wire NKD ;
wire NKE ;
wire NKF ;
wire NKG ;
wire NKH ;
wire NKI ;
wire NKJ ;
wire NKK ;
wire NKL ;
wire NKM ;
wire NKN ;
wire NKO ;
wire NKP ;
wire NLA ;
wire NLB ;
wire NLC ;
wire NLD ;
wire NLE ;
wire NLF ;
wire NLG ;
wire NLH ;
wire NLI ;
wire NLJ ;
wire NLK ;
wire NLL ;
wire NLM ;
wire NLN ;
wire NLO ;
wire NLP ;
wire NMA ;
wire NMB ;
wire NMC ;
wire NMD ;
wire NME ;
wire NMF ;
wire NMG ;
wire NMH ;
wire NMI ;
wire NMJ ;
wire NMK ;
wire NML ;
wire NMM ;
wire NMN ;
wire NMO ;
wire NMP ;
wire NNA ;
wire NNB ;
wire NNC ;
wire NND ;
wire NNE ;
wire NNF ;
wire NNG ;
wire NNH ;
wire NNI ;
wire NNJ ;
wire NNK ;
wire NNL ;
wire NNM ;
wire NNN ;
wire NNO ;
wire NNP ;
wire NOA ;
wire NOB ;
wire NOC ;
wire NOD ;
wire NOE ;
wire NOF ;
wire NOG ;
wire NOH ;
wire NOI ;
wire NOJ ;
wire NOK ;
wire NOL ;
wire NOM ;
wire NON ;
wire NOO ;
wire NOP ;
wire NPA ;
wire NPB ;
wire NPC ;
wire NPD ;
wire NPE ;
wire NPF ;
wire NPG ;
wire NPH ;
wire NPI ;
wire NPJ ;
wire NPK ;
wire NPL ;
wire NPM ;
wire NPN ;
wire NPO ;
wire NPP ;              

wire RAA ;
wire RAB ;
wire RAC ;
wire RAD ;
wire RAE ;
wire RAF ;
wire RAG ;
wire RAH ;
wire RAI ;
wire RAJ ;
wire RAK ;
wire RAL ;
wire RAM ;
wire RAN ;
wire RAO ;
wire RAP ;
wire RBA ;
wire RBB ;
wire RBC ;
wire RBD ;
wire RBE ;
wire RBF ;
wire RBG ;
wire RBH ;
wire RBI ;
wire RBJ ;
wire RBK ;
wire RBL ;
wire RBM ;
wire RBN ;
wire RBO ;
wire RBP ;
wire RCA ;
wire RCB ;
wire RCC ;
wire RCD ;
wire RCE ;
wire RCF ;
wire RCG ;
wire RCH ;
wire RCI ;
wire RCJ ;
wire RCK ;
wire RCL ;
wire RCM ;
wire RCN ;
wire RCO ;
wire RCP ;
wire RDA ;
wire RDB ;
wire RDC ;
wire RDD ;
wire RDE ;
wire RDF ;
wire RDG ;
wire RDH ;
wire RDI ;
wire RDJ ;
wire RDK ;
wire RDL ;
wire RDM ;
wire RDN ;
wire RDO ;
wire RDP ;
wire REA ;
wire REB ;
wire REC ;
wire RED ;
wire REE ;
wire REFF  ;
wire REG ;
wire REH ;
wire REI ;
wire REJ ;
wire REK ;
wire REL ;
wire REM ;
wire REN ;
wire REO ;
wire REP ;
wire RFA ;
wire RFB ;
wire RFC ;
wire RFD ;
wire RFE ;
wire RFF ;
wire RFG ;
wire RFH ;
wire RFI ;
wire RFJ ;
wire RFK ;
wire RFL ;
wire RFM ;
wire RFN ;
wire RFO ;
wire RFP ;
wire RGA ;
wire RGB ;
wire RGC ;
wire RGD ;
wire RGE ;
wire RGF ;
wire RGG ;
wire RGH ;
wire RGI ;
wire RGJ ;
wire RGK ;
wire RGL ;
wire RGM ;
wire RGN ;
wire RGO ;
wire RGP ;
wire RHA ;
wire RHB ;
wire RHC ;
wire RHD ;
wire RHE ;
wire RHF ;
wire RHG ;
wire RHH ;
wire RHI ;
wire RHJ ;
wire RHK ;
wire RHL ;
wire RHM ;
wire RHN ;
wire RHO ;
wire RHP ;
wire RIA ;
wire RIB ;
wire RIC ;
wire RID ;
wire RIE ;
wire RIF ;
wire RIG ;
wire RIH ;
wire RII ;
wire RIJ ;
wire RIK ;
wire RIL ;
wire RIM ;
wire RIN ;
wire RIO ;
wire RIP ;
wire RJA ;
wire RJB ;
wire RJC ;
wire RJD ;
wire RJE ;
wire RJF ;
wire RJG ;
wire RJH ;
wire RJI ;
wire RJJ ;
wire RJK ;
wire RJL ;
wire RJM ;
wire RJN ;
wire RJO ;
wire RJP ;
wire RKA ;
wire RKB ;
wire RKC ;
wire RKD ;
wire RKE ;
wire RKF ;
wire RKG ;
wire RKH ;
wire RKI ;
wire RKJ ;
wire RKK ;
wire RKL ;
wire RKM ;
wire RKN ;
wire RKO ;
wire RKP ;
wire RKA ;
wire RKB ;
wire RKC ;
wire RKD ;
wire RKE ;
wire RKF ;
wire RKG ;
wire RKH ;
wire RKI ;
wire RKJ ;
wire RKK ;
wire RKL ;
wire RKM ;
wire RKN ;
wire RKO ;
wire RKP ;
wire RLA ;
wire RLB ;
wire RLC ;
wire RLD ;
wire RLE ;
wire RLF ;
wire RLG ;
wire RLH ;
wire RLI ;
wire RLJ ;
wire RLK ;
wire RLL ;
wire RLM ;
wire RLN ;
wire RLO ;
wire RLP ;
wire RMA ;
wire RMB ;
wire RMC ;
wire RMD ;
wire RME ;
wire RMF ;
wire RMG ;
wire RMH ;
wire RMI ;
wire RMJ ;
wire RMK ;
wire RML ;
wire RMM ;
wire RMN ;
wire RMO ;
wire RMP ;
wire RNA ;
wire RNB ;
wire RNC ;
wire RND ;
wire RNE ;
wire RNF ;
wire RNG ;
wire RNH ;
wire RNI ;
wire RNJ ;
wire RNK ;
wire RNL ;
wire RNM ;
wire RNN ;
wire RNO ;
wire RNP ;
wire ROA ;
wire ROB ;
wire ROC ;
wire ROD ;
wire ROE ;
wire ROF ;
wire ROG ;
wire ROH ;
wire ROI ;
wire ROJ ;
wire ROK ;
wire ROL ;
wire ROM ;
wire RON ;
wire ROO ;
wire ROP ;
wire RPA ;
wire RPB ;
wire RPC ;
wire RPD ;
wire RPE ;
wire RPF ;
wire RPG ;
wire RPH ;
wire RPI ;
wire RPJ ;
wire RPK ;
wire RPL ;
wire RPM ;
wire RPN ;
wire RPO ;
wire RPP ;

wire SAA ;
wire SAB ;
wire SAC ;
wire SAD ;
wire SAE ;
wire SAF ;
wire SAG ;
wire SAH ;
wire SAI ;
wire SAJ ;
wire SAK ;
wire SAL ;
wire SAM ;
wire SAN ;
wire SAO ;
wire SAP ;
wire SBA ;
wire SBB ;
wire SBC ;
wire SBD ;
wire SBE ;
wire SBF ;
wire SBG ;
wire SBH ;
wire SBI ;
wire SBJ ;
wire SBK ;
wire SBL ;
wire SBM ;
wire SBN ;
wire SBO ;
wire SBP ;
wire SCA ;
wire SCB ;
wire SCC ;
wire SCD ;
wire SCE ;
wire SCF ;
wire SCG ;
wire SCH ;
wire SCI ;
wire SCJ ;
wire SCK ;
wire SCL ;
wire SCM ;
wire SCN ;
wire SCO ;
wire SCP ;
wire SDA ;
wire SDB ;
wire SDC ;
wire SDD ;
wire SDE ;
wire SDF ;
wire SDG ;
wire SDH ;
wire SDI ;
wire SDJ ;
wire SDK ;
wire SDL ;
wire SDM ;
wire SDN ;
wire SDO ;
wire SDP ;
wire SEA ;
wire SEB ;
wire SEC ;
wire SED ;
wire SEE ;
wire SEF ;
wire SEG ;
wire SEH ;
wire SEI ;
wire SEJ ;
wire SEK ;
wire SEL ;
wire SEM ;
wire SEN ;
wire SEO ;
wire SEP ;
wire SFA ;
wire SFB ;
wire SFC ;
wire SFD ;
wire SFE ;
wire SFF ;
wire SFG ;
wire SFH ;
wire SFI ;
wire SFJ ;
wire SFK ;
wire SFL ;
wire SFM ;
wire SFN ;
wire SFO ;
wire SFP ;
wire SGA ;
wire SGB ;
wire SGC ;
wire SGD ;
wire SGE ;
wire SGF ;
wire SGG ;
wire SGH ;
wire SGI ;
wire SGJ ;
wire SGK ;
wire SGL ;
wire SGM ;
wire SGN ;
wire SGO ;
wire SGP ;
wire SHA ;
wire SHB ;
wire SHC ;
wire SHD ;
wire SHE ;
wire SHF ;
wire SHG ;
wire SHH ;
wire SHI ;
wire SHJ ;
wire SHK ;
wire SHL ;
wire SHM ;
wire SHN ;
wire SHO ;
wire SHP ;
wire SIA ;
wire SIB ;
wire SIC ;
wire SID ;
wire SIE ;
wire SIF ;
wire SIG ;
wire SIH ;
wire SII ;
wire SIJ ;
wire SIK ;
wire SIL ;
wire SIM ;
wire SIN ;
wire SIO ;
wire SIP ;
wire SJA ;
wire SJB ;
wire SJC ;
wire SJD ;
wire SJE ;
wire SJF ;
wire SJG ;
wire SJH ;
wire SJI ;
wire SJJ ;
wire SJK ;
wire SJL ;
wire SJM ;
wire SJN ;
wire SJO ;
wire SJP ;
wire SKA ;
wire SKB ;
wire SKC ;
wire SKD ;
wire SKE ;
wire SKF ;
wire SKG ;
wire SKH ;
wire SKI ;
wire SKJ ;
wire SKK ;
wire SKL ;
wire SKM ;
wire SKN ;
wire SKO ;
wire SKP ;
wire SKA ;
wire SKB ;
wire SKC ;
wire SKD ;
wire SKE ;
wire SKF ;
wire SKG ;
wire SKH ;
wire SKI ;
wire SKJ ;
wire SKK ;
wire SKL ;
wire SKM ;
wire SKN ;
wire SKO ;
wire SKP ;
wire SLA ;
wire SLB ;
wire SLC ;
wire SLD ;
wire SLE ;
wire SLF ;
wire SLG ;
wire SLH ;
wire SLI ;
wire SLJ ;
wire SLK ;
wire SLL ;
wire SLM ;
wire SLN ;
wire SLO ;
wire SLP ;
wire SMA ;
wire SMB ;
wire SMC ;
wire SMD ;
wire SME ;
wire SMF ;
wire SMG ;
wire SMH ;
wire SMI ;
wire SMJ ;
wire SMK ;
wire SML ;
wire SMM ;
wire SMN ;
wire SMO ;
wire SMP ;
wire SNA ;
wire SNB ;
wire SNC ;
wire SND ;
wire SNE ;
wire SNF ;
wire SNG ;
wire SNH ;
wire SNI ;
wire SNJ ;
wire SNK ;
wire SNL ;
wire SNM ;
wire SNN ;
wire SNO ;
wire SNP ;
wire SOA ;
wire SOB ;
wire SOC ;
wire SOD ;
wire SOE ;
wire SOF ;
wire SOG ;
wire SOH ;
wire SOI ;
wire SOJ ;
wire SOK ;
wire SOL ;
wire SOM ;
wire SON ;
wire SOO ;
wire SOP ;
wire SPA ;
wire SPB ;
wire SPC ;
wire SPD ;
wire SPE ;
wire SPF ;
wire SPG ;
wire SPH ;
wire SPI ;
wire SPJ ;
wire SPK ;
wire SPL ;
wire SPM ;
wire SPN ;
wire SPO ;
wire SPP ;

wire XAA ;
wire XAB ;
wire XAC ;
wire XAD ;
wire XAE ;
wire XAF ;
wire XAG ;
wire XAH ;
wire XAI ;
wire XAJ ;
wire XAK ;
wire XAL ;
wire XAM ;
wire XAN ;
wire XAO ;
wire XAP ;
wire XBA ;
wire XBB ;
wire XBC ;
wire XBD ;
wire XBE ;
wire XBF ;
wire XBG ;
wire XBH ;
wire XBI ;
wire XBJ ;
wire XBK ;
wire XBL ;
wire XBM ;
wire XBN ;
wire XBO ;
wire XBP ;
wire XCA ;
wire XCB ;
wire XCC ;
wire XCD ;
wire XCE ;
wire XCF ;
wire XCG ;
wire XCH ;
wire XCI ;
wire XCJ ;
wire XCK ;
wire XCL ;
wire XCM ;
wire XCN ;
wire XCO ;
wire XCP ;
wire XDA ;
wire XDB ;
wire XDC ;
wire XDD ;
wire XDE ;
wire XDF ;
wire XDG ;
wire XDH ;
wire XDI ;
wire XDJ ;
wire XDK ;
wire XDL ;
wire XDM ;
wire XDN ;
wire XDO ;
wire XDP ;
wire XEA ;
wire XEB ;
wire XEC ;
wire XED ;
wire XEE ;
wire XEF ;
wire XEG ;
wire XEH ;
wire XEI ;
wire XEJ ;
wire XEK ;
wire XEL ;
wire XEM ;
wire XEN ;
wire XEO ;
wire XEP ;
wire XFA ;
wire XFB ;
wire XFC ;
wire XFD ;
wire XFE ;
wire XFF ;
wire XFG ;
wire XFH ;
wire XFI ;
wire XFJ ;
wire XFK ;
wire XFL ;
wire XFM ;
wire XFN ;
wire XFO ;
wire XFP ;
wire XGA ;
wire XGB ;
wire XGC ;
wire XGD ;
wire XGE ;
wire XGF ;
wire XGG ;
wire XGH ;
wire XGI ;
wire XGJ ;
wire XGK ;
wire XGL ;
wire XGM ;
wire XGN ;
wire XGO ;
wire XGP ;
wire XHA ;
wire XHB ;
wire XHC ;
wire XHD ;
wire XHE ;
wire XHF ;
wire XHG ;
wire XHH ;
wire XHI ;
wire XHJ ;
wire XHK ;
wire XHL ;
wire XHM ;
wire XHN ;
wire XHO ;
wire XHP ;
wire XIA ;
wire XIB ;
wire XIC ;
wire XID ;
wire XIE ;
wire XIF ;
wire XIG ;
wire XIH ;
wire XII ;
wire XIJ ;
wire XIK ;
wire XIL ;
wire XIM ;
wire XIN ;
wire XIO ;
wire XIP ;
wire XJA ;
wire XJB ;
wire XJC ;
wire XJD ;
wire XJE ;
wire XJF ;
wire XJG ;
wire XJH ;
wire XJI ;
wire XJJ ;
wire XJK ;
wire XJL ;
wire XJM ;
wire XJN ;
wire XJO ;
wire XJP ;
wire XKA ;
wire XKB ;
wire XKC ;
wire XKD ;
wire XKE ;
wire XKF ;
wire XKG ;
wire XKH ;
wire XKI ;
wire XKJ ;
wire XKK ;
wire XKL ;
wire XKM ;
wire XKN ;
wire XKO ;
wire XKP ;
wire XKA ;
wire XKB ;
wire XKC ;
wire XKD ;
wire XKE ;
wire XKF ;
wire XKG ;
wire XKH ;
wire XKI ;
wire XKJ ;
wire XKK ;
wire XKL ;
wire XKM ;
wire XKN ;
wire XKO ;
wire XKP ;
wire XLA ;
wire XLB ;
wire XLC ;
wire XLD ;
wire XLE ;
wire XLF ;
wire XLG ;
wire XLH ;
wire XLI ;
wire XLJ ;
wire XLK ;
wire XLL ;
wire XLM ;
wire XLN ;
wire XLO ;
wire XLP ;
wire XMA ;
wire XMB ;
wire XMC ;
wire XMD ;
wire XME ;
wire XMF ;
wire XMG ;
wire XMH ;
wire XMI ;
wire XMJ ;
wire XMK ;
wire XML ;
wire XMM ;
wire XMN ;
wire XMO ;
wire XMP ;
wire XNA ;
wire XNB ;
wire XNC ;
wire XND ;
wire XNE ;
wire XNF ;
wire XNG ;
wire XNH ;
wire XNI ;
wire XNJ ;
wire XNK ;
wire XNL ;
wire XNM ;
wire XNN ;
wire XNO ;
wire XNP ;
wire XOA ;
wire XOB ;
wire XOC ;
wire XOD ;
wire XOE ;
wire XOF ;
wire XOG ;
wire XOH ;
wire XOI ;
wire XOJ ;
wire XOK ;
wire XOL ;
wire XOM ;
wire XON ;
wire XOO ;
wire XOP ;
wire XPA ;
wire XPB ;
wire XPC ;
wire XPD ;
wire XPE ;
wire XPF ;
wire XPG ;
wire XPH ;
wire XPI ;
wire XPJ ;
wire XPK ;
wire XPL ;
wire XPM ;
wire XPN ;
wire XPO ;
wire XPP ;

wire YAA ;
wire YAB ;
wire YAC ;
wire YAD ;
wire YAE ;
wire YAF ;
wire YAG ;
wire YAH ;
wire YAI ;
wire YAJ ;
wire YAK ;
wire YAL ;
wire YAM ;
wire YAN ;
wire YAO ;
wire YAP ;
wire YBA ;
wire YBB ;
wire YBC ;
wire YBD ;
wire YBE ;
wire YBF ;
wire YBG ;
wire YBH ;
wire YBI ;
wire YBJ ;
wire YBK ;
wire YBL ;
wire YBM ;
wire YBN ;
wire YBO ;
wire YBP ;
wire YCA ;
wire YCB ;
wire YCC ;
wire YCD ;
wire YCE ;
wire YCF ;
wire YCG ;
wire YCH ;
wire YCI ;
wire YCJ ;
wire YCK ;
wire YCL ;
wire YCM ;
wire YCN ;
wire YCO ;
wire YCP ;
wire YDA ;
wire YDB ;
wire YDC ;
wire YDD ;
wire YDE ;
wire YDF ;
wire YDG ;
wire YDH ;
wire YDI ;
wire YDJ ;
wire YDK ;
wire YDL ;
wire YDM ;
wire YDN ;
wire YDO ;
wire YDP ;
wire YEA ;
wire YEB ;
wire YEC ;
wire YED ;
wire YEE ;
wire YEF ;
wire YEG ;
wire YEH ;
wire YEI ;
wire YEJ ;
wire YEK ;
wire YEL ;
wire YEM ;
wire YEN ;
wire YEO ;
wire YEP ;
wire YFA ;
wire YFB ;
wire YFC ;
wire YFD ;
wire YFE ;
wire YFF ;
wire YFG ;
wire YFH ;
wire YFI ;
wire YFJ ;
wire YFK ;
wire YFL ;
wire YFM ;
wire YFN ;
wire YFO ;
wire YFP ;
wire YGA ;
wire YGB ;
wire YGC ;
wire YGD ;
wire YGE ;
wire YGF ;
wire YGG ;
wire YGH ;
wire YGI ;
wire YGJ ;
wire YGK ;
wire YGL ;
wire YGM ;
wire YGN ;
wire YGO ;
wire YGP ;
wire YHA ;
wire YHB ;
wire YHC ;
wire YHD ;
wire YHE ;
wire YHF ;
wire YHG ;
wire YHH ;
wire YHI ;
wire YHJ ;
wire YHK ;
wire YHL ;
wire YHM ;
wire YHN ;
wire YHO ;
wire YHP ;
wire YIA ;
wire YIB ;
wire YIC ;
wire YID ;
wire YIE ;
wire YIF ;
wire YIG ;
wire YIH ;
wire YII ;
wire YIJ ;
wire YIK ;
wire YIL ;
wire YIM ;
wire YIN ;
wire YIO ;
wire YIP ;
wire YJA ;
wire YJB ;
wire YJC ;
wire YJD ;
wire YJE ;
wire YJF ;
wire YJG ;
wire YJH ;
wire YJI ;
wire YJJ ;
wire YJK ;
wire YJL ;
wire YJM ;
wire YJN ;
wire YJO ;
wire YJP ;
wire YKA ;
wire YKB ;
wire YKC ;
wire YKD ;
wire YKE ;
wire YKF ;
wire YKG ;
wire YKH ;
wire YKI ;
wire YKJ ;
wire YKK ;
wire YKL ;
wire YKM ;
wire YKN ;
wire YKO ;
wire YKP ;
wire YKA ;
wire YKB ;
wire YKC ;
wire YKD ;
wire YKE ;
wire YKF ;
wire YKG ;
wire YKH ;
wire YKI ;
wire YKJ ;
wire YKK ;
wire YKL ;
wire YKM ;
wire YKN ;
wire YKO ;
wire YKP ;
wire YLA ;
wire YLB ;
wire YLC ;
wire YLD ;
wire YLE ;
wire YLF ;
wire YLG ;
wire YLH ;
wire YLI ;
wire YLJ ;
wire YLK ;
wire YLL ;
wire YLM ;
wire YLN ;
wire YLO ;
wire YLP ;
wire YMA ;
wire YMB ;
wire YMC ;
wire YMD ;
wire YME ;
wire YMF ;
wire YMG ;
wire YMH ;
wire YMI ;
wire YMJ ;
wire YMK ;
wire YML ;
wire YMM ;
wire YMN ;
wire YMO ;
wire YMP ;
wire YNA ;
wire YNB ;
wire YNC ;
wire YND ;
wire YNE ;
wire YNF ;
wire YNG ;
wire YNH ;
wire YNI ;
wire YNJ ;
wire YNK ;
wire YNL ;
wire YNM ;
wire YNN ;
wire YNO ;
wire YNP ;
wire YOA ;
wire YOB ;
wire YOC ;
wire YOD ;
wire YOE ;
wire YOF ;
wire YOG ;
wire YOH ;
wire YOI ;
wire YOJ ;
wire YOK ;
wire YOL ;
wire YOM ;
wire YON ;
wire YOO ;
wire YOP ;
wire YPA ;
wire YPB ;
wire YPC ;
wire YPD ;
wire YPE ;
wire YPF ;
wire YPG ;
wire YPH ;
wire YPI ;
wire YPJ ;
wire YPK ;
wire YPL ;
wire YPM ;
wire YPN ;
wire YPO ;
wire YPP ;              
assign ZZI = 1'b1;
assign ZZO = 1'b0;
assign uaa = ~UAA;  //complement 
assign uab = ~UAB;  //complement 
assign uac = ~UAC;  //complement 
assign uad = ~UAD;  //complement 
assign uae = ~UAE;  //complement 
assign uaf = ~UAF;  //complement 
assign GAA = uaf & uae ; 
assign gaa = ~GAA ; //complement 
assign GAB = uaf & UAE ; 
assign gab = ~GAB ;  //complement 
assign GAC = UAF & uae ; 
assign gac = ~GAC ;  //complement 
assign GAD = UAF & UAE; 
assign gad = ~GAD; 
assign UBD = ~ubd;  //complement 
assign UBE = ~ube;  //complement 
assign UBF = ~ubf;  //complement 
assign UBA = ~uba;  //complement 
assign UBB = ~ubb;  //complement 
assign UBC = ~ubc;  //complement 
assign GBA = ubf & ube ; 
assign gba = ~GBA ; //complement 
assign GBB = ubf & UBE ; 
assign gbb = ~GBB ;  //complement 
assign GBC = UBF & ube ; 
assign gbc = ~GBC ;  //complement 
assign GBD = UBF & UBE; 
assign gbd = ~GBD; 
assign uca = ~UCA;  //complement 
assign ucb = ~UCB;  //complement 
assign ucc = ~UCC;  //complement 
assign GCA = ucf & uce ; 
assign gca = ~GCA ; //complement 
assign GCB = ucf & UCE ; 
assign gcb = ~GCB ;  //complement 
assign GCC = UCF & uce ; 
assign gcc = ~GCC ;  //complement 
assign GCD = UCF & UCE; 
assign gcd = ~GCD; 
assign ucd = ~UCD;  //complement 
assign uce = ~UCE;  //complement 
assign ucf = ~UCF;  //complement 
assign UDD = ~udd;  //complement 
assign UDE = ~ude;  //complement 
assign UDF = ~udf;  //complement 
assign GDA = udf & ude ; 
assign gda = ~GDA ; //complement 
assign GDB = udf & UDE ; 
assign gdb = ~GDB ;  //complement 
assign GDC = UDF & ude ; 
assign gdc = ~GDC ;  //complement 
assign GDD = UDF & UDE; 
assign gdd = ~GDD; 
assign UDA = ~uda;  //complement 
assign UDB = ~udb;  //complement 
assign UDC = ~udc;  //complement 
assign vaa = ~VAA;  //complement 
assign oaa = ~OAA;  //complement 
assign waa = ~WAA;  //complement 
assign wea = ~WEA;  //complement 
assign wia = ~WIA;  //complement 
assign wma = ~WMA;  //complement 
assign vai = ~VAI;  //complement 
assign oai = ~OAI;  //complement 
assign wai = ~WAI;  //complement 
assign wei = ~WEI;  //complement 
assign wii = ~WII;  //complement 
assign wmi = ~WMI;  //complement 
assign vba = ~VBA;  //complement 
assign oba = ~OBA;  //complement 
assign wba = ~WBA;  //complement 
assign wfa = ~WFA;  //complement 
assign wja = ~WJA;  //complement 
assign wna = ~WNA;  //complement 
assign vbi = ~VBI;  //complement 
assign obi = ~OBI;  //complement 
assign wbi = ~WBI;  //complement 
assign wfi = ~WFI;  //complement 
assign wji = ~WJI;  //complement 
assign wni = ~WNI;  //complement 
assign vca = ~VCA;  //complement 
assign oca = ~OCA;  //complement 
assign wca = ~WCA;  //complement 
assign wga = ~WGA;  //complement 
assign wka = ~WKA;  //complement 
assign woa = ~WOA;  //complement 
assign vci = ~VCI;  //complement 
assign oci = ~OCI;  //complement 
assign wci = ~WCI;  //complement 
assign wgi = ~WGI;  //complement 
assign wki = ~WKI;  //complement 
assign woi = ~WOI;  //complement 
assign vda = ~VDA;  //complement 
assign oda = ~ODA;  //complement 
assign wda = ~WDA;  //complement 
assign wha = ~WHA;  //complement 
assign wla = ~WLA;  //complement 
assign wpa = ~WPA;  //complement 
assign vdi = ~VDI;  //complement 
assign odi = ~ODI;  //complement 
assign wdi = ~WDI;  //complement 
assign whi = ~WHI;  //complement 
assign wli = ~WLI;  //complement 
assign wpi = ~WPI;  //complement 
assign KAA =  WEA & ZZI & TFA  |  VAA & ZZI & TGA  ; 
assign kaa = ~KAA;  //complement 
assign KAI =  WEI & ZZI & TFA  |  VAI & ZZI & TGA  ; 
assign kai = ~KAI;  //complement 
assign taa = ~TAA;  //complement 
assign tba = ~TBA;  //complement 
assign tca = ~TCA;  //complement 
assign tda = ~TDA;  //complement 
assign KBA =  WFA & ZZI & TFB  |  VBA & ZZI & TGB  ; 
assign kba = ~KBA;  //complement 
assign KBI =  WFI & ZZI & TFB  |  VBI & ZZI & TGB  ; 
assign kbi = ~KBI;  //complement 
assign OKJ = ~okj;  //complement 
assign uag = ~UAG;  //complement 
assign uah = ~UAH;  //complement 
assign udg = ~UDG;  //complement 
assign udh = ~UDH;  //complement 
assign OEA = ~oea;  //complement 
assign OEI = ~oei;  //complement 
assign OFA = ~ofa;  //complement 
assign OFI = ~ofi;  //complement 
assign KCA =  WGA & ZZI & TFC  |  VCA & ZZI & TGC  ; 
assign kca = ~KCA;  //complement 
assign KCI =  WGI & ZZI & TFC  |  VCI & ZZI & TGC  ; 
assign kci = ~KCI;  //complement 
assign QHA = ~qha;  //complement 
assign qae = ~QAE;  //complement 
assign qbe = ~QBE;  //complement 
assign qce = ~QCE;  //complement 
assign qde = ~QDE;  //complement 
assign OGA = ~oga;  //complement 
assign OGI = ~ogi;  //complement 
assign OHA = ~oha;  //complement 
assign OHI = ~ohi;  //complement 
assign ubg = ~UBG;  //complement 
assign ubh = ~UBH;  //complement 
assign ucg = ~UCG;  //complement 
assign uch = ~UCH;  //complement 
assign jad = qca & qba ; 
assign JAD = ~jad ; //complement 
assign qba = ~QBA;  //complement 
assign qca = ~QCA;  //complement 
assign qci = ~QCI;  //complement 
assign qda = ~QDA;  //complement 
assign QAA = ~qaa;  //complement 
assign QAB = ~qab;  //complement 
assign KDA =  WHA & ZZI & TFD  |  VDA & ZZI & TGD  ; 
assign kda = ~KDA;  //complement 
assign KDI =  WHI & ZZI & TFD  |  VDI & ZZI & TGD  ; 
assign kdi = ~KDI;  //complement 
assign qpa = ~QPA;  //complement 
assign qpb = ~QPB;  //complement 
assign JAC =  QPA & PAA & PAB  ; 
assign jac = ~JAC;  //complement 
assign JAA =  ZZI & QPA  ; 
assign jaa = ~JAA;  //complement 
assign JAB =  PAA & QPA  ; 
assign jab = ~JAB;  //complement 
assign QAC = ~qac;  //complement 
assign QAD = ~qad;  //complement 
assign paa = ~PAA;  //complement 
assign pad = ~PAD;  //complement 
assign pag = ~PAG;  //complement 
assign pab = ~PAB;  //complement 
assign pae = ~PAE;  //complement 
assign pah = ~PAH;  //complement 
assign pac = ~PAC;  //complement 
assign paf = ~PAF;  //complement 
assign pai = ~PAI;  //complement 
assign uea = ~UEA;  //complement 
assign ueb = ~UEB;  //complement 
assign uec = ~UEC;  //complement 
assign ued = ~UED;  //complement 
assign uee = ~UEE;  //complement 
assign uef = ~UEF;  //complement 
assign GEA = uef & uee ; 
assign gea = ~GEA ; //complement 
assign GEB = uef & UEE ; 
assign geb = ~GEB ;  //complement 
assign GEC = UEF & uee ; 
assign gec = ~GEC ;  //complement 
assign GED = UEF & UEE; 
assign ged = ~GED; 
assign UFD = ~ufd;  //complement 
assign UFE = ~ufe;  //complement 
assign UFF = ~uff;  //complement 
assign UFA = ~ufa;  //complement 
assign UFB = ~ufb;  //complement 
assign UFC = ~ufc;  //complement 
assign GFA = uff & ufe ; 
assign gfa = ~GFA ; //complement 
assign GFB = uff & UFE ; 
assign gfb = ~GFB ;  //complement 
assign GFC = UFF & ufe ; 
assign gfc = ~GFC ;  //complement 
assign GFD = UFF & UFE; 
assign gfd = ~GFD; 
assign uga = ~UGA;  //complement 
assign ugb = ~UGB;  //complement 
assign ugc = ~UGC;  //complement 
assign GGA = ugf & uge ; 
assign gga = ~GGA ; //complement 
assign GGB = ugf & UGE ; 
assign ggb = ~GGB ;  //complement 
assign GGC = UGF & uge ; 
assign ggc = ~GGC ;  //complement 
assign GGD = UGF & UGE; 
assign ggd = ~GGD; 
assign ugd = ~UGD;  //complement 
assign uge = ~UGE;  //complement 
assign ugf = ~UGF;  //complement 
assign UHD = ~uhd;  //complement 
assign UHE = ~uhe;  //complement 
assign UHF = ~uhf;  //complement 
assign GHA = uhf & uhe ; 
assign gha = ~GHA ; //complement 
assign GHB = uhf & UHE ; 
assign ghb = ~GHB ;  //complement 
assign GHC = UHF & uhe ; 
assign ghc = ~GHC ;  //complement 
assign GHD = UHF & UHE; 
assign ghd = ~GHD; 
assign UHA = ~uha;  //complement 
assign UHB = ~uhb;  //complement 
assign UHC = ~uhc;  //complement 
assign vab = ~VAB;  //complement 
assign oab = ~OAB;  //complement 
assign wab = ~WAB;  //complement 
assign web = ~WEB;  //complement 
assign wib = ~WIB;  //complement 
assign wmb = ~WMB;  //complement 
assign vaj = ~VAJ;  //complement 
assign oaj = ~OAJ;  //complement 
assign waj = ~WAJ;  //complement 
assign wej = ~WEJ;  //complement 
assign wij = ~WIJ;  //complement 
assign wmj = ~WMJ;  //complement 
assign vbb = ~VBB;  //complement 
assign obb = ~OBB;  //complement 
assign wbb = ~WBB;  //complement 
assign wfb = ~WFB;  //complement 
assign wjb = ~WJB;  //complement 
assign wnb = ~WNB;  //complement 
assign vbj = ~VBJ;  //complement 
assign obj = ~OBJ;  //complement 
assign wbj = ~WBJ;  //complement 
assign wfj = ~WFJ;  //complement 
assign wjj = ~WJJ;  //complement 
assign wnj = ~WNJ;  //complement 
assign vcb = ~VCB;  //complement 
assign ocb = ~OCB;  //complement 
assign wcb = ~WCB;  //complement 
assign wgb = ~WGB;  //complement 
assign wkb = ~WKB;  //complement 
assign wob = ~WOB;  //complement 
assign vcj = ~VCJ;  //complement 
assign ocj = ~OCJ;  //complement 
assign wcj = ~WCJ;  //complement 
assign wgj = ~WGJ;  //complement 
assign wkj = ~WKJ;  //complement 
assign woj = ~WOJ;  //complement 
assign vdb = ~VDB;  //complement 
assign odb = ~ODB;  //complement 
assign wdb = ~WDB;  //complement 
assign whb = ~WHB;  //complement 
assign wlb = ~WLB;  //complement 
assign wpb = ~WPB;  //complement 
assign vdj = ~VDJ;  //complement 
assign odj = ~ODJ;  //complement 
assign wdj = ~WDJ;  //complement 
assign whj = ~WHJ;  //complement 
assign wlj = ~WLJ;  //complement 
assign wpj = ~WPJ;  //complement 
assign KAB =  WEB & ZZI & TFA  |  VAB & ZZI & TGA  ; 
assign kab = ~KAB;  //complement 
assign KAJ =  WEJ & ZZI & TFA  |  VAJ & ZZI & TGA  ; 
assign kaj = ~KAJ;  //complement 
assign eca = ~ECA;  //complement 
assign eda = ~EDA;  //complement 
assign eea = ~EEA;  //complement 
assign ecb = ~ECB;  //complement 
assign edb = ~EDB;  //complement 
assign eeb = ~EEB;  //complement 
assign ecc = ~ECC;  //complement 
assign edc = ~EDC;  //complement 
assign eec = ~EEC;  //complement 
assign tab = ~TAB;  //complement 
assign tbb = ~TBB;  //complement 
assign tcb = ~TCB;  //complement 
assign tdb = ~TDB;  //complement 
assign jga = qec & ZZI ; 
assign JGA = ~jga ; //complement 
assign jge = qec & qjz ; 
assign JGE = ~jge ;  //complement 
assign JJA =  eda & edb & edc & QQI  ; 
assign jja = ~JJA;  //complement  
assign JJB =  EDA & edb & edc & QQJ  ; 
assign jjb = ~JJB;  //complement 
assign JJC =  eda & EDB & edc & QQK  ; 
assign jjc = ~JJC;  //complement  
assign JJD =  EDA & EDB & edc & QQL  ; 
assign jjd = ~JJD;  //complement 
assign KBB =  WFB & ZZI & TFB  |  VBB & ZZI & TGB  ; 
assign kbb = ~KBB;  //complement 
assign KBJ =  WFJ & ZZI & TFB  |  VBJ & ZZI & TGB  ; 
assign kbj = ~KBJ;  //complement 
assign JGC =  EEB & EEA & QEC  ; 
assign jgc = ~JGC;  //complement 
assign JGB =  EEA & QEC & QEC  ; 
assign jgb = ~JGB;  //complement 
assign JJE =  eda & edb & EDC & QQM  ; 
assign jje = ~JJE;  //complement  
assign JJF =  EDA & edb & EDC & QQN  ; 
assign jjf = ~JJF;  //complement 
assign JJG =  eda & EDB & EDC & QQO  ; 
assign jjg = ~JJG;  //complement  
assign ueg = ~UEG;  //complement 
assign ueh = ~UEH;  //complement 
assign uhg = ~UHG;  //complement 
assign uhh = ~UHH;  //complement 
assign jbd = qcb & qbb ; 
assign JBD = ~jbd ; //complement 
assign JGF =  ZZI & EEA & QEC  |  QJZ  ; 
assign jgf = ~JGF;  //complement 
assign JGG =  EEB & EEA & QEC  |  QJZ  ; 
assign jgg = ~JGG;  //complement 
assign OEB = ~oeb;  //complement 
assign OEJ = ~oej;  //complement 
assign OFB = ~ofb;  //complement 
assign OFJ = ~ofj;  //complement 
assign KCB =  WGB & ZZI & TFC  |  VCB & ZZI & TGC  ; 
assign kcb = ~KCB;  //complement 
assign KCJ =  WGJ & ZZI & TFC  |  VCJ & ZZI & TGC  ; 
assign kcj = ~KCJ;  //complement 
assign QHB = ~qhb;  //complement 
assign OGB = ~ogb;  //complement 
assign OGJ = ~ogj;  //complement 
assign OHB = ~ohb;  //complement 
assign OHJ = ~ohj;  //complement 
assign ufg = ~UFG;  //complement 
assign ufh = ~UFH;  //complement 
assign ugg = ~UGG;  //complement 
assign ugh = ~UGH;  //complement 
assign qbb = ~QBB;  //complement 
assign qcb = ~QCB;  //complement 
assign qcj = ~QCJ;  //complement 
assign QDB = ~qdb;  //complement 
assign OKK = ~okk;  //complement 
assign OKL = ~okl;  //complement 
assign OKM = ~okm;  //complement 
assign OKN = ~okn;  //complement 
assign KDB =  WHB & ZZI & TFD  |  VDB & ZZI & TGD  ; 
assign kdb = ~KDB;  //complement 
assign KDJ =  WHJ & ZZI & TFD  |  VDJ & ZZI & TGD  ; 
assign kdj = ~KDJ;  //complement 
assign JBC =  QPB & PBA & PBB  ; 
assign jbc = ~JBC;  //complement 
assign JBA =  ZZI & QPB  ; 
assign jba = ~JBA;  //complement 
assign JBB =  PBA & QPB  ; 
assign jbb = ~JBB;  //complement 
assign pba = ~PBA;  //complement 
assign pbd = ~PBD;  //complement 
assign pbg = ~PBG;  //complement 
assign pbb = ~PBB;  //complement 
assign pbe = ~PBE;  //complement 
assign pbh = ~PBH;  //complement 
assign pbc = ~PBC;  //complement 
assign pbf = ~PBF;  //complement 
assign pbi = ~PBI;  //complement 
assign uia = ~UIA;  //complement 
assign uib = ~UIB;  //complement 
assign uic = ~UIC;  //complement 
assign uid = ~UID;  //complement 
assign uie = ~UIE;  //complement 
assign uif = ~UIF;  //complement 
assign GIA = uif & uie ; 
assign gia = ~GIA ; //complement 
assign GIB = uif & UIE ; 
assign gib = ~GIB ;  //complement 
assign GIC = UIF & uie ; 
assign gic = ~GIC ;  //complement 
assign GID = UIF & UIE; 
assign gid = ~GID; 
assign UJD = ~ujd;  //complement 
assign UJE = ~uje;  //complement 
assign UJF = ~ujf;  //complement 
assign UJA = ~uja;  //complement 
assign UJB = ~ujb;  //complement 
assign UJC = ~ujc;  //complement 
assign GJA = ujf & uje ; 
assign gja = ~GJA ; //complement 
assign GJB = ujf & UJE ; 
assign gjb = ~GJB ;  //complement 
assign GJC = UJF & uje ; 
assign gjc = ~GJC ;  //complement 
assign GJD = UJF & UJE; 
assign gjd = ~GJD; 
assign uka = ~UKA;  //complement 
assign ukb = ~UKB;  //complement 
assign ukc = ~UKC;  //complement 
assign GKA = ukf & uke ; 
assign gka = ~GKA ; //complement 
assign GKB = ukf & UKE ; 
assign gkb = ~GKB ;  //complement 
assign GKC = UKF & uke ; 
assign gkc = ~GKC ;  //complement 
assign GKD = UKF & UKE; 
assign gkd = ~GKD; 
assign ukd = ~UKD;  //complement 
assign uke = ~UKE;  //complement 
assign ukf = ~UKF;  //complement 
assign ULD = ~uld;  //complement 
assign ULE = ~ule;  //complement 
assign ULF = ~ulf;  //complement 
assign GLA = ulf & ule ; 
assign gla = ~GLA ; //complement 
assign GLB = ulf & ULE ; 
assign glb = ~GLB ;  //complement 
assign GLC = ULF & ule ; 
assign glc = ~GLC ;  //complement 
assign GLD = ULF & ULE; 
assign gld = ~GLD; 
assign ULA = ~ula;  //complement 
assign ULB = ~ulb;  //complement 
assign ULC = ~ulc;  //complement 
assign vac = ~VAC;  //complement 
assign oac = ~OAC;  //complement 
assign wac = ~WAC;  //complement 
assign wec = ~WEC;  //complement 
assign wic = ~WIC;  //complement 
assign wmc = ~WMC;  //complement 
assign vak = ~VAK;  //complement 
assign oak = ~OAK;  //complement 
assign wak = ~WAK;  //complement 
assign wek = ~WEK;  //complement 
assign wik = ~WIK;  //complement 
assign wmk = ~WMK;  //complement 
assign vbc = ~VBC;  //complement 
assign obc = ~OBC;  //complement 
assign wbc = ~WBC;  //complement 
assign wfc = ~WFC;  //complement 
assign wjc = ~WJC;  //complement 
assign wnc = ~WNC;  //complement 
assign vbk = ~VBK;  //complement 
assign obk = ~OBK;  //complement 
assign wbk = ~WBK;  //complement 
assign wfk = ~WFK;  //complement 
assign wjk = ~WJK;  //complement 
assign wnk = ~WNK;  //complement 
assign vcc = ~VCC;  //complement 
assign occ = ~OCC;  //complement 
assign wcc = ~WCC;  //complement 
assign wgc = ~WGC;  //complement 
assign wkc = ~WKC;  //complement 
assign woc = ~WOC;  //complement 
assign vck = ~VCK;  //complement 
assign ock = ~OCK;  //complement 
assign wck = ~WCK;  //complement 
assign wgk = ~WGK;  //complement 
assign wkk = ~WKK;  //complement 
assign wok = ~WOK;  //complement 
assign vdc = ~VDC;  //complement 
assign odc = ~ODC;  //complement 
assign wdc = ~WDC;  //complement 
assign whc = ~WHC;  //complement 
assign wlc = ~WLC;  //complement 
assign wpc = ~WPC;  //complement 
assign vdk = ~VDK;  //complement 
assign odk = ~ODK;  //complement 
assign wdk = ~WDK;  //complement 
assign whk = ~WHK;  //complement 
assign wlk = ~WLK;  //complement 
assign wpk = ~WPK;  //complement 
assign KAC =  WEC & ZZI & TFA  |  VAC & ZZI & TGA  ; 
assign kac = ~KAC;  //complement 
assign KAK =  WEK & ZZI & TFA  |  VAK & ZZI & TGA  ; 
assign kak = ~KAK;  //complement 
assign qqa = ~QQA;  //complement 
assign qqe = ~QQE;  //complement 
assign qqb = ~QQB;  //complement 
assign qqf = ~QQF;  //complement 
assign tac = ~TAC;  //complement 
assign tbc = ~TBC;  //complement 
assign tcc = ~TCC;  //complement 
assign tdc = ~TDC;  //complement 
assign qqi = ~QQI;  //complement 
assign qqj = ~QQJ;  //complement 
assign KBC =  WFC & ZZI & TFB  |  VBC & ZZI & TGB  ; 
assign kbc = ~KBC;  //complement 
assign KBK =  WFK & ZZI & TFB  |  VBK & ZZI & TGB  ; 
assign kbk = ~KBK;  //complement 
assign qqk = ~QQK;  //complement 
assign JJJ =  QJH & qjm & QJK  |  QJI & qjm & QJK  ; 
assign jjj = ~JJJ;  //complement 
assign uig = ~UIG;  //complement 
assign uih = ~UIH;  //complement 
assign ulg = ~ULG;  //complement 
assign ulh = ~ULH;  //complement 
assign qjh = ~QJH;  //complement 
assign okb = ~OKB;  //complement 
assign qji = ~QJI;  //complement 
assign okc = ~OKC;  //complement 
assign OEC = ~oec;  //complement 
assign OEK = ~oek;  //complement 
assign OFC = ~ofc;  //complement 
assign OFK = ~ofk;  //complement 
assign KCC =  WGC & ZZI & TFC  |  VCC & ZZI & TGC  ; 
assign kcc = ~KCC;  //complement 
assign KCK =  WGK & ZZI & TFC  |  VCK & ZZI & TGC  ; 
assign kck = ~KCK;  //complement 
assign QHC = ~qhc;  //complement 
assign qjk = ~QJK;  //complement 
assign OGC = ~ogc;  //complement 
assign OGK = ~ogk;  //complement 
assign OHC = ~ohc;  //complement 
assign OHK = ~ohk;  //complement 
assign ujg = ~UJG;  //complement 
assign ujh = ~UJH;  //complement 
assign ukg = ~UKG;  //complement 
assign ukh = ~UKH;  //complement 
assign jcd = qcc & qbc ; 
assign JCD = ~jcd ; //complement 
assign qbc = ~QBC;  //complement 
assign qcc = ~QCC;  //complement 
assign qck = ~QCK;  //complement 
assign qdc = ~QDC;  //complement 
assign KDC =  WHC & ZZI & TFD  |  VDC & ZZI & TGD  ; 
assign kdc = ~KDC;  //complement 
assign KDK =  WHK & ZZI & TFD  |  VDK & ZZI & TGD  ; 
assign kdk = ~KDK;  //complement 
assign qpc = ~QPC;  //complement 
assign JCC =  QPC & PCA & PCB  ; 
assign jcc = ~JCC;  //complement 
assign JCA =  ZZI & QPC  ; 
assign jca = ~JCA;  //complement 
assign JCB =  PCA & QPC  ; 
assign jcb = ~JCB;  //complement 
assign OKO = ~oko;  //complement 
assign OKP = ~okp;  //complement 
assign OKQ = ~okq;  //complement 
assign pca = ~PCA;  //complement 
assign pcd = ~PCD;  //complement 
assign pcg = ~PCG;  //complement 
assign pcb = ~PCB;  //complement 
assign pce = ~PCE;  //complement 
assign pch = ~PCH;  //complement 
assign pcc = ~PCC;  //complement 
assign pcf = ~PCF;  //complement 
assign pci = ~PCI;  //complement 
assign uma = ~UMA;  //complement 
assign umb = ~UMB;  //complement 
assign umc = ~UMC;  //complement 
assign umd = ~UMD;  //complement 
assign ume = ~UME;  //complement 
assign umf = ~UMF;  //complement 
assign GMA = umf & ume ; 
assign gma = ~GMA ; //complement 
assign GMB = umf & UME ; 
assign gmb = ~GMB ;  //complement 
assign GMC = UMF & ume ; 
assign gmc = ~GMC ;  //complement 
assign GMD = UMF & UME; 
assign gmd = ~GMD; 
assign UND = ~und;  //complement 
assign UNE = ~une;  //complement 
assign UNF = ~unf;  //complement 
assign UNA = ~una;  //complement 
assign UNB = ~unb;  //complement 
assign UNC = ~unc;  //complement 
assign GNA = unf & une ; 
assign gna = ~GNA ; //complement 
assign GNB = unf & UNE ; 
assign gnb = ~GNB ;  //complement 
assign GNC = UNF & une ; 
assign gnc = ~GNC ;  //complement 
assign GND = UNF & UNE; 
assign gnd = ~GND; 
assign uoa = ~UOA;  //complement 
assign uob = ~UOB;  //complement 
assign uoc = ~UOC;  //complement 
assign GOA = uof & uoe ; 
assign goa = ~GOA ; //complement 
assign GOB = uof & UOE ; 
assign gob = ~GOB ;  //complement 
assign GOC = UOF & uoe ; 
assign goc = ~GOC ;  //complement 
assign GOD = UOF & UOE; 
assign god = ~GOD; 
assign uod = ~UOD;  //complement 
assign uoe = ~UOE;  //complement 
assign uof = ~UOF;  //complement 
assign UPD = ~upd;  //complement 
assign UPE = ~upe;  //complement 
assign UPF = ~upf;  //complement 
assign GPA = upf & upe ; 
assign gpa = ~GPA ; //complement 
assign GPB = upf & UPE ; 
assign gpb = ~GPB ;  //complement 
assign GPC = UPF & upe ; 
assign gpc = ~GPC ;  //complement 
assign GPD = UPF & UPE; 
assign gpd = ~GPD; 
assign UPA = ~upa;  //complement 
assign UPB = ~upb;  //complement 
assign UPC = ~upc;  //complement 
assign vad = ~VAD;  //complement 
assign oad = ~OAD;  //complement 
assign wad = ~WAD;  //complement 
assign wed = ~WED;  //complement 
assign wid = ~WID;  //complement 
assign wmd = ~WMD;  //complement 
assign val = ~VAL;  //complement 
assign oal = ~OAL;  //complement 
assign wal = ~WAL;  //complement 
assign wel = ~WEL;  //complement 
assign wil = ~WIL;  //complement 
assign wml = ~WML;  //complement 
assign vbd = ~VBD;  //complement 
assign obd = ~OBD;  //complement 
assign wbd = ~WBD;  //complement 
assign wfd = ~WFD;  //complement 
assign wjd = ~WJD;  //complement 
assign wnd = ~WND;  //complement 
assign vbl = ~VBL;  //complement 
assign obl = ~OBL;  //complement 
assign wbl = ~WBL;  //complement 
assign wfl = ~WFL;  //complement 
assign wjl = ~WJL;  //complement 
assign wnl = ~WNL;  //complement 
assign vcd = ~VCD;  //complement 
assign ocd = ~OCD;  //complement 
assign wcd = ~WCD;  //complement 
assign wgd = ~WGD;  //complement 
assign wkd = ~WKD;  //complement 
assign wod = ~WOD;  //complement 
assign vcl = ~VCL;  //complement 
assign ocl = ~OCL;  //complement 
assign wcl = ~WCL;  //complement 
assign wgl = ~WGL;  //complement 
assign wkl = ~WKL;  //complement 
assign wol = ~WOL;  //complement 
assign vdd = ~VDD;  //complement 
assign odd = ~ODD;  //complement 
assign wdd = ~WDD;  //complement 
assign whd = ~WHD;  //complement 
assign wld = ~WLD;  //complement 
assign wpd = ~WPD;  //complement 
assign vdl = ~VDL;  //complement 
assign odl = ~ODL;  //complement 
assign wdl = ~WDL;  //complement 
assign whl = ~WHL;  //complement 
assign wll = ~WLL;  //complement 
assign wpl = ~WPL;  //complement 
assign KAD =  WED & ZZI & TFA  |  VAD & ZZI & TGA  ; 
assign kad = ~KAD;  //complement 
assign KAL =  WEL & ZZI & TFA  |  VAL & ZZI & TGA  ; 
assign kal = ~KAL;  //complement 
assign tea = ~TEA;  //complement 
assign teb = ~TEB;  //complement 
assign tec = ~TEC;  //complement 
assign ted = ~TED;  //complement 
assign qqc = ~QQC;  //complement 
assign qqg = ~QQG;  //complement 
assign qqd = ~QQD;  //complement 
assign qqh = ~QQH;  //complement 
assign tad = ~TAD;  //complement 
assign tbd = ~TBD;  //complement 
assign tcd = ~TCD;  //complement 
assign tdd = ~TDD;  //complement 
assign JJH =  ECA & ECB & EEC  |  QJA  ; 
assign jjh = ~JJH; //complement 
assign JJI =  ECA & ECB & EEC  |  QJA  ; 
assign jji = ~JJI;  //complement 
assign qql = ~QQL;  //complement 
assign qqm = ~QQM;  //complement 
assign KBD =  WFD & ZZI & TFB  |  VBD & ZZI & TGB  ; 
assign kbd = ~KBD;  //complement 
assign KBL =  WFL & ZZI & TFB  |  VBL & ZZI & TGB  ; 
assign kbl = ~KBL;  //complement 
assign JJS = efb & efa ; 
assign jjs = ~JJS ; //complement 
assign JJT = efb & EFA ; 
assign jjt = ~JJT ;  //complement 
assign JJU = EFB & efa ; 
assign jju = ~JJU ;  //complement 
assign JJV = EFB & EFA; 
assign jjv = ~JJV; 
assign qqn = ~QQN;  //complement 
assign qqo = ~QQO;  //complement 
assign umg = ~UMG;  //complement 
assign umh = ~UMH;  //complement 
assign upg = ~UPG;  //complement 
assign uph = ~UPH;  //complement 
assign JJW = efb & efa ; 
assign jjw = ~JJW ; //complement 
assign JJX = efb & EFA ; 
assign jjx = ~JJX ;  //complement 
assign JJY = EFB & efa ; 
assign jjy = ~JJY ;  //complement 
assign JJZ = EFB & EFA; 
assign jjz = ~JJZ; 
assign efa = ~EFA;  //complement 
assign efb = ~EFB;  //complement 
assign OED = ~oed;  //complement 
assign OEL = ~oel;  //complement 
assign OFD = ~ofd;  //complement 
assign OFL = ~ofl;  //complement 
assign KCD =  WGD & ZZI & TFC  |  VCD & ZZI & TGC  ; 
assign kcd = ~KCD;  //complement 
assign KCL =  WGL & ZZI & TFC  |  VCL & ZZI & TGC  ; 
assign kcl = ~KCL;  //complement 
assign QHD = ~qhd;  //complement 
assign qeb = ~QEB;  //complement 
assign qef = ~QEF;  //complement 
assign OGD = ~ogd;  //complement 
assign OGL = ~ogl;  //complement 
assign OHD = ~ohd;  //complement 
assign OHL = ~ohl;  //complement 
assign ung = ~UNG;  //complement 
assign unh = ~UNH;  //complement 
assign uog = ~UOG;  //complement 
assign uoh = ~UOH;  //complement 
assign jdd = qcd & qbd ; 
assign JDD = ~jdd ; //complement 
assign qbd = ~QBD;  //complement 
assign qcd = ~QCD;  //complement 
assign qcl = ~QCL;  //complement 
assign qdd = ~QDD;  //complement 
assign KDD =  WHD & ZZI & TFD  |  VDD & ZZI & TGD  ; 
assign kdd = ~KDD;  //complement 
assign KDL =  WHL & ZZI & TFD  |  VDL & ZZI & TGD  ; 
assign kdl = ~KDL;  //complement 
assign qka = ~QKA;  //complement 
assign qkb = ~QKB;  //complement 
assign JDC =  QPD & PDA & PDB  ; 
assign jdc = ~JDC;  //complement 
assign JDA =  ZZI & QPD  ; 
assign jda = ~JDA;  //complement 
assign JDB =  PDA & QPD  ; 
assign jdb = ~JDB;  //complement 
assign OKR = ~okr;  //complement 
assign OKS = ~oks;  //complement 
assign okt = ~OKT;  //complement 
assign qpd = ~QPD;  //complement 
assign pda = ~PDA;  //complement 
assign pdd = ~PDD;  //complement 
assign pdg = ~PDG;  //complement 
assign pdb = ~PDB;  //complement 
assign pde = ~PDE;  //complement 
assign pdh = ~PDH;  //complement 
assign pdc = ~PDC;  //complement 
assign pdf = ~PDF;  //complement 
assign pdi = ~PDI;  //complement 
assign uai = ~UAI;  //complement 
assign uaj = ~UAJ;  //complement 
assign uak = ~UAK;  //complement 
assign ual = ~UAL;  //complement 
assign uam = ~UAM;  //complement 
assign uan = ~UAN;  //complement 
assign GAE = uan & uam ; 
assign gae = ~GAE ; //complement 
assign GAF = uan & UAM ; 
assign gaf = ~GAF ;  //complement 
assign GAG = UAN & uam ; 
assign gag = ~GAG ;  //complement 
assign GAH = UAN & UAM; 
assign gah = ~GAH; 
assign UBL = ~ubl;  //complement 
assign UBM = ~ubm;  //complement 
assign UBN = ~ubn;  //complement 
assign UBI = ~ubi;  //complement 
assign UBJ = ~ubj;  //complement 
assign UBK = ~ubk;  //complement 
assign GBE = ubn & ubm ; 
assign gbe = ~GBE ; //complement 
assign GBF = ubn & UBM ; 
assign gbf = ~GBF ;  //complement 
assign GBG = UBN & ubm ; 
assign gbg = ~GBG ;  //complement 
assign GBH = UBN & UBM; 
assign gbh = ~GBH; 
assign uci = ~UCI;  //complement 
assign ucj = ~UCJ;  //complement 
assign uck = ~UCK;  //complement 
assign GCE = ucn & ucm ; 
assign gce = ~GCE ; //complement 
assign GCF = ucn & UCM ; 
assign gcf = ~GCF ;  //complement 
assign GCG = UCN & ucm ; 
assign gcg = ~GCG ;  //complement 
assign GCH = UCN & UCM; 
assign gch = ~GCH; 
assign ucl = ~UCL;  //complement 
assign ucm = ~UCM;  //complement 
assign ucn = ~UCN;  //complement 
assign UDL = ~udl;  //complement 
assign UDM = ~udm;  //complement 
assign UDN = ~udn;  //complement 
assign GDE = udn & udm ; 
assign gde = ~GDE ; //complement 
assign GDF = udn & UDM ; 
assign gdf = ~GDF ;  //complement 
assign GDG = UDN & udm ; 
assign gdg = ~GDG ;  //complement 
assign GDH = UDN & UDM; 
assign gdh = ~GDH; 
assign UDI = ~udi;  //complement 
assign UDJ = ~udj;  //complement 
assign UDK = ~udk;  //complement 
assign vae = ~VAE;  //complement 
assign oae = ~OAE;  //complement 
assign wae = ~WAE;  //complement 
assign wee = ~WEE;  //complement 
assign wie = ~WIE;  //complement 
assign wme = ~WME;  //complement 
assign vam = ~VAM;  //complement 
assign oam = ~OAM;  //complement 
assign wam = ~WAM;  //complement 
assign wem = ~WEM;  //complement 
assign wim = ~WIM;  //complement 
assign wmm = ~WMM;  //complement 
assign vbe = ~VBE;  //complement 
assign obe = ~OBE;  //complement 
assign wbe = ~WBE;  //complement 
assign wfe = ~WFE;  //complement 
assign wje = ~WJE;  //complement 
assign wne = ~WNE;  //complement 
assign vbm = ~VBM;  //complement 
assign obm = ~OBM;  //complement 
assign wbm = ~WBM;  //complement 
assign wfm = ~WFM;  //complement 
assign wjm = ~WJM;  //complement 
assign wnm = ~WNM;  //complement 
assign vce = ~VCE;  //complement 
assign oce = ~OCE;  //complement 
assign wce = ~WCE;  //complement 
assign wge = ~WGE;  //complement 
assign wke = ~WKE;  //complement 
assign woe = ~WOE;  //complement 
assign vcm = ~VCM;  //complement 
assign ocm = ~OCM;  //complement 
assign wcm = ~WCM;  //complement 
assign wgm = ~WGM;  //complement 
assign wkm = ~WKM;  //complement 
assign wom = ~WOM;  //complement 
assign vde = ~VDE;  //complement 
assign ode = ~ODE;  //complement 
assign wde = ~WDE;  //complement 
assign whe = ~WHE;  //complement 
assign wle = ~WLE;  //complement 
assign wpe = ~WPE;  //complement 
assign vdm = ~VDM;  //complement 
assign odm = ~ODM;  //complement 
assign wdm = ~WDM;  //complement 
assign whm = ~WHM;  //complement 
assign wlm = ~WLM;  //complement 
assign wpm = ~WPM;  //complement 
assign KAE =  WEE & ZZI & TFE  |  VAE & ZZI & TGE  ; 
assign kae = ~KAE;  //complement 
assign KAM =  WEM & ZZI & TFE  |  VAM & ZZI & TGE  ; 
assign kam = ~KAM;  //complement 
assign daa = ~DAA;  //complement 
assign daf = ~DAF;  //complement 
assign dak = ~DAK;  //complement 
assign dab = ~DAB;  //complement 
assign dag = ~DAG;  //complement 
assign dal = ~DAL;  //complement 
assign dam = ~DAM;  //complement 
assign dah = ~DAH;  //complement 
assign dac = ~DAC;  //complement 
assign tae = ~TAE;  //complement 
assign tbe = ~TBE;  //complement 
assign tce = ~TCE;  //complement 
assign tde = ~TDE;  //complement 
assign JEE =  qla & DAA & DAB & DAC & DAD  ; 
assign jee = ~JEE;  //complement  
assign JEC =  qla & DAA & DAB  ; 
assign jec = ~JEC;  //complement 
assign jha = dac; 
assign JHA = ~jha; //complement 
assign jhb = dad; 
assign JHB = ~jhb;  //complement 
assign JEA = qla & ZZI ; 
assign jea = ~JEA ;  //complement 
assign JEB = qla & DAA; 
assign jeb = ~JEB; 
assign dan = ~DAN;  //complement 
assign dai = ~DAI;  //complement 
assign dad = ~DAD;  //complement 
assign KBE =  WFE & ZZI & TFF  |  VBE & ZZI & TGF  ; 
assign kbe = ~KBE;  //complement 
assign KBM =  WFM & ZZI & TFF  |  VBM & ZZI & TGF  ; 
assign kbm = ~KBM;  //complement 
assign JNA = dag & daf ; 
assign jna = ~JNA ; //complement 
assign JNB = dag & DAK ; 
assign jnb = ~JNB ;  //complement 
assign JNC = DAG & daf ; 
assign jnc = ~JNC ;  //complement 
assign JND = DAG & DAK; 
assign jnd = ~JND; 
assign JEF =  DAA & DAB & DAC & DAD & DAE  ; 
assign jef = ~JEF;  //complement  
assign JED =  qla & DAA & DAB & DAC  ; 
assign jed = ~JED;  //complement 
assign dao = ~DAO;  //complement 
assign daj = ~DAJ;  //complement 
assign dae = ~DAE;  //complement 
assign uao = ~UAO;  //complement 
assign uap = ~UAP;  //complement 
assign udo = ~UDO;  //complement 
assign udp = ~UDP;  //complement 
assign JIA =  dag & daf & QJM  ; 
assign jia = ~JIA;  //complement 
assign JIB =  dag & DAF & QJM  ; 
assign jib = ~JIB;  //complement 
assign JIC =  DAG & daf & QJM  ; 
assign jic = ~JIC;  //complement 
assign JID =  DAG & DAF & QJM  ; 
assign jid = ~JID;  //complement 
assign eaa = ~EAA;  //complement 
assign KCE =  WGE & ZZI & TFG  |  VCE & ZZI & TGG  ; 
assign kce = ~KCE;  //complement 
assign KCM =  WGM & ZZI & TFG  |  VCM & ZZI & TGG  ; 
assign kcm = ~KCM;  //complement 
assign eab = ~EAB;  //complement 
assign eac = ~EAC;  //complement 
assign OEE = ~oee;  //complement 
assign OEM = ~oem;  //complement 
assign OFE = ~ofe;  //complement 
assign OFM = ~ofm;  //complement 
assign ubo = ~UBO;  //complement 
assign ubp = ~UBP;  //complement 
assign uco = ~UCO;  //complement 
assign ucp = ~UCP;  //complement 
assign eae = ~EAE;  //complement 
assign ead = ~EAD;  //complement 
assign OGE = ~oge;  //complement 
assign OGM = ~ogm;  //complement 
assign OHE = ~ohe;  //complement 
assign OHM = ~ohm;  //complement 
assign KDE =  WHE & ZZI & TFH  |  VDE & ZZI & TGH  ; 
assign kde = ~KDE;  //complement 
assign KDM =  WHM & ZZI & TFH  |  VDM & ZZI & TGH  ; 
assign kdm = ~KDM;  //complement 
assign jma = dag & dak ; 
assign JMA = ~jma ; //complement 
assign jmb = dag & ZZI ; 
assign JMB = ~jmb ;  //complement 
assign JMC = DAK & DAG ; 
assign jmc = ~JMC ;  //complement 
assign jhc = dae; 
assign JHC = ~jhc;  //complement 
assign QLD = ~qld;  //complement 
assign JFB =  ZZO  |  ZZO  |  QLD & qjc & qju  ; 
assign jfb = ~JFB; //complement 
assign JFC =  ZZO  |  ZZO  |  QLD & qjc & qju  ; 
assign jfc = ~JFC;  //complement 
assign uei = ~UEI;  //complement 
assign uej = ~UEJ;  //complement 
assign uek = ~UEK;  //complement 
assign uel = ~UEL;  //complement 
assign uem = ~UEM;  //complement 
assign uen = ~UEN;  //complement 
assign GEE = uen & uem ; 
assign gee = ~GEE ; //complement 
assign GEF = uen & UEM ; 
assign gef = ~GEF ;  //complement 
assign GEG = UEN & uem ; 
assign geg = ~GEG ;  //complement 
assign GEH = UEN & UEM; 
assign geh = ~GEH; 
assign UFL = ~ufl;  //complement 
assign UFM = ~ufm;  //complement 
assign UFN = ~ufn;  //complement 
assign UFI = ~ufi;  //complement 
assign UFJ = ~ufj;  //complement 
assign UFK = ~ufk;  //complement 
assign GFE = ufn & ufm ; 
assign gfe = ~GFE ; //complement 
assign GFF = ufn & UFM ; 
assign gff = ~GFF ;  //complement 
assign GFG = UFN & ufm ; 
assign gfg = ~GFG ;  //complement 
assign GFH = UFN & UFM; 
assign gfh = ~GFH; 
assign ugi = ~UGI;  //complement 
assign ugj = ~UGJ;  //complement 
assign ugk = ~UGK;  //complement 
assign GGE = ugn & ugm ; 
assign gge = ~GGE ; //complement 
assign GGF = ugn & UGM ; 
assign ggf = ~GGF ;  //complement 
assign GGG = UGN & ugm ; 
assign ggg = ~GGG ;  //complement 
assign GGH = UGN & UGM; 
assign ggh = ~GGH; 
assign ugl = ~UGL;  //complement 
assign ugm = ~UGM;  //complement 
assign ugn = ~UGN;  //complement 
assign UHL = ~uhl;  //complement 
assign UHM = ~uhm;  //complement 
assign UHN = ~uhn;  //complement 
assign GHE = uhn & uhm ; 
assign ghe = ~GHE ; //complement 
assign GHF = uhn & UHM ; 
assign ghf = ~GHF ;  //complement 
assign GHG = UHN & uhm ; 
assign ghg = ~GHG ;  //complement 
assign GHH = UHN & UHM; 
assign ghh = ~GHH; 
assign UHI = ~uhi;  //complement 
assign UHJ = ~uhj;  //complement 
assign UHK = ~uhk;  //complement 
assign vaf = ~VAF;  //complement 
assign oaf = ~OAF;  //complement 
assign waf = ~WAF;  //complement 
assign wef = ~WEF;  //complement 
assign wif = ~WIF;  //complement 
assign wmf = ~WMF;  //complement 
assign van = ~VAN;  //complement 
assign oan = ~OAN;  //complement 
assign wan = ~WAN;  //complement 
assign wen = ~WEN;  //complement 
assign win = ~WIN;  //complement 
assign wmn = ~WMN;  //complement 
assign vbf = ~VBF;  //complement 
assign obf = ~OBF;  //complement 
assign wbf = ~WBF;  //complement 
assign wff = ~WFF;  //complement 
assign wjf = ~WJF;  //complement 
assign wnf = ~WNF;  //complement 
assign vbn = ~VBN;  //complement 
assign obn = ~OBN;  //complement 
assign wbn = ~WBN;  //complement 
assign wfn = ~WFN;  //complement 
assign wjn = ~WJN;  //complement 
assign wnn = ~WNN;  //complement 
assign vcf = ~VCF;  //complement 
assign ocf = ~OCF;  //complement 
assign wcf = ~WCF;  //complement 
assign wgf = ~WGF;  //complement 
assign wkf = ~WKF;  //complement 
assign wof = ~WOF;  //complement 
assign vcn = ~VCN;  //complement 
assign ocn = ~OCN;  //complement 
assign wcn = ~WCN;  //complement 
assign wgn = ~WGN;  //complement 
assign wkn = ~WKN;  //complement 
assign won = ~WON;  //complement 
assign vdf = ~VDF;  //complement 
assign odf = ~ODF;  //complement 
assign wdf = ~WDF;  //complement 
assign whf = ~WHF;  //complement 
assign wlf = ~WLF;  //complement 
assign wpf = ~WPF;  //complement 
assign vdn = ~VDN;  //complement 
assign odn = ~ODN;  //complement 
assign wdn = ~WDN;  //complement 
assign whn = ~WHN;  //complement 
assign wln = ~WLN;  //complement 
assign wpn = ~WPN;  //complement 
assign KAF =  WEF & ZZI & TFE  |  VAF & ZZI & TGE  ; 
assign kaf = ~KAF;  //complement 
assign KAN =  WEN & ZZI & TFE  |  VAN & ZZI & TGE  ; 
assign kan = ~KAN;  //complement 
assign OKI = ~oki;  //complement 
assign taf = ~TAF;  //complement 
assign tbf = ~TBF;  //complement 
assign tcf = ~TCF;  //complement 
assign tdf = ~TDF;  //complement 
assign dba = ~DBA;  //complement 
assign dbe = ~DBE;  //complement 
assign dbb = ~DBB;  //complement 
assign dbf = ~DBF;  //complement 
assign dbc = ~DBC;  //complement 
assign dbg = ~DBG;  //complement 
assign KBF =  WFF & ZZI & TFF  |  VBF & ZZI & TGF  ; 
assign kbf = ~KBF;  //complement 
assign KBN =  WFN & ZZI & TFF  |  VBN & ZZI & TGF  ; 
assign kbn = ~KBN;  //complement 
assign dbi = ~DBI;  //complement 
assign dbm = ~DBM;  //complement 
assign dbj = ~DBJ;  //complement 
assign dbn = ~DBN;  //complement 
assign dbk = ~DBK;  //complement 
assign dbo = ~DBO;  //complement 
assign ueo = ~UEO;  //complement 
assign uep = ~UEP;  //complement 
assign uho = ~UHO;  //complement 
assign uhp = ~UHP;  //complement 
assign qjd = ~QJD;  //complement 
assign okh = ~OKH;  //complement 
assign QEC = ~qec;  //complement 
assign QED = ~qed;  //complement 
assign QEE = ~qee;  //complement 
assign OEF = ~oef;  //complement 
assign OEN = ~oen;  //complement 
assign OFF = ~off;  //complement 
assign OFN = ~ofn;  //complement 
assign KCF =  WGF & ZZI & TFG  |  VCF & ZZI & TGG  ; 
assign kcf = ~KCF;  //complement 
assign KCN =  WGN & ZZI & TFG  |  VCN & ZZI & TGG  ; 
assign kcn = ~KCN;  //complement 
assign qjp = ~QJP;  //complement 
assign qjf = ~QJF;  //complement 
assign OGF = ~ogf;  //complement 
assign OGN = ~ogn;  //complement 
assign OHF = ~ohf;  //complement 
assign OHN = ~ohn;  //complement 
assign ufo = ~UFO;  //complement 
assign ufp = ~UFP;  //complement 
assign ugo = ~UGO;  //complement 
assign ugp = ~UGP;  //complement 
assign qjm = ~QJM;  //complement 
assign qjn = ~QJN;  //complement 
assign oka = ~OKA;  //complement 
assign qjc = ~QJC;  //complement 
assign qjt = ~QJT;  //complement 
assign qje = ~QJE;  //complement 
assign qjg = ~QJG;  //complement 
assign KDF =  WHF & ZZI & TFH  |  VDF & ZZI & TGH  ; 
assign kdf = ~KDF;  //complement 
assign KDN =  WHN & ZZI & TFH  |  VDN & ZZI & TGH  ; 
assign kdn = ~KDN;  //complement 
assign jpg = qjy & qlf ; 
assign JPG = ~jpg ; //complement 
assign jlx = tjd; 
assign JLX = ~jlx;  //complement 
assign jfa = qlg & qjt ; 
assign JFA = ~jfa ;  //complement 
assign jpe = qed & qeb ; 
assign JPE = ~jpe ;  //complement 
assign jpf = qed & qeb; 
assign JPF = ~jpf; 
assign qjo = ~QJO;  //complement 
assign qjl = ~QJL;  //complement 
assign tja = ~TJA;  //complement 
assign tjb = ~TJB;  //complement 
assign tjc = ~TJC;  //complement 
assign tjd = ~TJD;  //complement 
assign qlf = ~QLF;  //complement 
assign qlg = ~QLG;  //complement 
assign uii = ~UII;  //complement 
assign uij = ~UIJ;  //complement 
assign uik = ~UIK;  //complement 
assign uil = ~UIL;  //complement 
assign uim = ~UIM;  //complement 
assign uin = ~UIN;  //complement 
assign GIE = uin & uim ; 
assign gie = ~GIE ; //complement 
assign GIF = uin & UIM ; 
assign gif = ~GIF ;  //complement 
assign GIG = UIN & uim ; 
assign gig = ~GIG ;  //complement 
assign GIH = UIN & UIM; 
assign gih = ~GIH; 
assign UJL = ~ujl;  //complement 
assign UJM = ~ujm;  //complement 
assign UJN = ~ujn;  //complement 
assign UJI = ~uji;  //complement 
assign UJJ = ~ujj;  //complement 
assign UJK = ~ujk;  //complement 
assign GJE = ujn & ujm ; 
assign gje = ~GJE ; //complement 
assign GJF = ujn & UJM ; 
assign gjf = ~GJF ;  //complement 
assign GJG = UJN & ujm ; 
assign gjg = ~GJG ;  //complement 
assign GJH = UJN & UJM; 
assign gjh = ~GJH; 
assign uki = ~UKI;  //complement 
assign ukj = ~UKJ;  //complement 
assign ukk = ~UKK;  //complement 
assign GKE = ukn & ukm ; 
assign gke = ~GKE ; //complement 
assign GKF = ukn & UKM ; 
assign gkf = ~GKF ;  //complement 
assign GKG = UKN & ukm ; 
assign gkg = ~GKG ;  //complement 
assign GKH = UKN & UKM; 
assign gkh = ~GKH; 
assign ukl = ~UKL;  //complement 
assign ukm = ~UKM;  //complement 
assign ukn = ~UKN;  //complement 
assign ULL = ~ull;  //complement 
assign ULM = ~ulm;  //complement 
assign ULN = ~uln;  //complement 
assign GLE = uln & ulm ; 
assign gle = ~GLE ; //complement 
assign GLF = uln & ULM ; 
assign glf = ~GLF ;  //complement 
assign GLG = ULN & ulm ; 
assign glg = ~GLG ;  //complement 
assign GLH = ULN & ULM; 
assign glh = ~GLH; 
assign ULI = ~uli;  //complement 
assign ULJ = ~ulj;  //complement 
assign ULK = ~ulk;  //complement 
assign vag = ~VAG;  //complement 
assign oag = ~OAG;  //complement 
assign wag = ~WAG;  //complement 
assign weg = ~WEG;  //complement 
assign wig = ~WIG;  //complement 
assign wmg = ~WMG;  //complement 
assign vao = ~VAO;  //complement 
assign oao = ~OAO;  //complement 
assign wao = ~WAO;  //complement 
assign weo = ~WEO;  //complement 
assign wio = ~WIO;  //complement 
assign wmo = ~WMO;  //complement 
assign vbg = ~VBG;  //complement 
assign obg = ~OBG;  //complement 
assign wbg = ~WBG;  //complement 
assign wfg = ~WFG;  //complement 
assign wjg = ~WJG;  //complement 
assign wng = ~WNG;  //complement 
assign vbo = ~VBO;  //complement 
assign obo = ~OBO;  //complement 
assign wbo = ~WBO;  //complement 
assign wfo = ~WFO;  //complement 
assign wjo = ~WJO;  //complement 
assign wno = ~WNO;  //complement 
assign vcg = ~VCG;  //complement 
assign ocg = ~OCG;  //complement 
assign wcg = ~WCG;  //complement 
assign wgg = ~WGG;  //complement 
assign wkg = ~WKG;  //complement 
assign wog = ~WOG;  //complement 
assign vco = ~VCO;  //complement 
assign oco = ~OCO;  //complement 
assign wco = ~WCO;  //complement 
assign wgo = ~WGO;  //complement 
assign wko = ~WKO;  //complement 
assign woo = ~WOO;  //complement 
assign vdg = ~VDG;  //complement 
assign odg = ~ODG;  //complement 
assign wdg = ~WDG;  //complement 
assign whg = ~WHG;  //complement 
assign wlg = ~WLG;  //complement 
assign wpg = ~WPG;  //complement 
assign vdo = ~VDO;  //complement 
assign odo = ~ODO;  //complement 
assign wdo = ~WDO;  //complement 
assign who = ~WHO;  //complement 
assign wlo = ~WLO;  //complement 
assign wpo = ~WPO;  //complement 
assign KAG =  WEG & ZZI & TFE  |  VAG & ZZI & TGE  ; 
assign kag = ~KAG;  //complement 
assign KAO =  WEO & ZZI & TFE  |  VAO & ZZI & TGE  ; 
assign kao = ~KAO;  //complement 
assign tee = ~TEE;  //complement 
assign tef = ~TEF;  //complement 
assign teg = ~TEG;  //complement 
assign teh = ~TEH;  //complement 
assign tag = ~TAG;  //complement 
assign tbg = ~TBG;  //complement 
assign tcg = ~TCG;  //complement 
assign tdg = ~TDG;  //complement 
assign KBG =  WFG & ZZI & TFF  |  VBG & ZZI & TGF  ; 
assign kbg = ~KBG;  //complement 
assign KBO =  WFO & ZZI & TFF  |  VBO & ZZI & TGF  ; 
assign kbo = ~KBO;  //complement 
assign jla =  ZZI & ZZI & qde  ; 
assign JLA = ~jla;  //complement 
assign jlb =  ZZI & ZZI & qde  |  faa  ; 
assign JLB = ~jlb;  //complement 
assign faa = ~FAA;  //complement 
assign fba = ~FBA;  //complement 
assign qjv = ~QJV;  //complement 
assign qjw = ~QJW;  //complement 
assign uio = ~UIO;  //complement 
assign uip = ~UIP;  //complement 
assign ulo = ~ULO;  //complement 
assign ulp = ~ULP;  //complement 
assign JLF =  QDE & FBA & FBB & FBC & FBD & FBE  ; 
assign jlf = ~JLF;  //complement  
assign JLC =  QDE & FAA & FAB  ; 
assign jlc = ~JLC;  //complement 
assign fab = ~FAB;  //complement 
assign fbb = ~FBB;  //complement 
assign OEG = ~oeg;  //complement 
assign OEO = ~oeo;  //complement 
assign OFG = ~ofg;  //complement 
assign OFO = ~ofo;  //complement 
assign KCG =  WGG & ZZI & TFG  |  VCG & ZZI & TGG  ; 
assign kcg = ~KCG;  //complement 
assign KCO =  WGO & ZZI & TFG  |  VCO & ZZI & TGG  ; 
assign kco = ~KCO;  //complement 
assign JPC =  QJF & qed & qja & qjd & qjn & qjp  ; 
assign jpc = ~JPC;  //complement  
assign JPD =  qha & qhb & qhc & qhd & qlh  ; 
assign jpd = ~JPD;  //complement  
assign OGG = ~ogg;  //complement 
assign OGO = ~ogo;  //complement 
assign OHG = ~ohg;  //complement 
assign OHO = ~oho;  //complement 
assign ujo = ~UJO;  //complement 
assign ujp = ~UJP;  //complement 
assign uko = ~UKO;  //complement 
assign ukp = ~UKP;  //complement 
assign JXA = QJJ & QEE ; 
assign jxa = ~JXA ;  //complement 
assign QJA = ~qja;  //complement 
assign qjb = ~QJB;  //complement 
assign qjr = ~QJR;  //complement 
assign QJZ = ~qjz;  //complement 
assign oja = ~OJA;  //complement 
assign okg = ~OKG;  //complement 
assign ojd = ~OJD;  //complement 
assign QJJ = ~qjj;  //complement 
assign KDG =  WHG & ZZI & TFH  |  VDG & ZZI & TGH  ; 
assign kdg = ~KDG;  //complement 
assign KDO =  WHO & ZZI & TFH  |  VDO & ZZI & TGH  ; 
assign kdo = ~KDO;  //complement 
assign pea = ~PEA;  //complement 
assign pfa = ~PFA;  //complement 
assign pga = ~PGA;  //complement 
assign qjx = ~QJX;  //complement 
assign qjy = ~QJY;  //complement 
assign ojb = ~OJB;  //complement 
assign qju = ~QJU;  //complement 
assign ojf = ~OJF;  //complement 
assign pxa = ~PXA;  //complement 
assign pxb = ~PXB;  //complement 
assign pxc = ~PXC;  //complement 
assign peb = ~PEB;  //complement 
assign pfb = ~PFB;  //complement 
assign pgb = ~PGB;  //complement 
assign pec = ~PEC;  //complement 
assign pfc = ~PFC;  //complement 
assign pgc = ~PGC;  //complement 
assign qlh = ~QLH;  //complement 
assign QLJ = ~qlj;  //complement 
assign qjq = ~QJQ;  //complement 
assign qjs = ~QJS;  //complement 
assign umi = ~UMI;  //complement 
assign umj = ~UMJ;  //complement 
assign umk = ~UMK;  //complement 
assign uml = ~UML;  //complement 
assign umm = ~UMM;  //complement 
assign umn = ~UMN;  //complement 
assign GME = umn & umm ; 
assign gme = ~GME ; //complement 
assign GMF = umn & UMM ; 
assign gmf = ~GMF ;  //complement 
assign GMG = UMN & umm ; 
assign gmg = ~GMG ;  //complement 
assign GMH = UMN & UMM; 
assign gmh = ~GMH; 
assign UNL = ~unl;  //complement 
assign UNM = ~unm;  //complement 
assign UNN = ~unn;  //complement 
assign UNI = ~uni;  //complement 
assign UNJ = ~unj;  //complement 
assign UNK = ~unk;  //complement 
assign GNE = unn & unm ; 
assign gne = ~GNE ; //complement 
assign GNF = unn & UNM ; 
assign gnf = ~GNF ;  //complement 
assign GNG = UNN & unm ; 
assign gng = ~GNG ;  //complement 
assign GNH = UNN & UNM; 
assign gnh = ~GNH; 
assign uoi = ~UOI;  //complement 
assign uoj = ~UOJ;  //complement 
assign uok = ~UOK;  //complement 
assign GOE = uon & uom ; 
assign goe = ~GOE ; //complement 
assign GOF = uon & UOM ; 
assign gof = ~GOF ;  //complement 
assign GOG = UON & uom ; 
assign gog = ~GOG ;  //complement 
assign GOH = UON & UOM; 
assign goh = ~GOH; 
assign uol = ~UOL;  //complement 
assign uom = ~UOM;  //complement 
assign uon = ~UON;  //complement 
assign UPL = ~upl;  //complement 
assign UPM = ~upm;  //complement 
assign UPN = ~upn;  //complement 
assign GPE = upn & upm ; 
assign gpe = ~GPE ; //complement 
assign GPF = upn & UPM ; 
assign gpf = ~GPF ;  //complement 
assign GPG = UPN & upm ; 
assign gpg = ~GPG ;  //complement 
assign GPH = UPN & UPM; 
assign gph = ~GPH; 
assign UPI = ~upi;  //complement 
assign UPJ = ~upj;  //complement 
assign UPK = ~upk;  //complement 
assign vah = ~VAH;  //complement 
assign oah = ~OAH;  //complement 
assign wah = ~WAH;  //complement 
assign weh = ~WEH;  //complement 
assign wih = ~WIH;  //complement 
assign wmh = ~WMH;  //complement 
assign vap = ~VAP;  //complement 
assign oap = ~OAP;  //complement 
assign wap = ~WAP;  //complement 
assign wep = ~WEP;  //complement 
assign wip = ~WIP;  //complement 
assign wmp = ~WMP;  //complement 
assign vbh = ~VBH;  //complement 
assign obh = ~OBH;  //complement 
assign wbh = ~WBH;  //complement 
assign wfh = ~WFH;  //complement 
assign wjh = ~WJH;  //complement 
assign wnh = ~WNH;  //complement 
assign vbp = ~VBP;  //complement 
assign obp = ~OBP;  //complement 
assign wbp = ~WBP;  //complement 
assign wfp = ~WFP;  //complement 
assign wjp = ~WJP;  //complement 
assign wnp = ~WNP;  //complement 
assign vch = ~VCH;  //complement 
assign och = ~OCH;  //complement 
assign wch = ~WCH;  //complement 
assign wgh = ~WGH;  //complement 
assign wkh = ~WKH;  //complement 
assign woh = ~WOH;  //complement 
assign vcp = ~VCP;  //complement 
assign ocp = ~OCP;  //complement 
assign wcp = ~WCP;  //complement 
assign wgp = ~WGP;  //complement 
assign wkp = ~WKP;  //complement 
assign wop = ~WOP;  //complement 
assign vdh = ~VDH;  //complement 
assign odh = ~ODH;  //complement 
assign wdh = ~WDH;  //complement 
assign whh = ~WHH;  //complement 
assign wlh = ~WLH;  //complement 
assign wph = ~WPH;  //complement 
assign vdp = ~VDP;  //complement 
assign odp = ~ODP;  //complement 
assign wdp = ~WDP;  //complement 
assign whp = ~WHP;  //complement 
assign wlp = ~WLP;  //complement 
assign wpp = ~WPP;  //complement 
assign KAH =  WEH & ZZI & TFE  |  VAH & ZZI & TGE  ; 
assign kah = ~KAH;  //complement 
assign KAP =  WEP & ZZI & TFE  |  VAP & ZZI & TGE  ; 
assign kap = ~KAP;  //complement 
assign TFA = ~tfa;  //complement 
assign TFE = ~tfe;  //complement 
assign tga = ~TGA;  //complement 
assign tge = ~TGE;  //complement 
assign tah = ~TAH;  //complement 
assign tbh = ~TBH;  //complement 
assign tch = ~TCH;  //complement 
assign tdh = ~TDH;  //complement 
assign KBH =  WFH & ZZI & TFF  |  VBH & ZZI & TGF  ; 
assign kbh = ~KBH;  //complement 
assign KBP =  WFP & ZZI & TFF  |  VBP & ZZI & TGF  ; 
assign kbp = ~KBP;  //complement 
assign TFB = ~tfb;  //complement 
assign TFF = ~tff;  //complement 
assign tgb = ~TGB;  //complement 
assign tgf = ~TGF;  //complement 
assign fac = ~FAC;  //complement 
assign fbc = ~FBC;  //complement 
assign OKU = ~oku;  //complement 
assign OKV = ~okv;  //complement 
assign umo = ~UMO;  //complement 
assign ump = ~UMP;  //complement 
assign upo = ~UPO;  //complement 
assign upp = ~UPP;  //complement 
assign JLE =  QDE & FAA & FAB & FAC & FAD  ; 
assign jle = ~JLE;  //complement  
assign JLD =  QDE & FAA & FAB & FAC  ; 
assign jld = ~JLD;  //complement 
assign fad = ~FAD;  //complement 
assign fbd = ~FBD;  //complement 
assign OEH = ~oeh;  //complement 
assign OEP = ~oep;  //complement 
assign OFH = ~ofh;  //complement 
assign OFP = ~ofp;  //complement 
assign KCH =  WGH & ZZI & TFG  |  VCH & ZZI & TGG  ; 
assign kch = ~KCH;  //complement 
assign KCP =  WGP & ZZI & TFG  |  VCP & ZZI & TGG  ; 
assign kcp = ~KCP;  //complement 
assign TFC = ~tfc;  //complement 
assign TFG = ~tfg;  //complement 
assign tgc = ~TGC;  //complement 
assign tgg = ~TGG;  //complement 
assign fae = ~FAE;  //complement 
assign fbe = ~FBE;  //complement 
assign OGH = ~ogh;  //complement 
assign OGP = ~ogp;  //complement 
assign OHH = ~ohh;  //complement 
assign OHP = ~ohp;  //complement 
assign uno = ~UNO;  //complement 
assign unp = ~UNP;  //complement 
assign uoo = ~UOO;  //complement 
assign uop = ~UOP;  //complement 
assign tma = ~TMA;  //complement 
assign jxb = qlb; 
assign JXB = ~jxb; //complement 
assign QLB = ~qlb;  //complement 
assign KDH =  WHH & ZZI & TFH  |  VDH & ZZI & TGH  ; 
assign kdh = ~KDH;  //complement 
assign KDP =  WHP & ZZI & TFH  |  VDP & ZZI & TGH  ; 
assign kdp = ~KDP;  //complement 
assign TFD = ~tfd;  //complement 
assign TFH = ~tfh;  //complement 
assign tgd = ~TGD;  //complement 
assign tgh = ~TGH;  //complement 
assign QLA = ~qla;  //complement 
assign OKW = ~okw;  //complement 
assign OKX = ~okx;  //complement 
assign EBA = ~eba;  //complement 
assign EBB = ~ebb;  //complement 
assign EBC = ~ebc;  //complement 
assign iaa = ~IAA; //complement 
assign iab = ~IAB; //complement 
assign iac = ~IAC; //complement 
assign iad = ~IAD; //complement 
assign iae = ~IAE; //complement 
assign iaf = ~IAF; //complement 
assign iag = ~IAG; //complement 
assign iah = ~IAH; //complement 
assign iai = ~IAI; //complement 
assign iaj = ~IAJ; //complement 
assign iak = ~IAK; //complement 
assign ial = ~IAL; //complement 
assign iam = ~IAM; //complement 
assign ian = ~IAN; //complement 
assign iao = ~IAO; //complement 
assign iap = ~IAP; //complement 
assign iba = ~IBA; //complement 
assign ibb = ~IBB; //complement 
assign ibc = ~IBC; //complement 
assign ibd = ~IBD; //complement 
assign ibe = ~IBE; //complement 
assign ibf = ~IBF; //complement 
assign ibg = ~IBG; //complement 
assign ibh = ~IBH; //complement 
assign ibi = ~IBI; //complement 
assign ibj = ~IBJ; //complement 
assign ibk = ~IBK; //complement 
assign ibl = ~IBL; //complement 
assign ibm = ~IBM; //complement 
assign ibn = ~IBN; //complement 
assign ibo = ~IBO; //complement 
assign ibp = ~IBP; //complement 
assign ica = ~ICA; //complement 
assign icb = ~ICB; //complement 
assign icc = ~ICC; //complement 
assign icd = ~ICD; //complement 
assign ice = ~ICE; //complement 
assign icf = ~ICF; //complement 
assign icg = ~ICG; //complement 
assign ich = ~ICH; //complement 
assign ici = ~ICI; //complement 
assign icj = ~ICJ; //complement 
assign ick = ~ICK; //complement 
assign icl = ~ICL; //complement 
assign icm = ~ICM; //complement 
assign icn = ~ICN; //complement 
assign ico = ~ICO; //complement 
assign icp = ~ICP; //complement 
assign ida = ~IDA; //complement 
assign idb = ~IDB; //complement 
assign idc = ~IDC; //complement 
assign idd = ~IDD; //complement 
assign ide = ~IDE; //complement 
assign idf = ~IDF; //complement 
assign idg = ~IDG; //complement 
assign idh = ~IDH; //complement 
assign idi = ~IDI; //complement 
assign idj = ~IDJ; //complement 
assign idk = ~IDK; //complement 
assign idl = ~IDL; //complement 
assign idm = ~IDM; //complement 
assign idn = ~IDN; //complement 
assign ido = ~IDO; //complement 
assign idp = ~IDP; //complement 
assign iea = ~IEA; //complement 
assign ieb = ~IEB; //complement 
assign iec = ~IEC; //complement 
assign ied = ~IED; //complement 
assign iee = ~IEE; //complement 
assign ief = ~IEF; //complement 
assign ieg = ~IEG; //complement 
assign ieh = ~IEH; //complement 
assign iei = ~IEI; //complement 
assign iej = ~IEJ; //complement 
assign ifa = ~IFA; //complement 
assign ifb = ~IFB; //complement 
assign ifc = ~IFC; //complement 
assign ifd = ~IFD; //complement 
assign ife = ~IFE; //complement 
assign iga = ~IGA; //complement 
assign igb = ~IGB; //complement 
assign igc = ~IGC; //complement 
assign iha = ~IHA; //complement 
assign ihb = ~IHB; //complement 
assign ija = ~IJA; //complement 
assign ijb = ~IJB; //complement 
assign ijd = ~IJD; //complement 
assign ije = ~IJE; //complement 
assign ijf = ~IJF; //complement 
assign ijg = ~IJG; //complement 
assign izz = ~IZZ; //complement 
 
assign NAA = RAA | SAA | XAA | YAA;
assign NAB = RAB | SAB | XAB | YAB;
assign NAC = RAC | SAC | XAC | YAC;
assign NAD = RAD | SAD | XAD | YAD;
assign NAE = RAE | SAE | XAE | YAE;
assign NAF = RAF | SAF | XAF | YAF;
assign NAG = RAG | SAG | XAG | YAG;
assign NAH = RAH | SAH | XAH | YAH;
assign NAI = RAI | SAI | XAI | YAI;
assign NAJ = RAJ | SAJ | XAJ | YAJ;
assign NAK = RAK | SAK | XAK | YAK;
assign NAL = RAL | SAL | XAL | YAL;
assign NAM = RAM | SAM | XAM | YAM;
assign NAN = RAN | SAN | XAN | YAN;
assign NAO = RAO | SAO | XAO | YAO;
assign NAP = RAP | SAP | XAP | YAP;
assign NBA = RBA | SBA | XBA | YBA;
assign NBB = RBB | SBB | XBB | YBB;
assign NBC = RBC | SBC | XBC | YBC;
assign NBD = RBD | SBD | XBD | YBD;
assign NBE = RBE | SBE | XBE | YBE;
assign NBF = RBF | SBF | XBF | YBF;
assign NBG = RBG | SBG | XBG | YBG;
assign NBH = RBH | SBH | XBH | YBH;
assign NBI = RBI | SBI | XBI | YBI;
assign NBJ = RBJ | SBJ | XBJ | YBJ;
assign NBK = RBK | SBK | XBK | YBK;
assign NBL = RBL | SBL | XBL | YBL;
assign NBM = RBM | SBM | XBM | YBM;
assign NBN = RBN | SBN | XBN | YBN;
assign NBO = RBO | SBO | XBO | YBO;
assign NBP = RBP | SBP | XBP | YBP;
assign NCA = RCA | SCA | XCA | YCA;
assign NCB = RCB | SCB | XCB | YCB;
assign NCC = RCC | SCC | XCC | YCC;
assign NCD = RCD | SCD | XCD | YCD;
assign NCE = RCE | SCE | XCE | YCE;
assign NCF = RCF | SCF | XCF | YCF;
assign NCG = RCG | SCG | XCG | YCG;
assign NCH = RCH | SCH | XCH | YCH;
assign NCI = RCI | SCI | XCI | YCI;
assign NCJ = RCJ | SCJ | XCJ | YCJ;
assign NCK = RCK | SCK | XCK | YCK;
assign NCL = RCL | SCL | XCL | YCL;
assign NCM = RCM | SCM | XCM | YCM;
assign NCN = RCN | SCN | XCN | YCN;
assign NCO = RCO | SCO | XCO | YCO;
assign NCP = RCP | SCP | XCP | YCP;
assign NDA = RDA | SDA | XDA | YDA;
assign NDB = RDB | SDB | XDB | YDB;
assign NDC = RDC | SDC | XDC | YDC;
assign NDD = RDD | SDD | XDD | YDD;
assign NDE = RDE | SDE | XDE | YDE;
assign NDF = RDF | SDF | XDF | YDF;
assign NDG = RDG | SDG | XDG | YDG;
assign NDH = RDH | SDH | XDH | YDH;
assign NDI = RDI | SDI | XDI | YDI;
assign NDJ = RDJ | SDJ | XDJ | YDJ;
assign NDK = RDK | SDK | XDK | YDK;
assign NDL = RDL | SDL | XDL | YDL;
assign NDM = RDM | SDM | XDM | YDM;
assign NDN = RDN | SDN | XDN | YDN;
assign NDO = RDO | SDO | XDO | YDO;
assign NDP = RDP | SDP | XDP | YDP;
assign NEA = REA | SEA | XEA | YEA;
assign NEB = REB | SEB | XEB | YEB;
assign NEC = REC | SEC | XEC | YEC;
assign NED = RED | SED | XED | YED;
assign NEE = REE | SEE | XEE | YEE;
assign NEF = REFF  | SEF | XEF | YEF;
assign NEG = REG | SEG | XEG | YEG;
assign NEH = REH | SEH | XEH | YEH;
assign NEI = REI | SEI | XEI | YEI;
assign NEJ = REJ | SEJ | XEJ | YEJ;
assign NEK = REK | SEK | XEK | YEK;
assign NEL = REL | SEL | XEL | YEL;
assign NEM = REM | SEM | XEM | YEM;
assign NEN = REN | SEN | XEN | YEN;
assign NEO = REO | SEO | XEO | YEO;
assign NEP = REP | SEP | XEP | YEP;
assign NFA = RFA | SFA | XFA | YFA;
assign NFB = RFB | SFB | XFB | YFB;
assign NFC = RFC | SFC | XFC | YFC;
assign NFD = RFD | SFD | XFD | YFD;
assign NFE = RFE | SFE | XFE | YFE;
assign NFF = RFF | SFF | XFF | YFF;
assign NFG = RFG | SFG | XFG | YFG;
assign NFH = RFH | SFH | XFH | YFH;
assign NFI = RFI | SFI | XFI | YFI;
assign NFJ = RFJ | SFJ | XFJ | YFJ;
assign NFK = RFK | SFK | XFK | YFK;
assign NFL = RFL | SFL | XFL | YFL;
assign NFM = RFM | SFM | XFM | YFM;
assign NFN = RFN | SFN | XFN | YFN;
assign NFO = RFO | SFO | XFO | YFO;
assign NFP = RFP | SFP | XFP | YFP;
assign NGA = RGA | SGA | XGA | YGA;
assign NGB = RGB | SGB | XGB | YGB;
assign NGC = RGC | SGC | XGC | YGC;
assign NGD = RGD | SGD | XGD | YGD;
assign NGE = RGE | SGE | XGE | YGE;
assign NGF = RGF | SGF | XGF | YGF;
assign NGG = RGG | SGG | XGG | YGG;
assign NGH = RGH | SGH | XGH | YGH;
assign NGI = RGI | SGI | XGI | YGI;
assign NGJ = RGJ | SGJ | XGJ | YGJ;
assign NGK = RGK | SGK | XGK | YGK;
assign NGL = RGL | SGL | XGL | YGL;
assign NGM = RGM | SGM | XGM | YGM;
assign NGN = RGN | SGN | XGN | YGN;
assign NGO = RGO | SGO | XGO | YGO;
assign NGP = RGP | SGP | XGP | YGP;
assign NHA = RHA | SHA | XHA | YHA;
assign NHB = RHB | SHB | XHB | YHB;
assign NHC = RHC | SHC | XHC | YHC;
assign NHD = RHD | SHD | XHD | YHD;
assign NHE = RHE | SHE | XHE | YHE;
assign NHF = RHF | SHF | XHF | YHF;
assign NHG = RHG | SHG | XHG | YHG;
assign NHH = RHH | SHH | XHH | YHH;
assign NHI = RHI | SHI | XHI | YHI;
assign NHJ = RHJ | SHJ | XHJ | YHJ;
assign NHK = RHK | SHK | XHK | YHK;
assign NHL = RHL | SHL | XHL | YHL;
assign NHM = RHM | SHM | XHM | YHM;
assign NHN = RHN | SHN | XHN | YHN;
assign NHO = RHO | SHO | XHO | YHO;
assign NHP = RHP | SHP | XHP | YHP;
assign NIA = RIA | SIA | XIA | YIA;
assign NIB = RIB | SIB | XIB | YIB;
assign NIC = RIC | SIC | XIC | YIC;
assign NID = RID | SID | XID | YID;
assign NIE = RIE | SIE | XIE | YIE;
assign NIF = RIF | SIF | XIF | YIF;
assign NIG = RIG | SIG | XIG | YIG;
assign NIH = RIH | SIH | XIH | YIH;
assign NII = RII | SII | XII | YII;
assign NIJ = RIJ | SIJ | XIJ | YIJ;
assign NIK = RIK | SIK | XIK | YIK;
assign NIL = RIL | SIL | XIL | YIL;
assign NIM = RIM | SIM | XIM | YIM;
assign NIN = RIN | SIN | XIN | YIN;
assign NIO = RIO | SIO | XIO | YIO;
assign NIP = RIP | SIP | XIP | YIP;
assign NJA = RJA | SJA | XJA | YJA;
assign NJB = RJB | SJB | XJB | YJB;
assign NJC = RJC | SJC | XJC | YJC;
assign NJD = RJD | SJD | XJD | YJD;
assign NJE = RJE | SJE | XJE | YJE;
assign NJF = RJF | SJF | XJF | YJF;
assign NJG = RJG | SJG | XJG | YJG;
assign NJH = RJH | SJH | XJH | YJH;
assign NJI = RJI | SJI | XJI | YJI;
assign NJJ = RJJ | SJJ | XJJ | YJJ;
assign NJK = RJK | SJK | XJK | YJK;
assign NJL = RJL | SJL | XJL | YJL;
assign NJM = RJM | SJM | XJM | YJM;
assign NJN = RJN | SJN | XJN | YJN;
assign NJO = RJO | SJO | XJO | YJO;
assign NJP = RJP | SJP | XJP | YJP;
assign NKA = RKA | SKA | XKA | YKA;
assign NKB = RKB | SKB | XKB | YKB;
assign NKC = RKC | SKC | XKC | YKC;
assign NKD = RKD | SKD | XKD | YKD;
assign NKE = RKE | SKE | XKE | YKE;
assign NKF = RKF | SKF | XKF | YKF;
assign NKG = RKG | SKG | XKG | YKG;
assign NKH = RKH | SKH | XKH | YKH;
assign NKI = RKI | SKI | XKI | YKI;
assign NKJ = RKJ | SKJ | XKJ | YKJ;
assign NKK = RKK | SKK | XKK | YKK;
assign NKL = RKL | SKL | XKL | YKL;
assign NKM = RKM | SKM | XKM | YKM;
assign NKN = RKN | SKN | XKN | YKN;
assign NKO = RKO | SKO | XKO | YKO;
assign NKP = RKP | SKP | XKP | YKP;
assign NKA = RKA | SKA | XKA | YKA;
assign NKB = RKB | SKB | XKB | YKB;
assign NKC = RKC | SKC | XKC | YKC;
assign NKD = RKD | SKD | XKD | YKD;
assign NKE = RKE | SKE | XKE | YKE;
assign NKF = RKF | SKF | XKF | YKF;
assign NKG = RKG | SKG | XKG | YKG;
assign NKH = RKH | SKH | XKH | YKH;
assign NKI = RKI | SKI | XKI | YKI;
assign NKJ = RKJ | SKJ | XKJ | YKJ;
assign NKK = RKK | SKK | XKK | YKK;
assign NKL = RKL | SKL | XKL | YKL;
assign NKM = RKM | SKM | XKM | YKM;
assign NKN = RKN | SKN | XKN | YKN;
assign NKO = RKO | SKO | XKO | YKO;
assign NKP = RKP | SKP | XKP | YKP;
assign NLA = RLA | SLA | XLA | YLA;
assign NLB = RLB | SLB | XLB | YLB;
assign NLC = RLC | SLC | XLC | YLC;
assign NLD = RLD | SLD | XLD | YLD;
assign NLE = RLE | SLE | XLE | YLE;
assign NLF = RLF | SLF | XLF | YLF;
assign NLG = RLG | SLG | XLG | YLG;
assign NLH = RLH | SLH | XLH | YLH;
assign NLI = RLI | SLI | XLI | YLI;
assign NLJ = RLJ | SLJ | XLJ | YLJ;
assign NLK = RLK | SLK | XLK | YLK;
assign NLL = RLL | SLL | XLL | YLL;
assign NLM = RLM | SLM | XLM | YLM;
assign NLN = RLN | SLN | XLN | YLN;
assign NLO = RLO | SLO | XLO | YLO;
assign NLP = RLP | SLP | XLP | YLP;
assign NMA = RMA | SMA | XMA | YMA;
assign NMB = RMB | SMB | XMB | YMB;
assign NMC = RMC | SMC | XMC | YMC;
assign NMD = RMD | SMD | XMD | YMD;
assign NME = RME | SME | XME | YME;
assign NMF = RMF | SMF | XMF | YMF;
assign NMG = RMG | SMG | XMG | YMG;
assign NMH = RMH | SMH | XMH | YMH;
assign NMI = RMI | SMI | XMI | YMI;
assign NMJ = RMJ | SMJ | XMJ | YMJ;
assign NMK = RMK | SMK | XMK | YMK;
assign NML = RML | SML | XML | YML;
assign NMM = RMM | SMM | XMM | YMM;
assign NMN = RMN | SMN | XMN | YMN;
assign NMO = RMO | SMO | XMO | YMO;
assign NMP = RMP | SMP | XMP | YMP;
assign NNA = RNA | SNA | XNA | YNA;
assign NNB = RNB | SNB | XNB | YNB;
assign NNC = RNC | SNC | XNC | YNC;
assign NND = RND | SND | XND | YND;
assign NNE = RNE | SNE | XNE | YNE;
assign NNF = RNF | SNF | XNF | YNF;
assign NNG = RNG | SNG | XNG | YNG;
assign NNH = RNH | SNH | XNH | YNH;
assign NNI = RNI | SNI | XNI | YNI;
assign NNJ = RNJ | SNJ | XNJ | YNJ;
assign NNK = RNK | SNK | XNK | YNK;
assign NNL = RNL | SNL | XNL | YNL;
assign NNM = RNM | SNM | XNM | YNM;
assign NNN = RNN | SNN | XNN | YNN;
assign NNO = RNO | SNO | XNO | YNO;
assign NNP = RNP | SNP | XNP | YNP;
assign NOA = ROA | SOA | XOA | YOA;
assign NOB = ROB | SOB | XOB | YOB;
assign NOC = ROC | SOC | XOC | YOC;
assign NOD = ROD | SOD | XOD | YOD;
assign NOE = ROE | SOE | XOE | YOE;
assign NOF = ROF | SOF | XOF | YOF;
assign NOG = ROG | SOG | XOG | YOG;
assign NOH = ROH | SOH | XOH | YOH;
assign NOI = ROI | SOI | XOI | YOI;
assign NOJ = ROJ | SOJ | XOJ | YOJ;
assign NOK = ROK | SOK | XOK | YOK;
assign NOL = ROL | SOL | XOL | YOL;
assign NOM = ROM | SOM | XOM | YOM;
assign NON = RON | SON | XON | YON;
assign NOO = ROO | SOO | XOO | YOO;
assign NOP = ROP | SOP | XOP | YOP;
assign NPA = RPA | SPA | XPA | YPA;
assign NPB = RPB | SPB | XPB | YPB;
assign NPC = RPC | SPC | XPC | YPC;
assign NPD = RPD | SPD | XPD | YPD;
assign NPE = RPE | SPE | XPE | YPE;
assign NPF = RPF | SPF | XPF | YPF;
assign NPG = RPG | SPG | XPG | YPG;
assign NPH = RPH | SPH | XPH | YPH;
assign NPI = RPI | SPI | XPI | YPI;
assign NPJ = RPJ | SPJ | XPJ | YPJ;
assign NPK = RPK | SPK | XPK | YPK;
assign NPL = RPL | SPL | XPL | YPL;
assign NPM = RPM | SPM | XPM | YPM;
assign NPN = RPN | SPN | XPN | YPN;
assign NPO = RPO | SPO | XPO | YPO;
assign NPP = RPP | SPP | XPP | YPP;

always@(posedge IZZ )
   begin 
 UAA <= PAD & TEA |  DAH & tea ; 
 UAB <= PAE & TEA |  DAI & tea ; 
 UAC <= PFA & TEA |  DBE & tea ; 
 UAD <= PFB & TEA |  DBF & tea ; 
 UAE <= PAF & TEA |  DAJ & tea ; 
 UAF <= PFC & TEA |  DBG & tea ; 
 ubd <= pfb & TEA |  dbf & tea ; 
 ube <= paf & TEA |  daj & tea ; 
 ubf <= pfc & TEA |  dbg & tea ; 
 uba <= pad & TEA |  dah & tea ; 
 ubb <= pae & TEA |  dai & tea ; 
 ubc <= pfa & TEA |  dbe & tea ; 
 UCA <= DAM & tea |  PAD & TEA ; 
 UCB <= DAN & tea |  PAE & TEA ; 
 UCC <= DBI & tea |  PGA & TEA ; 
 UCD <= DBJ & tea |  PGB & TEA ; 
 UCE <= DAO & tea |  PAF & TEA ; 
 UCF <= DBK & tea |  PGC & TEA ; 
 udd <= dbn & tea |  pgb & TEA ; 
 ude <= dao & tea |  paf & TEA ; 
 udf <= dbo & tea |  pgc & TEA ; 
 uda <= dam & tea |  pad & TEA ; 
 udb <= dan & tea |  pae & TEA ; 
 udc <= dbm & tea |  pga & TEA ; 
 VAA <=  NAA & TAA  |  NEA & TBA  |  NIA & TCA  |  NMA & TDA  |  KAA  ; 
 OAA <=  NAA & TAA  |  NEA & TBA  |  NIA & TCA  |  NMA & TDA  |  KAA  ; 
 WAA <= IAA ; 
 WEA <= IAA ; 
 WIA <= IAA ; 
 WMA <= IAA ; 
 VAI <=  NAI & TAB  |  NEI & TBB  |  NII & TCB  |  NMI & TDB  |  KAI  ; 
 OAI <=  NAI & TAB  |  NEI & TBB  |  NII & TCB  |  NMI & TDB  |  KAI  ; 
 WAI <= IAI ; 
 WEI <= IAI ; 
 WII <= IAI ; 
 WMI <= IAI ; 
 VBA <=  NBA & TAC  |  NFA & TBC  |  NJA & TCC  |  NNA & TDC  |  KBA  ; 
 OBA <=  NBA & TAC  |  NFA & TBC  |  NJA & TCC  |  NNA & TDC  |  KBA  ; 
 WBA <= IBA ; 
 WFA <= IBA ; 
 WJA <= IBA ; 
 WNA <= IBA ; 
 VBI <=  NBI & TAD  |  NFI & TBD  |  NJI & TCD  |  NNI & TDD  |  KBI  ; 
 OBI <=  NBI & TAD  |  NFI & TBD  |  NJI & TCD  |  NNI & TDD  |  KBI  ; 
 WBI <= IBI ; 
 WFI <= IBI ; 
 WJI <= IBI ; 
 WNI <= IBI ; 
 VCA <=  NCA & TAE  |  NGA & TBE  |  NKA & TCE  |  NOA & TDE  |  KCA  ; 
 OCA <=  NCA & TAE  |  NGA & TBE  |  NKA & TCE  |  NOA & TDE  |  KCA  ; 
 WCA <= ICA ; 
 WGA <= ICA ; 
 WKA <= ICA ; 
 WOA <= ICA ; 
 VCI <=  NCI & TAF  |  NGI & TBF  |  NKI & TCF  |  NOI & TDF  |  KCI  ; 
 OCI <=  NCI & TAF  |  NGI & TBF  |  NKI & TCF  |  NOI & TDF  |  KCI  ; 
 WCI <= ICI ; 
 WGI <= ICI ; 
 WKI <= ICI ; 
 WOI <= ICI ; 
 VDA <=  NDA & TAG  |  NHA & TBG  |  NLA & TCG  |  NPA & TDG  |  KDA  ; 
 ODA <=  NDA & TAG  |  NHA & TBG  |  NLA & TCG  |  NPA & TDG  |  KDA  ; 
 WDA <= IDA ; 
 WHA <= IDA ; 
 WLA <= IDA ; 
 WPA <= IDA ; 
 VDI <=  NDI & TAH  |  NHI & TBH  |  NLI & TCH  |  NPI & TDH  |  KDI  ; 
 ODI <=  NDI & TAH  |  NHI & TBH  |  NLI & TCH  |  NPI & TDH  |  KDI  ; 
 WDI <= IDI ; 
 WHI <= IDI ; 
 WLI <= IDI ; 
 WPI <= IDI ; 
 TAA <= QED & JNA ; 
 TBA <= QED & JNB ; 
 TCA <= QED & JNC ; 
 TDA <= QED & JND ; 
 okj <= qjk ; 
 UAG <= QDA & ZZI ; 
 UAH <= QDA & ZZI ; 
 UDG <= QDA & ZZI ; 
 UDH <= QDA & ZZI ; 
 oea <= iaa ; 
 oei <= iai ; 
 ofa <= iba ; 
 ofi <= ibi ; 
 qha <=  qaa & qba & qca  |  jna  ; 
 QAE <= IGC ; 
 QBE <= QAE ; 
 QCE <= QBE ; 
 QDE <= QCE ; 
 oga <= ica ; 
 ogi <= ici ; 
 oha <= ida ; 
 ohi <= idi ; 
 UBG <= QDA & ZZI ; 
 UBH <= QDA & ZZI ; 
 UCG <= QDA & ZZI ; 
 UCH <= QDA & ZZI ; 
 QBA <= QAA ; 
 QCA <= QBA ; 
 QCI <= QBA ; 
 QDA <= QCA ; 
 qaa <=  igc  |  IGB  |  IGA  ; 
 qab <=  igc  |  IGB  |  iga  ; 
 QPA <=  JMA & TJD  |  QCA  ; 
 QPB <=  JMB & TJD  |  QCB  ; 
 qac <=  igc  |  igb  |  IGA  ; 
 qad <=  igc  |  igb  |  iga  ; 
 PAA <=  PAA & tja & jaa  |  JHA & TJA  |  paa & JAA  ; 
 PAD <=  PAA & tja & jaa  |  JHA & TJA  |  paa & JAA  ; 
 PAG <=  PAA & tja & jaa  |  JHA & TJA  |  paa & JAA  ; 
 PAB <=  PAB & tjb & jab  |  JHB & TJB  |  pab & JAB  ; 
 PAE <=  PAB & tjb & jab  |  JHB & TJB  |  pab & JAB  ; 
 PAH <=  PAB & tjb & jab  |  JHB & TJB  |  pab & JAB  ; 
 PAC <=  PAC & tjc & jac  |  JHC & TJC  |  pac & JAC  ; 
 PAF <=  PAC & tjc & jac  |  JHC & TJC  |  pac & JAC  ; 
 PAI <=  PAC & tjc & jac  |  JHC & TJC  |  pac & JAC  ; 
 UEA <= PBD & TEB |  DAH & teb ; 
 UEB <= PBE & TEB |  DAI & teb ; 
 UEC <= PFA & TEB |  DBE & teb ; 
 UED <= PFB & TEB |  DBF & teb ; 
 UEE <= PBF & TEB |  DAJ & teb ; 
 UEF <= PFC & TEB |  DBG & teb ; 
 ufd <= pfb & TEB |  dbf & teb ; 
 ufe <= pbf & TEB |  daj & teb ; 
 uff <= pfc & TEB |  dbg & teb ; 
 ufa <= pbd & TEB |  dah & teb ; 
 ufb <= pbe & TEB |  dai & teb ; 
 ufc <= pfa & TEB |  dbe & teb ; 
 UGA <= DAM & teb |  PBD & TEB ; 
 UGB <= DAN & teb |  PBE & TEB ; 
 UGC <= DBI & teb |  PGA & TEB ; 
 UGD <= DBJ & teb |  PGB & TEB ; 
 UGE <= DAO & teb |  PBF & TEB ; 
 UGF <= DBK & teb |  PGC & TEB ; 
 uhd <= dbn & teb |  pgb & TEB ; 
 uhe <= dao & teb |  pbf & TEB ; 
 uhf <= dbo & teb |  pgc & TEB ; 
 uha <= dam & teb |  pbd & TEB ; 
 uhb <= dan & teb |  pbe & TEB ; 
 uhc <= dbm & teb |  pga & TEB ; 
 VAB <=  NAB & TAA  |  NEB & TBA  |  NIB & TCA  |  NMB & TDA  |  KAB  ; 
 OAB <=  NAB & TAA  |  NEB & TBA  |  NIB & TCA  |  NMB & TDA  |  KAB  ; 
 WAB <= IAB ; 
 WEB <= IAB ; 
 WIB <= IAB ; 
 WMB <= IAB ; 
 VAJ <=  NAJ & TAB  |  NEJ & TBB  |  NIJ & TCB  |  NMJ & TDB  |  KAJ  ; 
 OAJ <=  NAJ & TAB  |  NEJ & TBB  |  NIJ & TCB  |  NMJ & TDB  |  KAJ  ; 
 WAJ <= IAJ ; 
 WEJ <= IAJ ; 
 WIJ <= IAJ ; 
 WMJ <= IAJ ; 
 VBB <=  NBB & TAC  |  NFB & TBC  |  NJB & TCC  |  NNB & TDC  |  KBB  ; 
 OBB <=  NBB & TAC  |  NFB & TBC  |  NJB & TCC  |  NNB & TDC  |  KBB  ; 
 WBB <= IBB ; 
 WFB <= IBB ; 
 WJB <= IBB ; 
 WNB <= IBB ; 
 VBJ <=  NBJ & TAD  |  NFJ & TBD  |  NJJ & TCD  |  NNJ & TDD  |  KBJ  ; 
 OBJ <=  NBJ & TAD  |  NFJ & TBD  |  NJJ & TCD  |  NNJ & TDD  |  KBJ  ; 
 WBJ <= IBJ ; 
 WFJ <= IBJ ; 
 WJJ <= IBJ ; 
 WNJ <= IBJ ; 
 VCB <=  NCB & TAE  |  NGB & TBE  |  NKB & TCE  |  NOB & TDE  |  KCB  ; 
 OCB <=  NCB & TAE  |  NGB & TBE  |  NKB & TCE  |  NOB & TDE  |  KCB  ; 
 WCB <= ICB ; 
 WGB <= ICB ; 
 WKB <= ICB ; 
 WOB <= ICB ; 
 VCJ <=  NCJ & TAF  |  NGJ & TBF  |  NKJ & TCF  |  NOJ & TDF  |  KCJ  ; 
 OCJ <=  NCJ & TAF  |  NGJ & TBF  |  NKJ & TCF  |  NOJ & TDF  |  KCJ  ; 
 WCJ <= ICJ ; 
 WGJ <= ICJ ; 
 WKJ <= ICJ ; 
 WOJ <= ICJ ; 
 VDB <=  NDB & TAG  |  NHB & TBG  |  NLB & TCG  |  NPB & TDG  |  KDB  ; 
 ODB <=  NDB & TAG  |  NHB & TBG  |  NLB & TCG  |  NPB & TDG  |  KDB  ; 
 WDB <= IDB ; 
 WHB <= IDB ; 
 WLB <= IDB ; 
 WPB <= IDB ; 
 VDJ <=  NDJ & TAH  |  NHJ & TBH  |  NLJ & TCH  |  NPJ & TDH  |  KDJ  ; 
 ODJ <=  NDJ & TAH  |  NHJ & TBH  |  NLJ & TCH  |  NPJ & TDH  |  KDJ  ; 
 WDJ <= IDJ ; 
 WHJ <= IDJ ; 
 WLJ <= IDJ ; 
 WPJ <= IDJ ; 
 ECA <=  ECA & jge  |  JGA & eca  ; 
 EDA <=  ECA & jge  |  JGA & eca  ; 
 EEA <=  ECA & jge  |  JGA & eca  ; 
 ECB <=  ECB & jgf  |  JGB & ecb  ; 
 EDB <=  ECB & jgf  |  JGB & ecb  ; 
 EEB <=  ECB & jgf  |  JGB & ecb  ; 
 ECC <=  ECC & jgg  |  JGC & ecc  ; 
 EDC <=  ECC & jgg  |  JGC & ecc  ; 
 EEC <=  ECC & jgg  |  JGC & ecc  ; 
 TAB <= QED & JNA ; 
 TBB <= QED & JNB ; 
 TCB <= QED & JNC ; 
 TDB <= QED & JND ; 
 UEG <= QDB & ZZI ; 
 UEH <= QDB & ZZI ; 
 UHG <= QDB & ZZI ; 
 UHH <= QDB & ZZI ; 
 oeb <= iab ; 
 oej <= iaj ; 
 ofb <= ibb ; 
 ofj <= ibj ; 
 qhb <=  qab & qbb & qcb  |  jnb  ; 
 ogb <= icb ; 
 ogj <= icj ; 
 ohb <= idb ; 
 ohj <= idj ; 
 UFG <= QDB & ZZI ; 
 UFH <= QDB & ZZI ; 
 UGG <= QDB & ZZI ; 
 UGH <= QDB & ZZI ; 
 QBB <= QAB ; 
 QCB <= QBB ; 
 QCJ <= QBB ; 
 qdb <= qcb ; 
 okk <= daa ; 
 okl <= dae ; 
 okm <= dak ; 
 okn <= dal ; 
 PBA <=  PBA & tja & jba  |  JHA & TJA  |  pba & JBA  ; 
 PBD <=  PBA & tja & jba  |  JHA & TJA  |  pba & JBA  ; 
 PBG <=  PBA & tja & jba  |  JHA & TJA  |  pba & JBA  ; 
 PBB <=  PBB & tjb & jbb  |  JHB & TJB  |  pbb & JBB  ; 
 PBE <=  PBB & tjb & jbb  |  JHB & TJB  |  pbb & JBB  ; 
 PBH <=  PBB & tjb & jbb  |  JHB & TJB  |  pbb & JBB  ; 
 PBC <=  PBC & tjc & jbc  |  JHC & TJC  |  pbc & JBC  ; 
 PBF <=  PBC & tjc & jbc  |  JHC & TJC  |  pbc & JBC  ; 
 PBI <=  PBC & tjc & jbc  |  JHC & TJC  |  pbc & JBC  ; 
 UIA <= PCD & TEC |  DAH & tec ; 
 UIB <= PCE & TEC |  DAI & tec ; 
 UIC <= PFA & TEC |  DBE & tec ; 
 UID <= PFB & TEC |  DBF & tec ; 
 UIE <= PCF & TEC |  DAJ & tec ; 
 UIF <= PFC & TEC |  DBG & tec ; 
 ujd <= pfb & TEC |  dbf & tec ; 
 uje <= pcf & TEC |  daj & tec ; 
 ujf <= pfc & TEC |  dbg & tec ; 
 uja <= pcd & TEC |  dah & tec ; 
 ujb <= pce & TEC |  dai & tec ; 
 ujc <= pfa & TEC |  dbe & tec ; 
 UKA <= DAM & tec |  PCD & TEC ; 
 UKB <= DAN & tec |  PCE & TEC ; 
 UKC <= DBI & tec |  PGA & TEC ; 
 UKD <= DBJ & tec |  PGB & TEC ; 
 UKE <= DAO & tec |  PCF & TEC ; 
 UKF <= DBK & tec |  PGC & TEC ; 
 uld <= dbn & tec |  pgb & TEC ; 
 ule <= dao & tec |  pcf & TEC ; 
 ulf <= dbo & tec |  pgc & TEC ; 
 ula <= dam & tec |  pcd & TEC ; 
 ulb <= dan & tec |  pce & TEC ; 
 ulc <= dbm & tec |  pga & TEC ; 
 VAC <=  NAC & TAA  |  NEC & TBA  |  NIC & TCA  |  NMC & TDA  |  KAC  ; 
 OAC <=  NAC & TAA  |  NEC & TBA  |  NIC & TCA  |  NMC & TDA  |  KAC  ; 
 WAC <= IAC ; 
 WEC <= IAC ; 
 WIC <= IAC ; 
 WMC <= IAC ; 
 VAK <=  NAK & TAB  |  NEK & TBB  |  NIK & TCB  |  NMK & TDB  |  KAK  ; 
 OAK <=  NAK & TAB  |  NEK & TBB  |  NIK & TCB  |  NMK & TDB  |  KAK  ; 
 WAK <= IAK ; 
 WEK <= IAK ; 
 WIK <= IAK ; 
 WMK <= IAK ; 
 VBC <=  NBC & TAC  |  NFC & TBC  |  NJC & TCC  |  NNC & TDC  |  KBC  ; 
 OBC <=  NBC & TAC  |  NFC & TBC  |  NJC & TCC  |  NNC & TDC  |  KBC  ; 
 WBC <= IBC ; 
 WFC <= IBC ; 
 WJC <= IBC ; 
 WNC <= IBC ; 
 VBK <=  NBK & TAD  |  NFK & TBD  |  NJK & TCD  |  NNK & TDD  |  KBK  ; 
 OBK <=  NBK & TAD  |  NFK & TBD  |  NJK & TCD  |  NNK & TDD  |  KBK  ; 
 WBK <= IBK ; 
 WFK <= IBK ; 
 WJK <= IBK ; 
 WNK <= IBK ; 
 VCC <=  NCC & TAE  |  NGC & TBE  |  NKC & TCE  |  NOC & TDE  |  KCC  ; 
 OCC <=  NCC & TAE  |  NGC & TBE  |  NKC & TCE  |  NOC & TDE  |  KCC  ; 
 WCC <= ICC ; 
 WGC <= ICC ; 
 WKC <= ICC ; 
 WOC <= ICC ; 
 VCK <=  NCK & TAF  |  NGK & TBF  |  NKK & TCF  |  NOK & TDF  |  KCK  ; 
 OCK <=  NCK & TAF  |  NGK & TBF  |  NKK & TCF  |  NOK & TDF  |  KCK  ; 
 WCK <= ICK ; 
 WGK <= ICK ; 
 WKK <= ICK ; 
 WOK <= ICK ; 
 VDC <=  NDC & TAG  |  NHC & TBG  |  NLC & TCG  |  NPC & TDG  |  KDC  ; 
 ODC <=  NDC & TAG  |  NHC & TBG  |  NLC & TCG  |  NPC & TDG  |  KDC  ; 
 WDC <= IDC ; 
 WHC <= IDC ; 
 WLC <= IDC ; 
 WPC <= IDC ; 
 VDK <=  NDK & TAH  |  NHK & TBH  |  NLK & TCH  |  NPK & TDH  |  KDK  ; 
 ODK <=  NDK & TAH  |  NHK & TBH  |  NLK & TCH  |  NPK & TDH  |  KDK  ; 
 WDK <= IDK ; 
 WHK <= IDK ; 
 WLK <= IDK ; 
 WPK <= IDK ; 
 QQA <=  QQA & jjh  |  ZZI & QCI  ; 
 QQE <=  QQE & jjh  |  QQA & QCI  ; 
 QQB <=  QQB & jjh  |  ZZI & QCJ  ; 
 QQF <=  QQF & jjh  |  QQB & QCJ  ; 
 TAC <= QED & JNA ; 
 TBC <= QED & JNB ; 
 TCC <= QED & JNC ; 
 TDC <= QED & JND ; 
 QQI <=  JJS & QQA  |  JJT & QQB  |  JJU & QQC  |  JJV & QQD  ; 
 QQJ <=  JJS & QQB  |  JJT & QQC  |  JJU & QQD  |  JJV & QQA  ; 
 QQK <=  JJS & QQC  |  JJT & QQD  |  JJU & QQA  |  JJV & QQB  ; 
 UIG <= QDC & ZZI ; 
 UIH <= QDC & ZZI ; 
 ULG <= QDC & ZZI ; 
 ULH <= QDC & ZZI ; 
 QJH <=  JJA  |  JJB  |  JJC  |  JJD  ; 
 OKB <=  JJA  |  JJB  |  JJC  |  JJD  ; 
 QJI <=  JJE  |  JJF  |  JJG  ; 
 OKC <=  JJE  |  JJF  |  JJG  ; 
 oec <= iac ; 
 oek <= iak ; 
 ofc <= ibc ; 
 ofk <= ibk ; 
 qhc <=  qac & qbc & qcc  |  jnc  ; 
 QJK <=  QJK & jlf & jji  |  QJG  ; 
 ogc <= icc ; 
 ogk <= ick ; 
 ohc <= idc ; 
 ohk <= idk ; 
 UJG <= QDC & ZZI ; 
 UJH <= QDC & ZZI ; 
 UKG <= QDC & ZZI ; 
 UKH <= QDC & ZZI ; 
 QBC <= QAC ; 
 QCC <= QBC ; 
 QCK <= QBC ; 
 QDC <= QCC ; 
 QPC <=  JMC & TJD  |  QCC  ; 
 oko <= dbi ; 
 okp <= dbj ; 
 okq <= dbk ; 
 PCA <=  PCA & tja & jca  |  JHA & TJA  |  pca & JCA  ; 
 PCD <=  PCA & tja & jca  |  JHA & TJA  |  pca & JCA  ; 
 PCG <=  PCA & tja & jca  |  JHA & TJA  |  pca & JCA  ; 
 PCB <=  PCB & tjb & jcb  |  JHB & TJB  |  pcb & JCB  ; 
 PCE <=  PCB & tjb & jcb  |  JHB & TJB  |  pcb & JCB  ; 
 PCH <=  PCB & tjb & jcb  |  JHB & TJB  |  pcb & JCB  ; 
 PCC <=  PCC & tjc & jcc  |  JHC & TJC  |  pcc & JCC  ; 
 PCF <=  PCC & tjc & jcc  |  JHC & TJC  |  pcc & JCC  ; 
 PCI <=  PCC & tjc & jcc  |  JHC & TJC  |  pcc & JCC  ; 
 UMA <= PDD & TED |  DAH & ted ; 
 UMB <= PDE & TED |  DAI & ted ; 
 UMC <= PFA & TED |  DBE & ted ; 
 UMD <= PFB & TED |  DBF & ted ; 
 UME <= PDF & TED |  DAJ & ted ; 
 UMF <= PFC & TED |  DBG & ted ; 
 und <= pfb & TED |  dbf & ted ; 
 une <= pdf & TED |  daj & ted ; 
 unf <= pec & TED |  dbg & ted ; 
 una <= pdd & TED |  dah & ted ; 
 unb <= pde & TED |  dai & ted ; 
 unc <= pfa & TED |  dbe & ted ; 
 UOA <= DAM & ted |  PDD & TED ; 
 UOB <= DAN & ted |  PDE & TED ; 
 UOC <= DBI & ted |  PGA & TED ; 
 UOD <= DBJ & ted |  PGB & TED ; 
 UOE <= DAO & ted |  PDF & TED ; 
 UOF <= DBK & ted |  PGC & TED ; 
 upd <= dbn & ted |  pgb & TED ; 
 upe <= dao & ted |  pdf & TED ; 
 upf <= dbo & ted |  pgc & TED ; 
 upa <= dam & ted |  pdd & TED ; 
 upb <= dan & ted |  pde & TED ; 
 upc <= dbm & ted |  pga & TED ; 
 VAD <=  NAD & TAA  |  NED & TBA  |  NID & TCA  |  NMD & TDA  |  KAD  ; 
 OAD <=  NAD & TAA  |  NED & TBA  |  NID & TCA  |  NMD & TDA  |  KAD  ; 
 WAD <= IAD ; 
 WED <= IAD ; 
 WID <= IAD ; 
 WMD <= IAD ; 
 VAL <=  NAL & TAB  |  NEL & TBB  |  NIL & TCB  |  NML & TDB  |  KAL  ; 
 OAL <=  NAL & TAB  |  NEL & TBB  |  NIL & TCB  |  NML & TDB  |  KAL  ; 
 WAL <= IAL ; 
 WEL <= IAL ; 
 WIL <= IAL ; 
 WML <= IAL ; 
 VBD <=  NBD & TAC  |  NFD & TBC  |  NJD & TCC  |  NND & TDC  |  KBD  ; 
 OBD <=  NBD & TAC  |  NFD & TBC  |  NJD & TCC  |  NND & TDC  |  KBD  ; 
 WBD <= IBD ; 
 WFD <= IBD ; 
 WJD <= IBD ; 
 WND <= IBD ; 
 VBL <=  NBL & TAD  |  NFL & TBD  |  NJL & TCD  |  NNL & TDD  |  KBL  ; 
 OBL <=  NBL & TAD  |  NFL & TBD  |  NJL & TCD  |  NNL & TDD  |  KBL  ; 
 WBL <= IBL ; 
 WFL <= IBL ; 
 WJL <= IBL ; 
 WNL <= IBL ; 
 VCD <=  NCD & TAE  |  NGD & TBE  |  NKD & TCE  |  NOD & TDE  |  KCD  ; 
 OCD <=  NCD & TAE  |  NGD & TBE  |  NKD & TCE  |  NOD & TDE  |  KCD  ; 
 WCD <= ICD ; 
 WGD <= ICD ; 
 WKD <= ICD ; 
 WOD <= ICD ; 
 VCL <=  NCL & TAF  |  NGL & TBF  |  NKL & TCF  |  NOL & TDF  |  KCL  ; 
 OCL <=  NCL & TAF  |  NGL & TBF  |  NKL & TCF  |  NOL & TDF  |  KCL  ; 
 WCL <= ICL ; 
 WGL <= ICL ; 
 WKL <= ICL ; 
 WOL <= ICL ; 
 VDD <=  NDD & TAG  |  NHD & TBG  |  NLD & TCG  |  NPD & TDG  |  KDD  ; 
 ODD <=  NDD & TAG  |  NHD & TBG  |  NLD & TCG  |  NPD & TDG  |  KDD  ; 
 WDD <= IDD ; 
 WHD <= IDD ; 
 WLD <= IDD ; 
 WPD <= IDD ; 
 VDL <=  NDL & TAH  |  NHL & TBH  |  NLL & TCH  |  NPL & TDH  |  KDL  ; 
 ODL <=  NDL & TAH  |  NHL & TBH  |  NLL & TCH  |  NPL & TDH  |  KDL  ; 
 WDL <= IDL ; 
 WHL <= IDL ; 
 WLL <= IDL ; 
 WPL <= IDL ; 
 TEA <= JAD ; 
 TEB <= JBD ; 
 TEC <= JCD ; 
 TED <= JDD ; 
 QQC <=  QQC & jjh  |  ZZI & QCK  ; 
 QQG <=  QQG & jjh  |  QQC & QCK  ; 
 QQD <=  QQD & jjh  |  ZZI & QCL  ; 
 QQH <=  QQH & jjh  |  QQD & QCL  ; 
 TAD <= QED & JNA ; 
 TBD <= QED & JNB ; 
 TCD <= QED & JNC ; 
 TDD <= QED & JND ; 
 QQL <=  JJW & QQH  |  JJX & QQE  |  JJY & QQF  |  JJZ & QQG  ; 
 QQM <=  JJW & QQE  |  JJX & QQF  |  JJY & QQG  |  JJZ & QQH  ; 
 QQN <=  JJW & QQF  |  JJX & QQG  |  JJY & QQH  |  JJZ & QQE  ; 
 QQO <=  JJW & QQG  |  JJX & QQH  |  JJY & QQE  |  JJZ & QQF  ; 
 UMG <= QDD & ZZI ; 
 UMH <= QDD & ZZI ; 
 UPG <= QDD & ZZI ; 
 UPH <= QDD & ZZI ; 
 EFA <=  EFA & jji  |  JIA & QKB  |  QKB & JIC  ; 
 EFB <=  EFB & jji  |  JIB & QKB  |  QKB & JIC  ; 
 oed <= iad ; 
 oel <= ial ; 
 ofd <= ibd ; 
 ofl <= ibl ; 
 qhd <=  qad & qbd & qcd  |  jnd  ; 
 QEB <=  QCA & JIA  |  QCB & JIB  |  QCC & JIC  |  QCD & JID  ; 
 QEF <=  QCA & JIA  |  QCB & JIB  |  QCC & JIC  |  QCD & JID  ; 
 ogd <= icd ; 
 ogl <= icl ; 
 ohd <= idd ; 
 ohl <= idl ; 
 UNG <= QDD & ZZI ; 
 UNH <= QDD & ZZI ; 
 UOG <= QDD & ZZI ; 
 UOH <= QDD & ZZI ; 
 QBD <= QAD ; 
 QCD <= QBD ; 
 QCL <= QBD ; 
 QDD <= QCD ; 
 QKA <= QJN & ZZI ; 
 QKB <= QJN & qka ; 
 okr <= pea ; 
 oks <= peb ; 
 OKT <= PEC ; 
 QPD <= QCD ; 
 PDA <=  PDA & tja & jda  |  JHA & TJA  |  pda & JDA  ; 
 PDD <=  PDA & tja & jda  |  JHA & TJA  |  pda & JDA  ; 
 PDG <=  PDA & tja & jda  |  JHA & TJA  |  pda & JDA  ; 
 PDB <=  PDB & tjb & jdb  |  JHB & TJB  |  pdb & JDB  ; 
 PDE <=  PDB & tjb & jdb  |  JHB & TJB  |  pdb & JDB  ; 
 PDH <=  PDB & tjb & jdb  |  JHB & TJB  |  pdb & JDB  ; 
 PDC <=  PDC & tjc & jdc  |  JHC & TJC  |  pdc & JDC  ; 
 PDF <=  PDC & tjc & jdc  |  JHC & TJC  |  pdc & JDC  ; 
 PDI <=  PDC & tjc & jdc  |  JHC & TJC  |  pdc & JDC  ; 
 UAI <= PAG & TEE |  DAH & tee ; 
 UAJ <= PAH & TEE |  DAI & tee ; 
 UAK <= PFA & TEE |  DBE & tee ; 
 UAL <= PFB & TEE |  DBF & tee ; 
 UAM <= PAI & TEE |  DAJ & tee ; 
 UAN <= PFC & TEE |  DBG & tee ; 
 ubl <= pfb & TEE |  dbf & tee ; 
 ubm <= pai & TEE |  daj & tee ; 
 ubn <= pfc & TEE |  dbg & tee ; 
 ubi <= pag & TEE |  dah & tee ; 
 ubj <= pah & TEE |  dai & tee ; 
 ubk <= pfa & TEE |  dbe & tee ; 
 UCI <= DAC & tee |  PAG & TEE ; 
 UCJ <= DAN & tee |  PAH & TEE ; 
 UCK <= DBI & tee |  PGA & TEE ; 
 UCL <= DBJ & tee |  PGB & TEE ; 
 UCM <= DAO & tee |  PAI & TEE ; 
 UCN <= DBK & tee |  PGC & TEE ; 
 udl <= dbn & tee |  pgb & TEE ; 
 udm <= dao & tee |  pai & TEE ; 
 udn <= dbo & tee |  pgc & TEE ; 
 udi <= dac & tee |  pag & TEE ; 
 udj <= dad & tee |  pah & TEE ; 
 udk <= dbm & tee |  pga & TEE ; 
 VAE <=  NAE & TAA  |  NEE & TBA  |  NIE & TCA  |  NME & TDA  |  KAE  ; 
 OAE <=  NAE & TAA  |  NEE & TBA  |  NIE & TCA  |  NME & TDA  |  KAE  ; 
 WAE <= IAE ; 
 WEE <= IAE ; 
 WIE <= IAE ; 
 WME <= IAE ; 
 VAM <=  NAM & TAB  |  NEM & TBB  |  NIM & TCB  |  NMM & TDB  |  KAM  ; 
 OAM <=  NAM & TAB  |  NEM & TBB  |  NIM & TCB  |  NMM & TDB  |  KAM  ; 
 WAM <= IAM ; 
 WEM <= IAM ; 
 WIM <= IAM ; 
 WMM <= IAM ; 
 VBE <=  NBE & TAC  |  NFE & TBC  |  NJE & TCC  |  NNE & TDC  |  KBE  ; 
 OBE <=  NBE & TAC  |  NFE & TBC  |  NJE & TCC  |  NNE & TDC  |  KBE  ; 
 WBE <= IBE ; 
 WFE <= IBE ; 
 WJE <= IBE ; 
 WNE <= IBE ; 
 VBM <=  NBM & TAD  |  NFM & TBD  |  NJM & TCD  |  NNM & TDD  |  KBM  ; 
 OBM <=  NBM & TAD  |  NFM & TBD  |  NJM & TCD  |  NNM & TDD  |  KBM  ; 
 WBM <= IBM ; 
 WFM <= IBM ; 
 WJM <= IBM ; 
 WNM <= IBM ; 
 VCE <=  NCE & TAE  |  NGE & TBE  |  NKE & TCE  |  NOE & TDE  |  KCE  ; 
 OCE <=  NCE & TAE  |  NGE & TBE  |  NKE & TCE  |  NOE & TDE  |  KCE  ; 
 WCE <= ICE ; 
 WGE <= ICE ; 
 WKE <= ICE ; 
 WOE <= ICE ; 
 VCM <=  NCM & TAF  |  NGM & TBF  |  NKM & TCF  |  NOM & TDF  |  KCM  ; 
 OCM <=  NCM & TAF  |  NGM & TBF  |  NKM & TCF  |  NOM & TDF  |  KCM  ; 
 WCM <= ICM ; 
 WGM <= ICM ; 
 WKM <= ICM ; 
 WOM <= ICM ; 
 VDE <=  NDE & TAG  |  NHE & TBG  |  NLE & TCG  |  NPE & TDG  |  KDE  ; 
 ODE <=  NDE & TAG  |  NHE & TBG  |  NLE & TCG  |  NPE & TDG  |  KDE  ; 
 WDE <= IDE ; 
 WHE <= IDE ; 
 WLE <= IDE ; 
 WPE <= IDE ; 
 VDM <=  NDM & TAH  |  NHM & TBH  |  NLM & TCH  |  NPM & TDH  |  KDM  ; 
 ODM <=  NDM & TAH  |  NHM & TBH  |  NLM & TCH  |  NPM & TDH  |  KDM  ; 
 WDM <= IDM ; 
 WHM <= IDM ; 
 WLM <= IDM ; 
 WPM <= IDM ; 
 DAA <=  DAA & qjt & jfb  |  IFA & QJC  |  EAA & JFB  ; 
 DAF <=  DAA & qjt & jfb  |  IFA & QJC  |  EAA & JFB  ; 
 DAK <=  DAA & qjt & jfb  |  IFA & QJC  |  EAA & JFB  ; 
 DAB <=  DAB & qjt & jfb  |  IFB & QJC  |  EAB & JFB  ; 
 DAG <=  DAB & qjt & jfb  |  IFB & QJC  |  EAB & JFB  ; 
 DAL <=  DAB & qjt & jfb  |  IFB & QJC  |  EAB & JFB  ; 
 DAM <=  DAC & qjt & jfb  |  IFC & QJC  |  EAC & JFB  ; 
 DAH <=  DAC & qjt & jfb  |  IFC & QJC  |  EAC & JFB  ; 
 DAC <=  DAC & qjt & jfb  |  IFC & QJC  |  EAC & JFB  ; 
 TAE <= QED & JNA ; 
 TBE <= QED & JNB ; 
 TCE <= QED & JNC ; 
 TDE <= QED & JND ; 
 DAN <=  DAD & qjt & jfc  |  IFD & QJC  |  EAD & JFC  ; 
 DAI <=  DAD & qjt & jfc  |  IFD & QJC  |  EAD & JFC  ; 
 DAD <=  DAD & qjt & jfc  |  IFD & QJC  |  EAD & JFC  ; 
 DAO <=  DAE & qjt & jfc  |  IFE & QJC  |  EAE & JFC  ; 
 DAJ <=  DAE & qjt & jfc  |  IFE & QJC  |  EAE & JFC  ; 
 DAE <=  DAE & qjt & jfc  |  IFE & QJC  |  EAE & JFC  ; 
 UAO <= QDA & ZZI ; 
 UAP <= QDA & ZZI ; 
 UDO <= QDA & ZZI ; 
 UDP <= QDA & ZZI ; 
 EAA <=  DAA & jxb & jea  |  daa & JEA  |  EAA & QLB  ; 
 EAB <=  DAB & jxb & jeb  |  dab & JEB  |  EAB & QLB  ; 
 EAC <=  DAC & jxb & jec  |  dac & JEC  |  EAC & QLB  ; 
 oee <= iae ; 
 oem <= iam ; 
 ofe <= ibe ; 
 ofm <= ibm ; 
 UBO <= QDA & ZZI ; 
 UBP <= QDA & ZZI ; 
 UCO <= QDA & ZZI ; 
 UCP <= QDA & ZZI ; 
 EAE <=  DAE & jxb & jee  |  dae & JEE  |  EAE & QLB  ; 
 EAD <=  DAD & jxb & jed  |  dad & JED  |  EAD & QLB  ; 
 oge <= ice ; 
 ogm <= icm ; 
 ohe <= ide ; 
 ohm <= idm ; 
 qld <= ijf & jpe ; 
 UEI <= PBG & TEF |  DAH & tef ; 
 UEJ <= PBH & TEF |  DAI & tef ; 
 UEK <= PFA & TEF |  DBE & tef ; 
 UEL <= PFB & TEF |  DBF & tef ; 
 UEM <= PBI & TEF |  DAJ & tef ; 
 UEN <= PFC & TEF |  DBG & tef ; 
 ufl <= pfb & TEF |  dbf & tef ; 
 ufm <= pbi & TEF |  daj & tef ; 
 ufn <= pfc & TEF |  dbg & tef ; 
 ufi <= pbg & TEF |  dah & tef ; 
 ufj <= pbh & TEF |  dai & tef ; 
 ufk <= pfa & TEF |  dbe & tef ; 
 UGI <= DAM & tef |  PBG & TEF ; 
 UGJ <= DAN & tef |  PBH & TEF ; 
 UGK <= DBI & tef |  PGA & TEF ; 
 UGL <= DBJ & tef |  PGB & TEF ; 
 UGM <= DAO & tef |  PBI & TEF ; 
 UGN <= DBK & tef |  PGC & TEF ; 
 uhl <= dbn & tef |  pgb & TEF ; 
 uhm <= dao & tef |  pbi & TEF ; 
 uhn <= dbo & tef |  pgc & TEF ; 
 uhi <= dac & tef |  pbg & TEF ; 
 uhj <= dan & tef |  pbh & TEF ; 
 uhk <= dbm & tef |  pga & TEF ; 
 VAF <=  NAF & TAA  |  NEF & TBA  |  NIF & TCA  |  NMF & TDA  |  KAF  ; 
 OAF <=  NAF & TAA  |  NEF & TBA  |  NIF & TCA  |  NMF & TDA  |  KAF  ; 
 WAF <= IAF ; 
 WEF <= IAF ; 
 WIF <= IAF ; 
 WMF <= IAF ; 
 VAN <=  NAN & TAB  |  NEN & TBB  |  NIN & TCB  |  NMN & TDB  |  KAN  ; 
 OAN <=  NAN & TAB  |  NEN & TBB  |  NIN & TCB  |  NMN & TDB  |  KAN  ; 
 WAN <= IAN ; 
 WEN <= IAN ; 
 WIN <= IAN ; 
 WMN <= IAN ; 
 VBF <=  NBF & TAC  |  NFF & TBC  |  NJF & TCC  |  NNF & TDC  |  KBF  ; 
 OBF <=  NBF & TAC  |  NFF & TBC  |  NJF & TCC  |  NNF & TDC  |  KBF  ; 
 WBF <= IBF ; 
 WFF <= IBF ; 
 WJF <= IBF ; 
 WNF <= IBF ; 
 VBN <=  NBN & TAD  |  NFN & TBD  |  NJN & TCD  |  NNN & TDD  |  KBN  ; 
 OBN <=  NBN & TAD  |  NFN & TBD  |  NJN & TCD  |  NNN & TDD  |  KBN  ; 
 WBN <= IBN ; 
 WFN <= IBN ; 
 WJN <= IBN ; 
 WNN <= IBN ; 
 VCF <=  NCF & TAE  |  NGF & TBE  |  NKF & TCE  |  NOF & TDE  |  KCF  ; 
 OCF <=  NCF & TAE  |  NGF & TBE  |  NKF & TCE  |  NOF & TDE  |  KCF  ; 
 WCF <= ICF ; 
 WGF <= ICF ; 
 WKF <= ICF ; 
 WOF <= ICF ; 
 VCN <=  NCN & TAF  |  NGN & TBF  |  NKN & TCF  |  NON & TDF  |  KCN  ; 
 OCN <=  NCN & TAF  |  NGN & TBF  |  NKN & TCF  |  NON & TDF  |  KCN  ; 
 WCN <= ICN ; 
 WGN <= ICN ; 
 WKN <= ICN ; 
 WON <= ICN ; 
 VDF <=  NDF & TAG  |  NHF & TBG  |  NLF & TCG  |  NPF & TDG  |  KDF  ; 
 ODF <=  NDF & TAG  |  NHF & TBG  |  NLF & TCG  |  NPF & TDG  |  KDF  ; 
 WDF <= IDF ; 
 WHF <= IDF ; 
 WLF <= IDF ; 
 WPF <= IDF ; 
 VDN <=  NDN & TAH  |  NHN & TBH  |  NLN & TCH  |  NPN & TDH  |  KDN  ; 
 ODN <=  NDN & TAH  |  NHN & TBH  |  NLN & TCH  |  NPN & TDH  |  KDN  ; 
 WDN <= IDN ; 
 WHN <= IDN ; 
 WLN <= IDN ; 
 WPN <= IDN ; 
 oki <= qje ; 
 TAF <= QED & JNA ; 
 TBF <= QED & JNB ; 
 TCF <= QED & JNC ; 
 TDF <= QED & JND ; 
 DBA <=  DBA & jfa  |  IEA & IED  |  IEE & IEH  |  EBA & QLF  ; 
 DBE <=  DBA & jfa  |  IEA & IED  |  IEE & IEH  |  EBA & QLF  ; 
 DBB <=  DBB & jfa  |  IEB & IED  |  IEF & IEH  |  EBB & QLF  ; 
 DBF <=  DBB & jfa  |  IEB & IED  |  IEF & IEH  |  EBB & QLF  ; 
 DBC <=  DBC & jfa  |  IEC & IED  |  IEG & IEH  |  EBC & QLF  ; 
 DBG <=  DBC & jfa  |  IEC & IED  |  IEG & IEH  |  EBC & QLF  ; 
 DBI <=  DBA & jfa  |  IEA & IEI  |  IEE & IEJ  |  EBA & QLF  ; 
 DBM <=  DBA & jfa  |  IEA & IEI  |  IEE & IEJ  |  EBA & QLF  ; 
 DBJ <=  DBB & jfa  |  IEB & IEI  |  IEF & IEJ  |  EBB & QLG  ; 
 DBN <=  DBB & jfa  |  IEB & IEI  |  IEF & IEJ  |  EBB & QLG  ; 
 DBK <=  DBC & jfa  |  IEC & IEI  |  IEG & IEJ  |  EBC & QLG  ; 
 DBO <=  DBC & jfa  |  IEC & IEI  |  IEG & IEJ  |  EBC & QLG  ; 
 UEO <= QDB & ZZI ; 
 UEP <= QDB & ZZI ; 
 UHO <= QDB & ZZI ; 
 UHP <= QDB & ZZI ; 
 QJD <=  ijd & ije & QJD  |  JEF & JPF  ; 
 OKH <=  ijd & ije & QJD  |  JEF & JPF  ; 
 qec <=  QJE & jjj  |  ijd & jpc  |  jpd  ; 
 qed <=  QJE & jjj  |  ijd & jpc  |  jpd  ; 
 qee <=  QJE & jjj  |  ijd & jpc  |  jpd  ; 
 oef <= iaf ; 
 oen <= ian ; 
 off <= ibf ; 
 ofn <= ibn ; 
 QJP <=  QJP & jpg & ija  |  IJE & ija  ; 
 QJF <=  QJF & jpe  |  IHB  |  IJD  |  QJG  ; 
 ogf <= icf ; 
 ogn <= icn ; 
 ohf <= idf ; 
 ohn <= idn ; 
 UFO <= QDB & ZZI ; 
 UFP <= QDB & ZZI ; 
 UGO <= QDB & ZZI ; 
 UGP <= QDB & ZZI ; 
 QJM <=  QJM & qeb & ija  |  IJE & ija  ; 
 QJN <=  QJM & qeb & ija  |  IJE & ija  ; 
 OKA <=  QJM & qeb & ija  |  IJE & ija  ; 
 QJC <=  IJB & IJG  |  ZZO & qja  |  ZZO & QJU  ; 
 QJT <=  IJB & IJG  |  QJW & qja  |  IJF & QJU  ; 
 QJE <=  QJE & jlf  |  IJE  ; 
 QJG <=  IJE & jlf  ; 
 QJO <=  QJQ  |  QJO & qjx  ; 
 QJL <=  IJE  ; 
 TJA <= QJL ; 
 TJB <= QJL ; 
 TJC <= QJL ; 
 TJD <= QJL ; 
 QLF <= qju & IJF ; 
 QLG <= qju & IJF ; 
 UII <= PCG & TEG |  DAH & teg ; 
 UIJ <= PCH & TEG |  DAI & teg ; 
 UIK <= PEA & TEG |  DBE & teg ; 
 UIL <= PEB & TEG |  DBF & teg ; 
 UIM <= PCI & TEG |  DAJ & teg ; 
 UIN <= PFC & TEG |  DBG & teg ; 
 ujl <= pfb & TEG |  dbf & teg ; 
 ujm <= pci & TEG |  daj & teg ; 
 ujn <= pfc & TEG |  dbg & teg ; 
 uji <= pcg & TEG |  dah & teg ; 
 ujj <= pch & TEG |  dai & teg ; 
 ujk <= pfa & TEG |  dbe & teg ; 
 UKI <= DAM & teg |  PCG & TEG ; 
 UKJ <= DAN & teg |  PCH & TEG ; 
 UKK <= DBI & teg |  PGA & TEG ; 
 UKL <= DBJ & teg |  PGB & TEG ; 
 UKM <= DAO & teg |  PCI & TEG ; 
 UKN <= DBK & teg |  PGC & TEG ; 
 ull <= dbn & teg |  pgb & TEG ; 
 ulm <= dao & teg |  pci & TEG ; 
 uln <= dbo & teg |  pgc & TEG ; 
 uli <= dam & teg |  pcg & TEG ; 
 ulj <= dan & teg |  pch & TEG ; 
 ulk <= dbm & teg |  pga & TEG ; 
 VAG <=  NAG & TAA  |  NEG & TBA  |  NIG & TCA  |  NMG & TDA  |  KAG  ; 
 OAG <=  NAG & TAA  |  NEG & TBA  |  NIG & TCA  |  NMG & TDA  |  KAG  ; 
 WAG <= IAG ; 
 WEG <= IAG ; 
 WIG <= IAG ; 
 WMG <= IAG ; 
 VAO <=  NAO & TAB  |  NEO & TBB  |  NIO & TCB  |  NMO & TDB  |  KAO  ; 
 OAO <=  NAO & TAB  |  NEO & TBB  |  NIO & TCB  |  NMO & TDB  |  KAO  ; 
 WAO <= IAO ; 
 WEO <= IAO ; 
 WIO <= IAO ; 
 WMO <= IAO ; 
 VBG <=  NBG & TAC  |  NFG & TBC  |  NJG & TCC  |  NNG & TDC  |  KBG  ; 
 OBG <=  NBG & TAC  |  NFG & TBC  |  NJG & TCC  |  NNG & TDC  |  KBG  ; 
 WBG <= IBG ; 
 WFG <= IBG ; 
 WJG <= IBG ; 
 WNG <= IBG ; 
 VBO <=  NBO & TAD  |  NFO & TBD  |  NJO & TCD  |  NNO & TDD  |  KBO  ; 
 OBO <=  NBO & TAD  |  NFO & TBD  |  NJO & TCD  |  NNO & TDD  |  KBO  ; 
 WBO <= IBO ; 
 WFO <= IBO ; 
 WJO <= IBO ; 
 WNO <= IBO ; 
 VCG <=  NCG & TAE  |  NGG & TBE  |  NKG & TCE  |  NOG & TDE  |  KCG  ; 
 OCG <=  NCG & TAE  |  NGG & TBE  |  NKG & TCE  |  NOG & TDE  |  KCG  ; 
 WCG <= ICG ; 
 WGG <= ICG ; 
 WKG <= ICG ; 
 WOG <= ICG ; 
 VCO <=  NCO & TAF  |  NGO & TBF  |  NKO & TCF  |  NOO & TDF  |  KCO  ; 
 OCO <=  NCO & TAF  |  NGO & TBF  |  NKO & TCF  |  NOO & TDF  |  KCO  ; 
 WCO <= ICO ; 
 WGO <= ICO ; 
 WKO <= ICO ; 
 WOO <= ICO ; 
 VDG <=  NDG & TAG  |  NHG & TBG  |  NLG & TCG  |  NPG & TDG  |  KDG  ; 
 ODG <=  NDG & TAG  |  NHG & TBG  |  NLG & TCG  |  NPG & TDG  |  KDG  ; 
 WDG <= IDG ; 
 WHG <= IDG ; 
 WLG <= IDG ; 
 WPG <= IDG ; 
 VDO <=  NDO & TAH  |  NHO & TBH  |  NLO & TCH  |  NPO & TDH  |  KDO  ; 
 ODO <=  NDO & TAH  |  NHO & TBH  |  NLO & TCH  |  NPO & TDH  |  KDO  ; 
 WDO <= IDO ; 
 WHO <= IDO ; 
 WLO <= IDO ; 
 WPO <= IDO ; 
 TEE <= JAD ; 
 TEF <= JBD ; 
 TEG <= JCD ; 
 TEH <= JDD ; 
 TAG <= QED & JNA ; 
 TBG <= QED & JNB ; 
 TCG <= QED & JNC ; 
 TDG <= QED & JND ; 
 FAA <=  FAA & jlx & jla  |  JLA & faa  ; 
 FBA <=  FAA & jlx & jla  |  JLA & faa  ; 
 QJV <= QJU & ZZI ; 
 QJW <= QJU & qjv ; 
 UIO <= QDC & ZZI ; 
 UIP <= QDC & ZZI ; 
 ULO <= QDC & ZZI ; 
 ULP <= QDC & ZZI ; 
 FAB <=  FAB & tjd & jlb  |  JLB & fab  ; 
 FBB <=  FAB & tjd & jlb  |  JLB & fab  ; 
 oeg <= iag ; 
 oeo <= iao ; 
 ofg <= ibg ; 
 ofo <= ibo ; 
 ogg <= icg ; 
 ogo <= ico ; 
 ohg <= idg ; 
 oho <= ido ; 
 UJO <= QDC & ZZI ; 
 UJP <= QDC & ZZI ; 
 UKO <= QDC & ZZI ; 
 UKP <= QDC & ZZI ; 
 qja <= ijb ; 
 QJB <= QJA ; 
 QJR <= QJQ ; 
 qjz <= ijb ; 
 OJA <= JPE ; 
 OKG <= JPC ; 
 OJD <= JLF ; 
 qjj <= ijb ; 
 PEA <=  PEA & qjx  |  QJX & PXA  ; 
 PFA <=  PEA & qjx  |  QJX & PXA  ; 
 PGA <=  PEA & qjx  |  QJX & PXA  ; 
 QJX <= qjs & QJO ; 
 QJY <= qjs & QJO ; 
 OJB <=  QJU & ijd & ije  |  QJD & IHB  ; 
 QJU <=  QJU & ijd & ije  |  QJD & IHB  ; 
 OJF <=  QJU & ijd & ije  |  QJD & IHB  ; 
 PXA <= PXA & qjq |  DBA & QJQ ; 
 PXB <= PXB & qjq |  DBB & QJQ ; 
 PXC <= PXC & qjq |  DBC & QJQ ; 
 PEB <=  PEB & qjx  |  QJX & PXB  ; 
 PFB <=  PEB & qjx  |  QJX & PXB  ; 
 PGB <=  PEB & qjx  |  QJX & PXB  ; 
 PEC <=  PEC & qjx  |  QJX & PXC  ; 
 PFC <=  PEC & qjx  |  QJX & PXC  ; 
 PGC <=  PEC & qjx  |  QJX & PXC  ; 
 QLH <= QLJ ; 
 qlj <= ijf ; 
 QJQ <= QJE ; 
 QJS <= QJR ; 
 UMI <= PDG & TEH |  DAH & teh ; 
 UMJ <= PDH & TEH |  DAI & teh ; 
 UMK <= PFA & TEH |  DBE & teh ; 
 UML <= PFB & TEH |  DBF & teh ; 
 UMM <= PDI & TEH |  DAJ & teh ; 
 UMN <= PFC & TEH |  DBG & teh ; 
 unl <= pfb & TEH |  dbf & teh ; 
 unm <= pdi & TEH |  daj & teh ; 
 unn <= pfc & TEH |  dbg & teh ; 
 uni <= pdg & TEH |  dah & teh ; 
 unj <= pdh & TEH |  dai & teh ; 
 unk <= pfa & TEH |  dbe & teh ; 
 UOI <= DAM & teh |  PDG & TEH ; 
 UOJ <= DAN & teh |  PDH & TEH ; 
 UOK <= DBI & teh |  PGA & TEH ; 
 UOL <= DBJ & teh |  PGB & TEH ; 
 UOM <= DAO & teh |  PDI & TEH ; 
 UON <= DBK & teh |  PGC & TEH ; 
 upl <= dbn & teh |  pgb & TEH ; 
 upm <= dao & teh |  pdi & TEH ; 
 upn <= dbo & teh |  pgc & TEH ; 
 upi <= dam & teh |  pdg & TEH ; 
 upj <= dan & teh |  pdh & TEH ; 
 upk <= dbm & teh |  pga & TEH ; 
 VAH <=  NAH & TAA  |  NEH & TBA  |  NIH & TCA  |  NMH & TDA  |  KAH  ; 
 OAH <=  NAH & TAA  |  NEH & TBA  |  NIH & TCA  |  NMH & TDA  |  KAH  ; 
 WAH <= IAH ; 
 WEH <= IAH ; 
 WIH <= IAH ; 
 WMH <= IAH ; 
 VAP <=  NAP & TAB  |  NEP & TBB  |  NIP & TCB  |  NMP & TDB  |  KAP  ; 
 OAP <=  NAP & TAB  |  NEP & TBB  |  NIP & TCB  |  NMP & TDB  |  KAP  ; 
 WAP <= IAP ; 
 WEP <= IAP ; 
 WIP <= IAP ; 
 WMP <= IAP ; 
 VBH <=  NBH & TAC  |  NFH & TBC  |  NJH & TCC  |  NNH & TDC  |  KBH  ; 
 OBH <=  NBH & TAC  |  NFH & TBC  |  NJH & TCC  |  NNH & TDC  |  KBH  ; 
 WBH <= IBH ; 
 WFH <= IBH ; 
 WJH <= IBH ; 
 WNH <= IBH ; 
 VBP <=  NBP & TAD  |  NFP & TBD  |  NJP & TCD  |  NNP & TDD  |  KBP  ; 
 OBP <=  NBP & TAD  |  NFP & TBD  |  NJP & TCD  |  NNP & TDD  |  KBP  ; 
 WBP <= IBP ; 
 WFP <= IBP ; 
 WJP <= IBP ; 
 WNP <= IBP ; 
 VCH <=  NCH & TAE  |  NGH & TBE  |  NKH & TCE  |  NOH & TDE  |  KCH  ; 
 OCH <=  NCH & TAE  |  NGH & TBE  |  NKH & TCE  |  NOH & TDE  |  KCH  ; 
 WCH <= ICH ; 
 WGH <= ICH ; 
 WKH <= ICH ; 
 WOH <= ICH ; 
 VCP <=  NCP & TAF  |  NGP & TBF  |  NKP & TCF  |  NOP & TDF  |  KCP  ; 
 OCP <=  NCP & TAF  |  NGP & TBF  |  NKP & TCF  |  NOP & TDF  |  KCP  ; 
 WCP <= ICP ; 
 WGP <= ICP ; 
 WKP <= ICP ; 
 WOP <= ICP ; 
 VDH <=  NDH & TAG  |  NHH & TBG  |  NLH & TCG  |  NPH & TDG  |  KDH  ; 
 ODH <=  NDH & TAG  |  NHH & TBG  |  NLH & TCG  |  NPH & TDG  |  KDH  ; 
 WDH <= IDH ; 
 WHH <= IDH ; 
 WLH <= IDH ; 
 WPH <= IDH ; 
 VDP <=  NDP & TAH  |  NHP & TBH  |  NLP & TCH  |  NPP & TDH  |  KDP  ; 
 ODP <=  NDP & TAH  |  NHP & TBH  |  NLP & TCH  |  NPP & TDH  |  KDP  ; 
 WDP <= IDP ; 
 WHP <= IDP ; 
 WLP <= IDP ; 
 WPP <= IDP ; 
 tfa <= qef & ZZI ; 
 tfe <= qef & ZZI ; 
 TGA <= qef & qee ; 
 TGE <= qef & qee ; 
 TAH <= QED & JNA ; 
 TBH <= QED & JNB ; 
 TCH <= QED & JNC ; 
 TDH <= QED & JND ; 
 tfb <= qef & ZZI ; 
 tff <= qef & ZZI ; 
 TGB <= qef & qee ; 
 TGF <= qef & qee ; 
 FAC <=  FAC & jlx & jlc  |  JLC & fac  ; 
 FBC <=  FAC & jlx & jlc  |  JLC & fac  ; 
 oku <= faa ; 
 okv <= fab ; 
 UMO <= QDD & ZZI ; 
 UMP <= QDD & ZZI ; 
 UPO <= QDD & ZZI ; 
 UPP <= QDD & ZZI ; 
 FAD <=  FAD & tjd & jld  |  JLD & fad  ; 
 FBD <=  FAD & tjd & jld  |  JLD & fad  ; 
 oeh <= iah ; 
 oep <= iap ; 
 ofh <= ibh ; 
 ofp <= ibp ; 
 tfc <= qef & ZZI ; 
 tfg <= qef & ZZI ; 
 TGC <= qef & qee ; 
 TGG <= qef & qee ; 
 FAE <=  FAE & tjd & jle  |  JLE & fae  ; 
 FBE <=  FAE & tjd & jle  |  JLE & fae  ; 
 ogh <= ich ; 
 ogp <= icp ; 
 ohh <= idh ; 
 ohp <= idp ; 
 UNO <= QDD & ZZI ; 
 UNP <= QDD & ZZI ; 
 UOO <= QDD & ZZI ; 
 UOP <= QDD & ZZI ; 
 TMA <= IHA ; 
 qlb <=  qjb & jxa  |  ZZI & IJF  |  QLD  |  IJD  ; 
 tfd <= qef & ZZI ; 
 tfh <= qef & ZZI ; 
 TGD <= qef & qee ; 
 TGH <= qef & qee ; 
 qla <=  qja  |  IJD  ; 
 okw <= fac ; 
 okx <= fad ; 
 eba <= dba & qlb |  eba & QLB ; 
 ebb <= dbb & qlb |  ebb & QLB ; 
 ebc <= dbc & qlb |  ebc & QLB ; 
end
ram_16x4 rinst_0(RAA,RAB,RAC,RAD,WAA,WAB,WAC,WAD,uaa,uab,uac,uad, GAA, UAG, IZZ); 
ram_16x4 rinst_1(SAA,SAB,SAC,SAD,WEA,WEB,WEC,WED,uaa,uab,uac,uad, GAB, UAG, IZZ); 
ram_16x4 rinst_2(XAA,XAB,XAC,XAD,WIA,WIB,WIC,WID,uaa,uab,uac,uad, GAC, UAG, IZZ); 
ram_16x4 rinst_3(RAI,RAJ,RAK,RAL,WAI,WAJ,WAK,WAL,UAA,UAB,UAC,UAD, GAA, UAH, IZZ); 
ram_16x4 rinst_4(SAI,SAJ,SAK,SAL,WEI,WEJ,WEK,WEL,UAA,UAB,UAC,UAD, GAB, UAH, IZZ); 
ram_16x4 rinst_5(RBA,RBB,RBC,RBD,WBA,WBB,WBC,WBD,uba,ubb,ubc,ubd, GBA, UBG, IZZ); 
ram_16x4 rinst_6(SBA,SBB,SBC,SBD,WFA,WFB,WFC,WFD,uba,ubb,ubc,ubd, GBB, UBG, IZZ); 
ram_16x4 rinst_7(XBA,XBB,XBC,XBD,WJA,WJB,WJC,WJD,uba,ubb,ubc,ubd, GBC, UBG, IZZ); 
ram_16x4 rinst_8(XBI,XBJ,XBK,XBL,WJI,WJJ,WJK,WJL,UBA,UBB,UBC,UBD, GBC, UBH, IZZ); 
ram_16x4 rinst_9(YBI,YBJ,YBK,YBL,WNI,WNJ,WNK,WNL,UBA,UBB,UBC,UBD, GBD, UBH, IZZ); 
ram_16x4 rinst_10(RCA,RCB,RCC,RCD,WCA,WCB,WCC,WCD,uca,ucb,ucc,ucd, GCA, UCG, IZZ); 
ram_16x4 rinst_11(SCA,SCB,SCC,SCD,WGA,WGB,WGC,WGD,uca,ucb,ucc,ucd, GCB, UCG, IZZ); 
ram_16x4 rinst_12(RCI,RCJ,RCK,RCL,WCI,WCJ,WCK,WCL,UCA,UCB,UCC,UCD, GCA, UCH, IZZ); 
ram_16x4 rinst_13(SCI,SCJ,SCK,SCL,WGI,WGJ,WGK,WGL,UCA,UCB,UCC,UCD, GCB, UCH, IZZ); 
ram_16x4 rinst_14(XCI,XCJ,XCK,XCL,WKI,WKJ,WKK,WKL,UCA,UCB,UCC,UCD, GCC, UCH, IZZ); 
ram_16x4 rinst_15(RDA,RDB,RDC,RDD,WDA,WDB,WDC,WDD,uda,udb,udc,udd, GDA, UDG, IZZ); 
ram_16x4 rinst_16(SDA,SDB,SDC,SDD,WHA,WHB,WHC,WHD,uda,udb,udc,udd, GDB, UDG, IZZ); 
ram_16x4 rinst_17(RDI,RDJ,RDK,RDL,WDI,WDJ,WDK,WDL,UDA,UDB,UDC,UDD, GDA, UDH, IZZ); 
ram_16x4 rinst_18(SDI,SDJ,SDK,SDL,WHI,WHJ,WHK,WHL,UDA,UDB,UDC,UDD, GDB, UDH, IZZ); 
ram_16x4 rinst_19(XDI,XDJ,XDK,XDL,WLI,WLJ,WLK,WLL,UDA,UDB,UDC,UDD, GDC, UDH, IZZ); 
ram_16x4 rinst_20(YAA,YAB,YAC,YAD,WMA,WMB,WMC,WMD,uaa,uab,uac,uad, GAD, UAG, IZZ); 
ram_16x4 rinst_21(XAI,XAJ,XAK,XAL,WII,WIJ,WIK,WIL,UAA,UAB,UAC,UAD, GAC, UAH, IZZ); 
ram_16x4 rinst_22(YAI,YAJ,YAK,YAL,WMI,WMJ,WMK,WML,UAA,UAB,UAC,UAD, GAD, UAH, IZZ); 
ram_16x4 rinst_23(YBA,YBB,YBC,YBD,WNA,WNB,WNC,WND,uba,ubb,ubc,ubd, GBD, UBG, IZZ); 
ram_16x4 rinst_24(RBI,RBJ,RBK,RBL,WBI,WBJ,WBK,WBL,UBA,UBB,UBC,UBD, GBA, UBH, IZZ); 
ram_16x4 rinst_25(SBI,SBJ,SBK,SBL,WFI,WFJ,WFK,WFL,UBA,UBB,UBC,UBD, GBB, UBH, IZZ); 
ram_16x4 rinst_26(XCA,XCB,XCC,XCD,WKA,WKB,WKC,WKD,uca,ucb,ucc,ucd, GCC, UCG, IZZ); 
ram_16x4 rinst_27(YCA,YCB,YCC,YCD,WOA,WOB,WOC,WOD,uca,ucb,ucc,ucd, GCD, UCG, IZZ); 
ram_16x4 rinst_28(YCI,YCJ,YCK,YCL,WOI,WOJ,WOK,WOL,UCA,UCB,UCC,UCD, GCD, UCH, IZZ); 
ram_16x4 rinst_29(XDA,XDB,XDC,XDD,WLA,WLB,WLC,WLD,uda,udb,udc,udd, GDC, UDG, IZZ); 
ram_16x4 rinst_30(YDA,YDB,YDC,YDD,WPA,WPB,WPC,WPD,uda,udb,udc,udd, GDD, UDG, IZZ); 
ram_16x4 rinst_31(YDI,YDJ,YDK,YDL,WPI,WPJ,WPK,WPL,UDA,UDB,UDC,UDD, GDD, UDH, IZZ); 
ram_16x4 rinst_32(REA,REB,REC,RED,WAA,WAB,WAC,WAD,uea,ueb,uec,ued, GEA, UEG, IZZ); 
ram_16x4 rinst_33(SEA,SEB,SEC,SED,WEA,WEB,WEC,WED,uea,ueb,uec,ued, GEB, UEG, IZZ); 
ram_16x4 rinst_34(XEA,XEB,XEC,XED,WIA,WIB,WIC,WID,uea,ueb,uec,ued, GEC, UEG, IZZ); 
ram_16x4 rinst_35(REI,REJ,REK,REL,WAI,WAJ,WAK,WAL,UEA,UEB,UEC,UED, GEA, UEH, IZZ); 
ram_16x4 rinst_36(SEI,SEJ,SEK,SEL,WEI,WEJ,WEK,WEL,UEA,UEB,UEC,UED, GEB, UEH, IZZ); 
ram_16x4 rinst_37(RFA,RFB,RFC,RFD,WBA,WBB,WBC,WBD,ufa,ufb,ufc,ufd, GFA, UFG, IZZ); 
ram_16x4 rinst_38(SFA,SFB,SFC,SFD,WFA,WFB,WFC,WFD,ufa,ufb,ufc,ufd, GFB, UFG, IZZ); 
ram_16x4 rinst_39(XFA,XFB,XFC,XFD,WJA,WJB,WJC,WJD,ufa,ufb,ufc,ufd, GFC, UFG, IZZ); 
ram_16x4 rinst_40(RFI,RFJ,RFK,RFL,WBI,WBJ,WBK,WBL,UFA,UFB,UFC,UFD, GFA, UFH, IZZ); 
ram_16x4 rinst_41(SFI,SFJ,SFK,SFL,WFI,WFJ,WFK,WFL,UFA,UFB,UFC,UFD, GFB, UFH, IZZ); 
ram_16x4 rinst_42(RGA,RGB,RGC,RGD,WCA,WCB,WCC,WCD,uga,ugb,ugc,ugd, GGA, UGG, IZZ); 
ram_16x4 rinst_43(SGA,SGB,SGC,SGD,WGA,WGB,WGC,WGD,uga,ugb,ugc,ugd, GGB, UGG, IZZ); 
ram_16x4 rinst_44(RGI,RGJ,RGK,RGL,WCI,WCJ,WCK,WCL,UGA,UGB,UGC,UGD, GGA, UGH, IZZ); 
ram_16x4 rinst_45(SGI,SGJ,SGK,SGL,WGI,WGJ,WGK,WGL,UGA,UGB,UGC,UGD, GGB, UGH, IZZ); 
ram_16x4 rinst_46(XGI,XGJ,XGK,XGL,WKI,WKJ,WKK,WKL,UGA,UGB,UGC,UGD, GGC, UGH, IZZ); 
ram_16x4 rinst_47(RHA,RHB,RHC,RHD,WDA,WDB,WDC,WDD,uha,uhb,uhc,uhd, GHA, UHG, IZZ); 
ram_16x4 rinst_48(SHA,SHB,SHC,SHD,WHA,WHB,WHC,WHD,uha,uhb,uhc,uhd, GHB, UHG, IZZ); 
ram_16x4 rinst_49(RHI,RHJ,RHK,RHL,WDI,WDJ,WDK,WDL,UHA,UHB,UHC,UHD, GHA, UHH, IZZ); 
ram_16x4 rinst_50(SHI,SHJ,SHK,SHL,WHI,WHJ,WHK,WHL,UHA,UHB,UHC,UHD, GHB, UHH, IZZ); 
ram_16x4 rinst_51(XHI,XHJ,XHK,XHL,WLI,WLJ,WLK,WLL,UHA,UHB,UHC,UHD, GHC, UHH, IZZ); 
ram_16x4 rinst_52(YEA,YEB,YEC,YED,WMA,WMB,WMC,WMD,uea,ueb,uec,ued, GED, UEG, IZZ); 
ram_16x4 rinst_53(XEI,XEJ,XEK,XEL,WII,WIJ,WIK,WIL,UEA,UEB,UEC,UED, GEC, UEH, IZZ); 
ram_16x4 rinst_54(YEI,YEJ,YEK,YEL,WMI,WMJ,WMK,WML,UEA,UEB,UEC,UED, GED, UEH, IZZ); 
ram_16x4 rinst_55(YFA,YFB,YFC,YFD,WNA,WNB,WNC,WND,ufa,ufb,ufc,ufd, GFD, UFG, IZZ); 
ram_16x4 rinst_56(XFI,XFJ,XFK,XFL,WJI,WJJ,WJK,WJL,UFA,UFB,UFC,UFD, GFC, UFH, IZZ); 
ram_16x4 rinst_57(YFI,YFJ,YFK,YFL,WNI,WNJ,WNK,WNL,UFA,UFB,UFC,UFD, GFD, UFH, IZZ); 
ram_16x4 rinst_58(XGA,XGB,XGC,XGD,WKA,WKB,WKC,WKD,uga,ugb,ugc,ugd, GGC, UGG, IZZ); 
ram_16x4 rinst_59(YGA,YGB,YGC,YGD,WOA,WOB,WOC,WOD,uga,ugb,ugc,ugd, GGD, UGG, IZZ); 
ram_16x4 rinst_60(YGI,YGJ,YGK,YGL,WOI,WOJ,WOK,WOL,UGA,UGB,UGC,UGD, GGD, UGH, IZZ); 
ram_16x4 rinst_61(XHA,XHB,XHC,XHD,WLA,WLB,WLC,WLD,uha,uhb,uhc,uhd, GHC, UHG, IZZ); 
ram_16x4 rinst_62(YHA,YHB,YHC,YHD,WPA,WPB,WPC,WPD,uha,uhb,uhc,uhd, GHD, UHG, IZZ); 
ram_16x4 rinst_63(YHI,YHJ,YHK,YHL,WPI,WPJ,WPK,WPL,UHA,UHB,UHC,UHD, GHD, UHH, IZZ); 
ram_16x4 rinst_64(RIA,RIB,RIC,RID,WAA,WAB,WAC,WAD,uia,uib,uic,uid, GIA, UIG, IZZ); 
ram_16x4 rinst_65(SIA,SIB,SIC,SID,WEA,WEB,WEC,WED,uia,uib,uic,uid, GIB, UIG, IZZ); 
ram_16x4 rinst_66(XIA,XIB,XIC,XID,WIA,WIB,WIC,WID,uia,uib,uic,uid, GIC, UIG, IZZ); 
ram_16x4 rinst_67(RII,RIJ,RIK,RIL,WAI,WAJ,WAK,WAL,UIA,UIB,UIC,UID, GIA, UIH, IZZ); 
ram_16x4 rinst_68(SII,SIJ,SIK,SIL,WEI,WEJ,WEK,WEL,UIA,UIB,UIC,UID, GIB, UIH, IZZ); 
ram_16x4 rinst_69(RJA,RJB,RJC,RJD,WBA,WBB,WBC,WBD,uja,ujb,ujc,ujd, GJA, UJG, IZZ); 
ram_16x4 rinst_70(SJA,SJB,SJC,SJD,WFA,WFB,WFC,WFD,uja,ujb,ujc,ujd, GJB, UJG, IZZ); 
ram_16x4 rinst_71(XJA,XJB,XJC,XJD,WJA,WJB,WJC,WJD,uja,ujb,ujc,ujd, GJC, UJG, IZZ); 
ram_16x4 rinst_72(RJI,RJJ,RJK,RJL,WBI,WBJ,WBK,WBL,UJA,UJB,UJC,UJD, GJA, UJH, IZZ); 
ram_16x4 rinst_73(SJI,SJJ,SJK,SJL,WFI,WFJ,WFK,WFL,UJA,UJB,UJC,UJD, GJB, UJH, IZZ); 
ram_16x4 rinst_74(RKA,RKB,RKC,RKD,WCA,WCB,WCC,WCD,uka,ukb,ukc,ukd, GKA, UKG, IZZ); 
ram_16x4 rinst_75(SKA,SKB,SKC,SKD,WGA,WGB,WGC,WGD,uka,ukb,ukc,ukd, GKB, UKG, IZZ); 
ram_16x4 rinst_76(RKI,RKJ,RKK,RKL,WCI,WCJ,WCK,WCL,UKA,UKB,UKC,UKD, GKA, UKH, IZZ); 
ram_16x4 rinst_77(SKI,SKJ,SKK,SKL,WGI,WGJ,WGK,WGL,UKA,UKB,UKC,UKD, GKB, UKH, IZZ); 
ram_16x4 rinst_78(XKI,XKJ,XKK,XKL,WKI,WKJ,WKK,WKL,UKA,UKB,UKC,UKD, GKC, UKH, IZZ); 
ram_16x4 rinst_79(RLA,RLB,RLC,RLD,WDA,WDB,WDC,WDD,ula,ulb,ulc,uld, GLA, ULG, IZZ); 
ram_16x4 rinst_80(SLA,SLB,SLC,SLD,WHA,WHB,WHC,WHD,ula,ulb,ulc,uld, GLB, ULG, IZZ); 
ram_16x4 rinst_81(RLI,RLJ,RLK,RLL,WDI,WDJ,WDK,WDL,ULA,ULB,ULC,ULD, GLA, ULH, IZZ); 
ram_16x4 rinst_82(SLI,SLJ,SLK,SLL,WHI,WHJ,WHK,WHL,ULA,ULB,ULC,ULD, GLB, ULH, IZZ); 
ram_16x4 rinst_83(XLI,XLJ,XLK,XLL,WLI,WLJ,WLK,WLL,ULA,ULB,ULC,ULD, GLC, ULH, IZZ); 
ram_16x4 rinst_84(YIA,YIB,YIC,YID,WMA,WMB,WMC,WMD,uia,uib,uic,uid, GID, UIG, IZZ); 
ram_16x4 rinst_85(XII,XIJ,XIK,XIL,WII,WIJ,WIK,WIL,UIA,UIB,UIC,UID, GIC, UIH, IZZ); 
ram_16x4 rinst_86(YII,YIJ,YIK,YIL,WMI,WMJ,WMK,WML,UIA,UIB,UIC,UID, GID, UIH, IZZ); 
ram_16x4 rinst_87(YJA,YJB,YJC,YJD,WNA,WNB,WNC,WND,uja,ujb,ujc,ujd, GJD, UJG, IZZ); 
ram_16x4 rinst_88(XJI,XJJ,XJK,XJL,WJI,WJJ,WJK,WJL,UJA,UJB,UJC,UJD, GJC, UJH, IZZ); 
ram_16x4 rinst_89(YJI,YJJ,YJK,YJL,WNI,WNJ,WNK,WNL,UJA,UJB,UJC,UJD, GJD, UJH, IZZ); 
ram_16x4 rinst_90(XKA,XKB,XKC,XKD,WKA,WKB,WKC,WKD,uka,ukb,ukc,ukd, GKC, UKG, IZZ); 
ram_16x4 rinst_91(YKA,YKB,YKC,YKD,WOA,WOB,WOC,WOD,uka,ukb,ukc,ukd, GKD, UKG, IZZ); 
ram_16x4 rinst_92(YKI,YKJ,YKK,YKL,WOI,WOJ,WOK,WOL,UKA,UKB,UKC,UKD, GKD, UKH, IZZ); 
ram_16x4 rinst_93(XLA,XLB,XLC,XLD,WLA,WLB,WLC,WLD,ula,ulb,ulc,uld, GLC, ULG, IZZ); 
ram_16x4 rinst_94(YLA,YLB,YLC,YLD,WPA,WPB,WPC,WPD,ula,ulb,ulc,uld, GLD, ULG, IZZ); 
ram_16x4 rinst_95(YLI,YLJ,YLK,YLL,WPI,WPJ,WPK,WPL,ULA,ULB,ULC,ULD, GLD, ULH, IZZ); 
ram_16x4 rinst_96(RMA,RMB,RMC,RMD,WAA,WAB,WAC,WAD,uma,umb,umc,umd, GMA, UMG, IZZ); 
ram_16x4 rinst_97(SMA,SMB,SMC,SMD,WEA,WEB,WEC,WED,uma,umb,umc,umd, GMB, UMG, IZZ); 
ram_16x4 rinst_98(XMA,XMB,XMC,XMD,WIA,WIB,WIC,WID,uma,umb,umc,umd, GMC, UMG, IZZ); 
ram_16x4 rinst_99(RMI,RMJ,RMK,RML,WAI,WAJ,WAK,WAL,UMA,UMB,UMC,UMD, GMA, UMH, IZZ); 
ram_16x4 rinst_100(SMI,SMJ,SMK,SML,WEI,WEJ,WEK,WEL,UMA,UMB,UMC,UMD, GMB, UMH, IZZ); 
ram_16x4 rinst_101(RNA,RNB,RNC,RND,WBA,WBB,WBC,WBD,una,unb,unc,und, GNA, UNG, IZZ); 
ram_16x4 rinst_102(SNA,SNB,SNC,SND,WFA,WFB,WFC,WFD,una,unb,unc,und, GNB, UNG, IZZ); 
ram_16x4 rinst_103(XNA,XNB,XNC,XND,WJA,WJB,WJC,WJD,una,unb,unc,und, GNC, UNG, IZZ); 
ram_16x4 rinst_104(RNI,RNJ,RNK,RNL,WBI,WBJ,WBK,WBL,UNA,UNB,UNC,UND, GNA, UNH, IZZ); 
ram_16x4 rinst_105(SNI,SNJ,SNK,SNL,WFI,WFJ,WFK,WFL,UNA,UNB,UNC,UND, GNB, UNH, IZZ); 
ram_16x4 rinst_106(ROA,ROB,ROC,ROD,WCA,WCB,WCC,WCD,uoa,uob,uoc,uod, GOA, UOG, IZZ); 
ram_16x4 rinst_107(SOA,SOB,SOC,SOD,WGA,WGB,WGC,WGD,uoa,uob,uoc,uod, GOB, UOG, IZZ); 
ram_16x4 rinst_108(ROI,ROJ,ROK,ROL,WCI,WCJ,WCK,WCL,UOA,UOB,UOC,UOD, GOA, UOH, IZZ); 
ram_16x4 rinst_109(SOI,SOJ,SOK,SOL,WGI,WGJ,WGK,WGL,UOA,UOB,UOC,UOD, GOB, UOH, IZZ); 
ram_16x4 rinst_110(XOI,XOJ,XOK,XOL,WKI,WKJ,WKK,WKL,UOA,UOB,UOC,UOD, GOC, UOH, IZZ); 
ram_16x4 rinst_111(RPA,RPB,RPC,RPD,WDA,WDB,WDC,WDD,upa,upb,upc,upd, GPA, UPG, IZZ); 
ram_16x4 rinst_112(SPA,SPB,SPC,SPD,WHA,WHB,WHC,WHD,upa,upb,upc,upd, GPB, UPG, IZZ); 
ram_16x4 rinst_113(RPI,RPJ,RPK,RPL,WDI,WDJ,WDK,WDL,UPA,UPB,UPC,UPD, GPA, UPH, IZZ); 
ram_16x4 rinst_114(SPI,SPJ,SPK,SPL,WHI,WHJ,WHK,WHL,UPA,UPB,UPC,UPD, GPB, UPH, IZZ); 
ram_16x4 rinst_115(XPI,XPJ,XPK,XPL,WLI,WLJ,WLK,WLL,UPA,UPB,UPC,UPD, GPC, UPH, IZZ); 
ram_16x4 rinst_116(YMA,YMB,YMC,YMD,WMA,WMB,WMC,WMD,uma,umb,umc,umd, GMD, UMG, IZZ); 
ram_16x4 rinst_117(XMI,XMJ,XMK,XML,WII,WIJ,WIK,WIL,UMA,UMB,UMC,UMD, GMC, UMH, IZZ); 
ram_16x4 rinst_118(YMI,YMJ,YMK,YML,WMI,WMJ,WMK,WML,UMA,UMB,UMC,UMD, GMD, UMH, IZZ); 
ram_16x4 rinst_119(YNA,YNB,YNC,YND,WNA,WNB,WNC,WND,una,unb,unc,und, GND, UNG, IZZ); 
ram_16x4 rinst_120(XNI,XNJ,XNK,XNL,WJI,WJJ,WJK,WJL,UNA,UNB,UNC,UND, GNC, UNH, IZZ); 
ram_16x4 rinst_121(YNI,YNJ,YNK,YNL,WNI,WNJ,WNK,WNL,UNA,UNB,UNC,UND, GND, UNH, IZZ); 
ram_16x4 rinst_122(XOA,XOB,XOC,XOD,WKA,WKB,WKC,WKD,uoa,uob,uoc,uod, GOC, UOG, IZZ); 
ram_16x4 rinst_123(YOA,YOB,YOC,YOD,WOA,WOB,WOC,WOD,uoa,uob,uoc,uod, GOD, UOG, IZZ); 
ram_16x4 rinst_124(YOI,YOJ,YOK,YOL,WOI,WOJ,WOK,WOL,UOA,UOB,UOC,UOD, GOD, UOH, IZZ); 
ram_16x4 rinst_125(XPA,XPB,XPC,XPD,WLA,WLB,WLC,WLD,upa,upb,upc,upd, GPC, UPG, IZZ); 
ram_16x4 rinst_126(YPA,YPB,YPC,YPD,WPA,WPB,WPC,WPD,upa,upb,upc,upd, GPD, UPG, IZZ); 
ram_16x4 rinst_127(YPI,YPJ,YPK,YPL,WPI,WPJ,WPK,WPL,UPA,UPB,UPC,UPD, GPD, UPH, IZZ); 
ram_16x4 rinst_128(RAE,RAF,RAG,RAH,WAE,WAF,WAG,WAH,uai,uaj,uak,ual, GAE, UAO, IZZ); 
ram_16x4 rinst_129(SAE,SAF,SAG,SAH,WEE,WEF,WEG,WEH,uai,uaj,uak,ual, GAF, UAO, IZZ); 
ram_16x4 rinst_130(XAE,XAF,XAG,XAH,WIE,WIF,WIG,WIH,uai,uaj,uak,ual, GAG, UAO, IZZ); 
ram_16x4 rinst_131(RAM,RAN,RAO,RAP,WAM,WAN,WAO,WAP,UAI,UAJ,UAK,UAL, GAE, UAP, IZZ); 
ram_16x4 rinst_132(SAM,SAN,SAO,SAP,WEM,WEN,WEO,WEP,UAI,UAJ,UAK,UAL, GAF, UAP, IZZ); 
ram_16x4 rinst_133(RBE,RBF,RBG,RBH,WBE,WBF,WBG,WBH,ubi,ubj,ubk,ubl, GBE, UBO, IZZ); 
ram_16x4 rinst_134(SBE,SBF,SBG,SBH,WFE,WFF,WFG,WFH,ubi,ubj,ubk,ubl, GBF, UBO, IZZ); 
ram_16x4 rinst_135(XBE,XBF,XBG,XBH,WJE,WJF,WJG,WJH,ubi,ubj,ubk,ubl, GBG, UBO, IZZ); 
ram_16x4 rinst_136(RBM,RBN,RBO,RBP,WBM,WBN,WBO,WBP,UBI,UBJ,UBK,UBL, GBE, UBP, IZZ); 
ram_16x4 rinst_137(SBM,SBN,SBO,SBP,WFM,WFN,WFO,WFP,UBI,UBJ,UBK,UBL, GBF, UBP, IZZ); 
ram_16x4 rinst_138(RCE,RCF,RCG,RCH,WCE,WCF,WCG,WCH,uci,ucj,uck,ucl, GCE, UCO, IZZ); 
ram_16x4 rinst_139(SCE,SCF,SCG,SCH,WGE,WGF,WGG,WGH,uci,ucj,uck,ucl, GCF, UCO, IZZ); 
ram_16x4 rinst_140(RCM,RCN,RCO,RCP,WCM,WCN,WCO,WCP,UCI,UCJ,UCK,UCL, GCE, UCP, IZZ); 
ram_16x4 rinst_141(SCM,SCN,SCO,SCP,WGM,WGN,WGO,WGP,UCI,UCJ,UCK,UCL, GCF, UCP, IZZ); 
ram_16x4 rinst_142(XCM,XCN,XCO,XCP,WKM,WKN,WKO,WKP,UCI,UCJ,UCK,UCL, GCG, UCP, IZZ); 
ram_16x4 rinst_143(RDE,RDF,RDG,RDH,WDE,WDF,WDG,WDH,udi,udj,udk,udl, GDE, UDO, IZZ); 
ram_16x4 rinst_144(SDE,SDF,SDG,SDH,WHE,WHF,WHG,WHH,udi,udj,udk,udl, GDF, UDO, IZZ); 
ram_16x4 rinst_145(RDM,RDN,RDO,RDP,WDM,WDN,WDO,WDP,UDI,UDJ,UDK,UDL, GDE, UDP, IZZ); 
ram_16x4 rinst_146(SDM,SDN,SDO,SDP,WHM,WHN,WHO,WHP,UDI,UDJ,UDK,UDL, GDF, UDP, IZZ); 
ram_16x4 rinst_147(XDM,XDN,XDO,XDP,WLM,WLN,WLO,WLP,UDI,UDJ,UDK,UDL, GDG, UDP, IZZ); 
ram_16x4 rinst_148(YAE,YAF,YAG,YAH,WME,WMF,WMG,WMH,uai,uaj,uak,ual, GAH, UAO, IZZ); 
ram_16x4 rinst_149(XAM,XAN,XAO,XAP,WIM,WIN,WIO,WIP,UAI,UAJ,UAK,UAL, GAG, UAP, IZZ); 
ram_16x4 rinst_150(YAM,YAN,YAO,YAP,WMM,WMN,WMO,WMP,UAI,UAJ,UAK,UAL, GAH, UAP, IZZ); 
ram_16x4 rinst_151(YBE,YBF,YBG,YBH,WNE,WNF,WNG,WNH,ubi,ubj,ubk,ubl, GBH, UBO, IZZ); 
ram_16x4 rinst_152(XBM,XBN,XBO,XBP,WJM,WJN,WJO,WJP,UBI,UBJ,UBK,UBL, GBG, UBP, IZZ); 
ram_16x4 rinst_153(YBM,YBN,YBO,YBP,WNM,WNN,WNO,WNP,UBI,UBJ,UBK,UBL, GBH, UBP, IZZ); 
ram_16x4 rinst_154(XCE,XCF,XCG,XCH,WKE,WKF,WKG,WKH,uci,ucj,uck,ucl, GCG, UCO, IZZ); 
ram_16x4 rinst_155(YCE,YCF,YCG,YCH,WOE,WOF,WOG,WOH,uci,ucj,uck,ucl, GCH, UCO, IZZ); 
ram_16x4 rinst_156(YCM,YCN,YCO,YCP,WOM,WON,WOO,WOP,UCI,UCJ,UCK,UCL, GCH, UCP, IZZ); 
ram_16x4 rinst_157(XDE,XDF,XDG,XDH,WLE,WLF,WLG,WLH,udi,udj,udk,udl, GDG, UDO, IZZ); 
ram_16x4 rinst_158(YDE,YDF,YDG,YDH,WPE,WPF,WPG,WPH,udi,udj,udk,udl, GDH, UDO, IZZ); 
ram_16x4 rinst_159(YDM,YDN,YDO,YDP,WPM,WPN,WPO,WPP,UDI,UDJ,UDK,UDL, GDH, UDP, IZZ); 
ram_16x4 rinst_160(REE,REFF ,REG,REH,WAE,WAF,WAG,WAH,uei,uej,uek,uel, GEE, UEO, IZZ); 
ram_16x4 rinst_161(SEE,SEF,SEG,SEH,WEE,WEF,WEG,WEH,uei,uej,uek,uel, GEF, UEO, IZZ); 
ram_16x4 rinst_162(XEE,XEF,XEG,XEH,WIE,WIF,WIG,WIH,uei,uej,uek,uel, GEG, UEO, IZZ); 
ram_16x4 rinst_163(REM,REN,REO,REP,WAM,WAN,WAO,WAP,UEI,UEJ,UEK,UEL, GEE, UEP, IZZ); 
ram_16x4 rinst_164(SEM,SEN,SEO,SEP,WEM,WEN,WEO,WEP,UEI,UEJ,UEK,UEL, GEF, UEP, IZZ); 
ram_16x4 rinst_165(RFE,RFF,RFG,RFH,WBE,WBF,WBG,WBH,ufi,ufj,ufk,ufl, GFE, UFO, IZZ); 
ram_16x4 rinst_166(SFE,SFF,SFG,SFH,WFE,WFF,WFG,WFH,ufi,ufj,ufk,ufl, GFF, UFO, IZZ); 
ram_16x4 rinst_167(XFE,XFF,XFG,XFH,WJE,WJF,WJG,WJH,ufi,ufj,ufk,ufl, GFG, UFO, IZZ); 
ram_16x4 rinst_168(RFM,RFN,RFO,RFP,WBM,WBN,WBO,WBP,UFI,UFJ,UFK,UFL, GFE, UFP, IZZ); 
ram_16x4 rinst_169(SFM,SFN,SFO,SFP,WFM,WFN,WFO,WFP,UFI,UFJ,UFK,UFL, GFF, UFP, IZZ); 
ram_16x4 rinst_170(RGE,RGF,RGG,RGH,WCE,WCF,WCG,WCH,ugi,ugj,ugk,ugl, GGE, UGO, IZZ); 
ram_16x4 rinst_171(SGE,SGF,SGG,SGH,WGE,WGF,WGG,WGH,ugi,ugj,ugk,ugl, GGF, UGO, IZZ); 
ram_16x4 rinst_172(RGM,RGN,RGO,RGP,WCM,WCN,WCO,WCP,UGI,UGJ,UGK,UGL, GGE, UGP, IZZ); 
ram_16x4 rinst_173(SGM,SGN,SGO,SGP,WGM,WGN,WGO,WGP,UGI,UGJ,UGK,UGL, GGF, UGP, IZZ); 
ram_16x4 rinst_174(XGM,XGN,XGO,XGP,WKM,WKN,WKO,WKP,UGI,UGJ,UGK,UGL, GGG, UGP, IZZ); 
ram_16x4 rinst_175(RHE,RHF,RHG,RHH,WDE,WDF,WDG,WDH,uhi,uhj,uhk,uhl, GHE, UHO, IZZ); 
ram_16x4 rinst_176(SHE,SHF,SHG,SHH,WHE,WHF,WHG,WHH,uhi,uhj,uhk,uhl, GHF, UHO, IZZ); 
ram_16x4 rinst_177(RHM,RHN,RHO,RHP,WDM,WDN,WDO,WDP,UHI,UHJ,UHK,UHL, GHE, UHP, IZZ); 
ram_16x4 rinst_178(SHM,SHN,SHO,SHP,WHM,WHN,WHO,WHP,UHI,UHJ,UHK,UHL, GHF, UHP, IZZ); 
ram_16x4 rinst_179(XHM,XHN,XHO,XHP,WLM,WLN,WLO,WLP,UHI,UHJ,UHK,UHL, GHG, UHP, IZZ); 
ram_16x4 rinst_180(YEE,YEF,YEG,YEH,WME,WMF,WMG,WMH,uei,uej,uek,uel, GEH, UEO, IZZ); 
ram_16x4 rinst_181(XEM,XEN,XEO,XEP,WIM,WIN,WIO,WIP,UEI,UEJ,UEK,UEL, GEG, UEP, IZZ); 
ram_16x4 rinst_182(YEM,YEN,YEO,YEP,WMM,WMN,WMO,WMP,UEI,UEJ,UEK,UEL, GEH, UEP, IZZ); 
ram_16x4 rinst_183(YFE,YFF,YFG,YFH,WNE,WNF,WNG,WNH,ufi,ufj,ufk,ufl, GFH, UFO, IZZ); 
ram_16x4 rinst_184(XFM,XFN,XFO,XFP,WJM,WJN,WJO,WJP,UFI,UFJ,UFK,UFL, GFG, UFP, IZZ); 
ram_16x4 rinst_185(YFM,YFN,YFO,YFP,WNM,WNN,WNO,WNP,UFI,UFJ,UFK,UFL, GFH, UFP, IZZ); 
ram_16x4 rinst_186(XGE,XGF,XGG,XGH,WKE,WKF,WKG,WKH,ugi,ugj,ugk,ugl, GGG, UGO, IZZ); 
ram_16x4 rinst_187(YGE,YGF,YGG,YGH,WOE,WOF,WOG,WOH,ugi,ugj,ugk,ugl, GGH, UGO, IZZ); 
ram_16x4 rinst_188(YGM,YGN,YGO,YGP,WOM,WON,WOO,WOP,UGI,UGJ,UGK,UGL, GGH, UGP, IZZ); 
ram_16x4 rinst_189(XHE,XHF,XHG,XHH,WLE,WLF,WLG,WLH,uhi,uhj,uhk,uhl, GHG, UHO, IZZ); 
ram_16x4 rinst_190(YHE,YHF,YHG,YHH,WPE,WPF,WPG,WPH,uhi,uhj,uhk,uhl, GHH, UHO, IZZ); 
ram_16x4 rinst_191(YHM,YHN,YHO,YHP,WPM,WPN,WPO,WPP,UHI,UHJ,UHK,UHL, GHH, UHP, IZZ); 
ram_16x4 rinst_192(RIE,RIF,RIG,RIH,WAE,WAF,WAG,WAH,uii,uij,uik,uil, GIE, UIO, IZZ); 
ram_16x4 rinst_193(SIE,SIF,SIG,SIH,WEE,WEF,WEG,WEH,uii,uij,uik,uil, GIF, UIO, IZZ); 
ram_16x4 rinst_194(XIE,XIF,XIG,XIH,WIE,WIF,WIG,WIH,uii,uij,uik,uil, GIG, UIO, IZZ); 
ram_16x4 rinst_195(RIM,RIN,RIO,RIP,WAM,WAN,WAO,WAP,UII,UIJ,UIK,UIL, GIE, UIP, IZZ); 
ram_16x4 rinst_196(SIM,SIN,SIO,SIP,WEM,WEN,WEO,WEP,UII,UIJ,UIK,UIL, GIF, UIP, IZZ); 
ram_16x4 rinst_197(RJE,RJF,RJG,RJH,WBE,WBF,WBG,WBH,uji,ujj,ujk,ujl, GJE, UJO, IZZ); 
ram_16x4 rinst_198(SJE,SJF,SJG,SJH,WFE,WFF,WFG,WFH,uji,ujj,ujk,ujl, GJF, UJO, IZZ); 
ram_16x4 rinst_199(XJE,XJF,XJG,XJH,WJE,WJF,WJG,WJH,uji,ujj,ujk,ujl, GJG, UJO, IZZ); 
ram_16x4 rinst_200(RJM,RJN,RJO,RJP,WBM,WBN,WBO,WBP,UJI,UJJ,UJK,UJL, GJE, UJP, IZZ); 
ram_16x4 rinst_201(SJM,SJN,SJO,SJP,WFM,WFN,WFO,WFP,UJI,UJJ,UJK,UJL, GJF, UJP, IZZ); 
ram_16x4 rinst_202(RKE,RKF,RKG,RKH,WCE,WCF,WCG,WCH,uki,ukj,ukk,ukl, GKE, UKO, IZZ); 
ram_16x4 rinst_203(SKE,SKF,SKG,SKH,WGE,WGF,WGG,WGH,uki,ukj,ukk,ukl, GKF, UKO, IZZ); 
ram_16x4 rinst_204(RKM,RKN,RKO,RKP,WCM,WCN,WCO,WCP,UKI,UKJ,UKK,UKL, GKE, UKP, IZZ); 
ram_16x4 rinst_205(SKM,SKN,SKO,SKP,WGM,WGN,WGO,WGP,UKI,UKJ,UKK,UKL, GKF, UKP, IZZ); 
ram_16x4 rinst_206(XKM,XKN,XKO,XKP,WKM,WKN,WKO,WKP,UKI,UKJ,UKK,UKL, GKG, UKP, IZZ); 
ram_16x4 rinst_207(RLE,RLF,RLG,RLH,WDE,WDF,WDG,WDH,uli,ulj,ulk,ull, GLE, ULO, IZZ); 
ram_16x4 rinst_208(SLE,SLF,SLG,SLH,WHE,WHF,WHG,WHH,uli,ulj,ulk,ull, GLF, ULO, IZZ); 
ram_16x4 rinst_209(RLM,RLN,RLO,RLP,WDM,WDN,WDO,WDP,ULI,ULJ,ULK,ULL, GLE, ULP, IZZ); 
ram_16x4 rinst_210(SLM,SLN,SLO,SLP,WHM,WHN,WHO,WHP,ULI,ULJ,ULK,ULL, GLF, ULP, IZZ); 
ram_16x4 rinst_211(XLM,XLN,XLO,XLP,WLM,WLN,WLO,WLP,ULI,ULJ,ULK,ULL, GLG, ULP, IZZ); 
ram_16x4 rinst_212(YIE,YIF,YIG,YIH,WME,WMF,WMG,WMH,uii,uij,uik,uil, GIH, UIO, IZZ); 
ram_16x4 rinst_213(XIM,XIN,XIO,XIP,WIM,WIN,WIO,WIP,UII,UIJ,UIK,UIL, GIG, UIP, IZZ); 
ram_16x4 rinst_214(YIM,YIN,YIO,YIP,WMM,WMN,WMO,WMP,UII,UIJ,UIK,UIL, GIH, UIP, IZZ); 
ram_16x4 rinst_215(YJE,YJF,YJG,YJH,WNE,WNF,WNG,WNH,uji,ujj,ujk,ujl, GJH, UJO, IZZ); 
ram_16x4 rinst_216(XJM,XJN,XJO,XJP,WJM,WJN,WJO,WJP,UJI,UJJ,UJK,UJL, GJG, UJP, IZZ); 
ram_16x4 rinst_217(YJM,YJN,YJO,YJP,WNM,WNN,WNO,WNP,UJI,UJJ,UJK,UJL, GJH, UJP, IZZ); 
ram_16x4 rinst_218(XKE,XKF,XKG,XKH,WKE,WKF,WKG,WKH,uki,ukj,ukk,ukl, GKG, UKO, IZZ); 
ram_16x4 rinst_219(YKE,YKF,YKG,YKH,WOE,WOF,WOG,WOH,uki,ukj,ukk,ukl, GKH, UKO, IZZ); 
ram_16x4 rinst_220(YKM,YKN,YKO,YKP,WOM,WON,WOO,WOP,UKI,UKJ,UKK,UKL, GKH, UKP, IZZ); 
ram_16x4 rinst_221(XLE,XLF,XLG,XLH,WLE,WLF,WLG,WLH,uli,ulj,ulk,ull, GLG, ULO, IZZ); 
ram_16x4 rinst_222(YLE,YLF,YLG,YLH,WPE,WPF,WPG,WPH,uli,ulj,ulk,ull, GLH, ULO, IZZ); 
ram_16x4 rinst_223(YLM,YLN,YLO,YLP,WPM,WPN,WPO,WPP,ULI,ULJ,ULK,ULL, GLH, ULP, IZZ); 
ram_16x4 rinst_224(RME,RMF,RMG,RMH,WAE,WAF,WAG,WAH,umi,umj,umk,uml, GME, UMO, IZZ); 
ram_16x4 rinst_225(SME,SMF,SMG,SMH,WEE,WEF,WEG,WEH,umi,umj,umk,uml, GMF, UMO, IZZ); 
ram_16x4 rinst_226(XME,XMF,XMG,XMH,WIE,WIF,WIG,WIH,umi,umj,umk,uml, GMG, UMO, IZZ); 
ram_16x4 rinst_227(RMM,RMN,RMO,RMP,WAM,WAN,WAO,WAP,UMI,UMJ,UMK,UML, GME, UMP, IZZ); 
ram_16x4 rinst_228(SMM,SMN,SMO,SMP,WEM,WEN,WEO,WEP,UMI,UMJ,UMK,UML, GMF, UMP, IZZ); 
ram_16x4 rinst_229(RNE,RNF,RNG,RNH,WBE,WBF,WBG,WBH,uni,unj,unk,unl, GNE, UNO, IZZ); 
ram_16x4 rinst_230(SNE,SNF,SNG,SNH,WFE,WFF,WFG,WFH,uni,unj,unk,unl, GNF, UNO, IZZ); 
ram_16x4 rinst_231(XNE,XNF,XNG,XNH,WJE,WJF,WJG,WJH,uni,unj,unk,unl, GNG, UNO, IZZ); 
ram_16x4 rinst_232(RNM,RNN,RNO,RNP,WBM,WBN,WBO,WBP,UNI,UNJ,UNK,UNL, GNE, UNP, IZZ); 
ram_16x4 rinst_233(SNM,SNN,SNO,SNP,WFM,WFN,WFO,WFP,UNI,UNJ,UNK,UNL, GNF, UNP, IZZ); 
ram_16x4 rinst_234(ROE,ROF,ROG,ROH,WCE,WCF,WCG,WCH,uoi,uoj,uok,uol, GOE, UOO, IZZ); 
ram_16x4 rinst_235(SOE,SOF,SOG,SOH,WGE,WGF,WGG,WGH,uoi,uoj,uok,uol, GOF, UOO, IZZ); 
ram_16x4 rinst_236(ROM,RON,ROO,ROP,WCM,WCN,WCO,WCP,UOI,UOJ,UOK,UOL, GOE, UOP, IZZ); 
ram_16x4 rinst_237(SOM,SON,SOO,SOP,WGM,WGN,WGO,WGP,UOI,UOJ,UOK,UOL, GOF, UOP, IZZ); 
ram_16x4 rinst_238(XOM,XON,XOO,XOP,WKM,WKN,WKO,WKP,UOI,UOJ,UOK,UOL, GOG, UOP, IZZ); 
ram_16x4 rinst_239(RPE,RPF,RPG,RPH,WDE,WDF,WDG,WDH,upi,upj,upk,upl, GPE, UPO, IZZ); 
ram_16x4 rinst_240(SPE,SPF,SPG,SPH,WHE,WHF,WHG,WHH,upi,upj,upk,upl, GPF, UPO, IZZ); 
ram_16x4 rinst_241(RPM,RPN,RPO,RPP,WDM,WDN,WDO,WDP,UPI,UPJ,UPK,UPL, GPE, UPP, IZZ); 
ram_16x4 rinst_242(SPM,SPN,SPO,SPP,WHM,WHN,WHO,WHP,UPI,UPJ,UPK,UPL, GPF, UPP, IZZ); 
ram_16x4 rinst_243(XPM,XPN,XPO,XPP,WLM,WLN,WLO,WLP,UPI,UPJ,UPK,UPL, GPG, UPP, IZZ); 
ram_16x4 rinst_244(YME,YMF,YMG,YMH,WME,WMF,WMG,WMH,umi,umj,umk,uml, GMH, UMO, IZZ); 
ram_16x4 rinst_245(XMM,XMN,XMO,XMP,WIM,WIN,WIO,WIP,UMI,UMJ,UMK,UML, GMG, UMP, IZZ); 
ram_16x4 rinst_246(YMM,YMN,YMO,YMP,WMM,WMN,WMO,WMP,UMI,UMJ,UMK,UML, GMH, UMP, IZZ); 
ram_16x4 rinst_247(YNE,YNF,YNG,YNH,WNE,WNF,WNG,WNH,uni,unj,unk,unl, GNH, UNO, IZZ); 
ram_16x4 rinst_248(XNM,XNN,XNO,XNP,WJM,WJN,WJO,WJP,UNI,UNJ,UNK,UNL, GNG, UNP, IZZ); 
ram_16x4 rinst_249(YNM,YNN,YNO,YNP,WNM,WNN,WNO,WNP,UNI,UNJ,UNK,UNL, GNH, UNP, IZZ); 
ram_16x4 rinst_250(XOE,XOF,XOG,XOH,WKE,WKF,WKG,WKH,uoi,uoj,uok,uol, GOG, UOO, IZZ); 
ram_16x4 rinst_251(YOE,YOF,YOG,YOH,WOE,WOF,WOG,WOH,uoi,uoj,uok,uol, GOH, UOO, IZZ); 
ram_16x4 rinst_252(YOM,YON,YOO,YOP,WOM,WON,WOO,WOP,UOI,UOJ,UOK,UOL, GOH, UOP, IZZ); 
ram_16x4 rinst_253(XPE,XPF,XPG,XPH,WLE,WLF,WLG,WLH,upi,upj,upk,upl, GPG, UPO, IZZ); 
ram_16x4 rinst_254(YPE,YPF,YPG,YPH,WPE,WPF,WPG,WPH,upi,upj,upk,upl, GPH, UPO, IZZ); 
ram_16x4 rinst_255(YPM,YPN,YPO,YPP,WPM,WPN,WPO,WPP,UPI,UPJ,UPK,UPL, GPH, UPP, IZZ); 
endmodule;
