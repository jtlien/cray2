module ia( IZZ,
 IAA, 
 IAB, 
 IAC, 
 IAD, 
 IAE, 
 IAF, 
 IAG, 
 IAH, 
 IAI, 
 IAJ, 
 IAK, 
 IAL, 
 IAM, 
 IAN, 
 IAO, 
 IAP, 
 IBA, 
 IBB, 
 IBC, 
 IBD, 
 IBE, 
 IBF, 
 IBG, 
 IBH, 
 IBI, 
 IBJ, 
 IBK, 
 IBL, 
 IBM, 
 IBN, 
 IBO, 
 IBP, 
 ICA, 
 ICB, 
 ICC, 
 ICD, 
 ICE, 
 ICF, 
 ICG, 
 ICH, 
 ICI, 
 ICJ, 
 ICK, 
 ICL, 
 ICM, 
 ICN, 
 ICO, 
 ICP, 
 IDA, 
 IDB, 
 IDC, 
 IDD, 
 IDE, 
 IDF, 
 IDG, 
 IDH, 
 IDI, 
 IDJ, 
 IDK, 
 IDL, 
 IDM, 
 IDN, 
 IDO, 
 IDP, 
 IEA, 
 IEB, 
 IEC, 
 IED, 
 IEE, 
 IEF, 
 IEG, 
 IEH, 
 IEI, 
 IEJ, 
 IEK, 
 IEL, 
 IEM, 
 IEN, 
 IEO, 
 IEP, 
 IEQ, 
 IER, 
 IES, 
 IET, 
 IEU, 
 IEV, 
 IEW, 
 IEX, 
 IFA, 
 IFB, 
 IFC, 
 IFD, 
 IGA, 
 IGB, 
 IGC, 
 IHA, 
 IHB, 
 IJB, 
 IJD, 
 IJE, 
 IJF, 
 OAA, 
 OAB, 
 OAC, 
 OAD, 
 OAE, 
 OAF, 
 OAG, 
 OAH, 
 OAI, 
 OAJ, 
 OAK, 
 OAL, 
 OAM, 
 OAN, 
 OAO, 
 OAP, 
 OAP, 
 OBA, 
 OBB, 
 OBC, 
 OBD, 
 OBE, 
 OBF, 
 OBG, 
 OBH, 
 OBI, 
 OBJ, 
 OBK, 
 OBL, 
 OBM, 
 OBN, 
 OBO, 
 OBP, 
 OCA, 
 OCB, 
 OCC, 
 OCD, 
 OCE, 
 OCF, 
 OCG, 
 OCH, 
 OCI, 
 OCJ, 
 OCK, 
 OCL, 
 OCM, 
 OCN, 
 OCO, 
 OCP, 
 ODA, 
 ODB, 
 ODC, 
 ODD, 
 ODE, 
 ODF, 
 ODG, 
 ODH, 
 ODI, 
 ODJ, 
 ODK, 
 ODL, 
 ODM, 
 ODN, 
 ODO, 
 ODP, 
 OEA, 
 OEB, 
 OEC, 
 OED, 
 OEE, 
 OEF, 
 OEG, 
 OEH, 
 OEI, 
 OEJ, 
 OEK, 
 OEL, 
 OEM, 
 OEN, 
 OEO, 
 OFA, 
 OFB, 
 OFC, 
 OFD, 
 OFE, 
 OFF, 
 OFG, 
 OFH, 
 OFI, 
 OFJ, 
 OFK, 
 OFL, 
 OFM, 
 OFN, 
 OFO, 
 OFP, 
 OGA, 
 OGB, 
 OGC, 
 OGD, 
 OGE, 
 OGF, 
 OGG, 
 OGH, 
 OGI, 
 OGJ, 
 OGK, 
 OGL, 
 OGM, 
 OGN, 
 OGO, 
 OGP, 
 OHA, 
 OHB, 
 OHC, 
 OHD, 
 OHE, 
 OHF, 
 OHG, 
 OHH, 
 OHI, 
 OHJ, 
 OHK, 
 OHL, 
 OHM, 
 OHN, 
 OHO, 
 OHP, 
 OJA, 
 OJB, 
 OJC, 
 OJD, 
 OJE, 
 OKA, 
 OKB, 
 OKC, 
 OKD, 
 OKE, 
 OKF, 
 OKG, 
 OKH, 
 OKI, 
 OKJ, 
 OKK, 
 OKL, 
 OKM, 
 OKN, 
 OKO, 
 OKP, 
 OKQ, 
 OKR, 
 OKS, 
 OKT, 
 OKU, 
 OKV, 
 OKW, 
OKX ); 
    
 input IZZ; 
 input IAA; 
 input IAB; 
 input IAC; 
 input IAD; 
 input IAE; 
 input IAF; 
 input IAG; 
 input IAH; 
 input IAI; 
 input IAJ; 
 input IAK; 
 input IAL; 
 input IAM; 
 input IAN; 
 input IAO; 
 input IAP; 
 input IBA; 
 input IBB; 
 input IBC; 
 input IBD; 
 input IBE; 
 input IBF; 
 input IBG; 
 input IBH; 
 input IBI; 
 input IBJ; 
 input IBK; 
 input IBL; 
 input IBM; 
 input IBN; 
 input IBO; 
 input IBP; 
 input ICA; 
 input ICB; 
 input ICC; 
 input ICD; 
 input ICE; 
 input ICF; 
 input ICG; 
 input ICH; 
 input ICI; 
 input ICJ; 
 input ICK; 
 input ICL; 
 input ICM; 
 input ICN; 
 input ICO; 
 input ICP; 
 input IDA; 
 input IDB; 
 input IDC; 
 input IDD; 
 input IDE; 
 input IDF; 
 input IDG; 
 input IDH; 
 input IDI; 
 input IDJ; 
 input IDK; 
 input IDL; 
 input IDM; 
 input IDN; 
 input IDO; 
 input IDP; 
 input IEA; 
 input IEB; 
 input IEC; 
 input IED; 
 input IEE; 
 input IEF; 
 input IEG; 
 input IEH; 
 input IEI; 
 input IEJ; 
 input IEK; 
 input IEL; 
 input IEM; 
 input IEN; 
 input IEO; 
 input IEP; 
 input IEQ; 
 input IER; 
 input IES; 
 input IET; 
 input IEU; 
 input IEV; 
 input IEW; 
 input IEX; 
 input IFA; 
 input IFB; 
 input IFC; 
 input IFD; 
 input IGA; 
 input IGB; 
 input IGC; 
 input IHA; 
 input IHB; 
 input IJB; 
 input IJD; 
 input IJE; 
 input IJF; 
 output OAA; 
 output OAB; 
 output OAC; 
 output OAD; 
 output OAE; 
 output OAF; 
 output OAG; 
 output OAH; 
 output OAI; 
 output OAJ; 
 output OAK; 
 output OAL; 
 output OAM; 
 output OAN; 
 output OAO; 
 output OAP; 
 output OAP; 
 output OBA; 
 output OBB; 
 output OBC; 
 output OBD; 
 output OBE; 
 output OBF; 
 output OBG; 
 output OBH; 
 output OBI; 
 output OBJ; 
 output OBK; 
 output OBL; 
 output OBM; 
 output OBN; 
 output OBO; 
 output OBP; 
 output OCA; 
 output OCB; 
 output OCC; 
 output OCD; 
 output OCE; 
 output OCF; 
 output OCG; 
 output OCH; 
 output OCI; 
 output OCJ; 
 output OCK; 
 output OCL; 
 output OCM; 
 output OCN; 
 output OCO; 
 output OCP; 
 output ODA; 
 output ODB; 
 output ODC; 
 output ODD; 
 output ODE; 
 output ODF; 
 output ODG; 
 output ODH; 
 output ODI; 
 output ODJ; 
 output ODK; 
 output ODL; 
 output ODM; 
 output ODN; 
 output ODO; 
 output ODP; 
 output OEA; 
 output OEB; 
 output OEC; 
 output OED; 
 output OEE; 
 output OEF; 
 output OEG; 
 output OEH; 
 output OEI; 
 output OEJ; 
 output OEK; 
 output OEL; 
 output OEM; 
 output OEN; 
 output OEO; 
 output OFA; 
 output OFB; 
 output OFC; 
 output OFD; 
 output OFE; 
 output OFF; 
 output OFG; 
 output OFH; 
 output OFI; 
 output OFJ; 
 output OFK; 
 output OFL; 
 output OFM; 
 output OFN; 
 output OFO; 
 output OFP; 
 output OGA; 
 output OGB; 
 output OGC; 
 output OGD; 
 output OGE; 
 output OGF; 
 output OGG; 
 output OGH; 
 output OGI; 
 output OGJ; 
 output OGK; 
 output OGL; 
 output OGM; 
 output OGN; 
 output OGO; 
 output OGP; 
 output OHA; 
 output OHB; 
 output OHC; 
 output OHD; 
 output OHE; 
 output OHF; 
 output OHG; 
 output OHH; 
 output OHI; 
 output OHJ; 
 output OHK; 
 output OHL; 
 output OHM; 
 output OHN; 
 output OHO; 
 output OHP; 
 output OJA; 
 output OJB; 
 output OJC; 
 output OJD; 
 output OJE; 
 output OKA; 
 output OKB; 
 output OKC; 
 output OKD; 
 output OKE; 
 output OKF; 
 output OKG; 
 output OKH; 
 output OKI; 
 output OKJ; 
 output OKK; 
 output OKL; 
 output OKM; 
 output OKN; 
 output OKO; 
 output OKP; 
 output OKQ; 
 output OKR; 
 output OKS; 
 output OKT; 
 output OKU; 
 output OKV; 
 output OKW; 
 output OKX; 
  
  
reg  AAA ;
reg  AAB ;
reg  AAC ;
reg  AAD ;
reg  AAE ;
reg  AAF ;
reg  AAG ;
reg  AAH ;
reg  AAI ;
reg  AAJ ;
reg  AAK ;
reg  AAL ;
reg  AAM ;
reg  AAN ;
reg  AAO ;
reg  AAP ;
reg  AAQ ;
reg  AAR ;
reg  AAS ;
reg  AAT ;
reg  AAU ;
reg  AAV ;
reg  AAW ;
reg  AAX ;
reg  ABA ;
reg  ABB ;
reg  ABC ;
reg  ABD ;
reg  ABE ;
reg  ABF ;
reg  ABG ;
reg  ABH ;
reg  ABI ;
reg  ABJ ;
reg  ABK ;
reg  ABL ;
reg  ABM ;
reg  ABN ;
reg  ABO ;
reg  ABP ;
reg  ABQ ;
reg  ABR ;
reg  ABS ;
reg  ABT ;
reg  ABU ;
reg  ABV ;
reg  ABW ;
reg  ABX ;
reg  ACA ;
reg  ACB ;
reg  ACC ;
reg  ACD ;
reg  ACE ;
reg  ACF ;
reg  ACG ;
reg  ACH ;
reg  ACI ;
reg  ACJ ;
reg  ACK ;
reg  ACL ;
reg  ACM ;
reg  ACN ;
reg  ACO ;
reg  ACP ;
reg  ACQ ;
reg  ACR ;
reg  ACS ;
reg  ACT ;
reg  ACU ;
reg  ACV ;
reg  ACW ;
reg  ACX ;
reg  ADA ;
reg  ADB ;
reg  ADC ;
reg  ADD ;
reg  ADE ;
reg  ADF ;
reg  ADG ;
reg  ADH ;
reg  ADI ;
reg  ADJ ;
reg  ADK ;
reg  ADL ;
reg  ADM ;
reg  ADN ;
reg  ADO ;
reg  ADP ;
reg  ADQ ;
reg  ADR ;
reg  ADS ;
reg  ADT ;
reg  ADU ;
reg  ADV ;
reg  ADW ;
reg  ADX ;
reg  AEA ;
reg  AEB ;
reg  AEC ;
reg  AED ;
reg  AEE ;
reg  AEF ;
reg  AEG ;
reg  AEH ;
reg  AEI ;
reg  AEJ ;
reg  AEK ;
reg  AEL ;
reg  AEM ;
reg  AEN ;
reg  AEO ;
reg  AEP ;
reg  AEQ ;
reg  AER ;
reg  AES ;
reg  AET ;
reg  AEU ;
reg  AEV ;
reg  AEW ;
reg  AEX ;
reg  AFA ;
reg  AFB ;
reg  AFC ;
reg  AFD ;
reg  AFE ;
reg  AFF ;
reg  AFG ;
reg  AFH ;
reg  AFI ;
reg  AFJ ;
reg  AFK ;
reg  AFL ;
reg  AFM ;
reg  AFN ;
reg  AFO ;
reg  AFP ;
reg  AFQ ;
reg  AFR ;
reg  AFS ;
reg  AFT ;
reg  AFU ;
reg  AFV ;
reg  AFW ;
reg  AFX ;
reg  AGA ;
reg  AGB ;
reg  AGC ;
reg  AGD ;
reg  AGE ;
reg  AGF ;
reg  AGG ;
reg  AGH ;
reg  AGI ;
reg  AGJ ;
reg  AGK ;
reg  AGL ;
reg  AGM ;
reg  AGN ;
reg  AGO ;
reg  AGP ;
reg  AGQ ;
reg  AGR ;
reg  AGS ;
reg  AGT ;
reg  AGU ;
reg  AGV ;
reg  AGW ;
reg  AGX ;
reg  AHA ;
reg  AHB ;
reg  AHC ;
reg  AHD ;
reg  AHE ;
reg  AHF ;
reg  AHG ;
reg  AHH ;
reg  AHI ;
reg  AHJ ;
reg  AHK ;
reg  AHL ;
reg  AHM ;
reg  AHN ;
reg  AHO ;
reg  AHP ;
reg  AHQ ;
reg  AHR ;
reg  AHS ;
reg  AHT ;
reg  AHU ;
reg  AHV ;
reg  AHW ;
reg  AHX ;
reg  AIA ;
reg  AIB ;
reg  AIC ;
reg  AID ;
reg  AIE ;
reg  AIF ;
reg  AIG ;
reg  AIH ;
reg  AII ;
reg  AIJ ;
reg  AIK ;
reg  AIL ;
reg  AIM ;
reg  AIN ;
reg  AIO ;
reg  AIP ;
reg  AIQ ;
reg  AIR ;
reg  AIS ;
reg  AIT ;
reg  AIU ;
reg  AIV ;
reg  AIW ;
reg  AIX ;
reg  CAA ;
reg  CAB ;
reg  CBA ;
reg  CBB ;
reg  CCA ;
reg  CCB ;
reg  CDA ;
reg  CDB ;
reg  DAA ;
reg  DAB ;
reg  DAC ;
reg  DAD ;
reg  DAE ;
reg  DAF ;
reg  DAG ;
reg  DAH ;
reg  DAI ;
reg  DAJ ;
reg  DAK ;
reg  DAL ;
reg  DBA ;
reg  DBB ;
reg  DBC ;
reg  DBE ;
reg  DBF ;
reg  DBG ;
reg  DBI ;
reg  DBJ ;
reg  DBK ;
reg  EAA ;
reg  EAB ;
reg  EAC ;
reg  EAD ;
reg  eba ;
reg  ebb ;
reg  ebc ;
reg  FAA ;
reg  FAB ;
reg  FAC ;
reg  FAD ;
reg  GAA ;
reg  GAB ;
reg  GAC ;
reg  HAA ;
reg  HAB ;
reg  HAC ;
reg  HBA ;
reg  HBB ;
reg  HBC ;
reg  HCA ;
reg  HCB ;
reg  HCC ;
reg  HDA ;
reg  HDB ;
reg  HDC ;
reg  HEA ;
reg  HEB ;
reg  HEC ;
reg  HFA ;
reg  HFB ;
reg  HFC ;
reg  HGA ;
reg  HGB ;
reg  HGC ;
reg  HHA ;
reg  HHB ;
reg  HHC ;
reg  HIA ;
reg  HIB ;
reg  HIC ;
reg  HID ;
reg  KDE ;
reg  OAA ;
reg  OAB ;
reg  OAC ;
reg  OAD ;
reg  OAE ;
reg  OAF ;
reg  OAG ;
reg  OAH ;
reg  OAI ;
reg  OAJ ;
reg  OAK ;
reg  OAL ;
reg  OAM ;
reg  OAN ;
reg  OAO ;
reg  OAP ;
reg  OBA ;
reg  OBB ;
reg  OBC ;
reg  OBD ;
reg  OBE ;
reg  OBF ;
reg  OBG ;
reg  OBH ;
reg  OBI ;
reg  OBJ ;
reg  OBK ;
reg  OBL ;
reg  OBM ;
reg  OBN ;
reg  OBO ;
reg  OBP ;
reg  OCA ;
reg  OCB ;
reg  OCC ;
reg  OCD ;
reg  OCE ;
reg  OCF ;
reg  OCG ;
reg  OCH ;
reg  OCI ;
reg  OCJ ;
reg  OCK ;
reg  OCL ;
reg  OCM ;
reg  OCN ;
reg  OCO ;
reg  OCP ;
reg  ODA ;
reg  ODB ;
reg  ODC ;
reg  ODD ;
reg  ODE ;
reg  ODF ;
reg  ODG ;
reg  ODH ;
reg  ODI ;
reg  ODJ ;
reg  ODK ;
reg  ODL ;
reg  ODM ;
reg  ODN ;
reg  ODO ;
reg  ODP ;
reg  oea ;
reg  oeb ;
reg  oec ;
reg  oed ;
reg  oee ;
reg  oef ;
reg  oeg ;
reg  oeh ;
reg  oei ;
reg  oej ;
reg  oek ;
reg  oel ;
reg  oem ;
reg  oen ;
reg  oeo ;
reg  oep ;
reg  ofa ;
reg  ofb ;
reg  ofc ;
reg  ofd ;
reg  ofe ;
reg  off ;
reg  ofg ;
reg  ofh ;
reg  ofi ;
reg  ofj ;
reg  ofk ;
reg  ofl ;
reg  ofm ;
reg  ofn ;
reg  ofo ;
reg  ofp ;
reg  oga ;
reg  ogb ;
reg  ogc ;
reg  ogd ;
reg  oge ;
reg  ogf ;
reg  ogg ;
reg  ogh ;
reg  ogi ;
reg  ogj ;
reg  ogk ;
reg  ogl ;
reg  ogm ;
reg  ogn ;
reg  ogo ;
reg  ogp ;
reg  oha ;
reg  ohb ;
reg  ohc ;
reg  ohd ;
reg  ohe ;
reg  ohf ;
reg  ohg ;
reg  ohh ;
reg  ohi ;
reg  ohj ;
reg  ohk ;
reg  ohl ;
reg  ohm ;
reg  ohn ;
reg  oho ;
reg  ohp ;
reg  OJA ;
reg  OJB ;
reg  OJC ;
reg  ojd ;
reg  oje ;
reg  OKA ;
reg  OKB ;
reg  OKC ;
reg  OKD ;
reg  OKE ;
reg  okf ;
reg  OKG ;
reg  OKH ;
reg  oki ;
reg  okj ;
reg  okk ;
reg  okl ;
reg  okm ;
reg  okn ;
reg  oko ;
reg  okp ;
reg  okq ;
reg  okr ;
reg  oks ;
reg  okt ;
reg  oku ;
reg  okv ;
reg  okw ;
reg  okx ;
reg  PAA ;
reg  PAB ;
reg  PAC ;
reg  PAD ;
reg  PAE ;
reg  PAF ;
reg  PBA ;
reg  PBB ;
reg  PBC ;
reg  PBD ;
reg  PBE ;
reg  PBF ;
reg  PCA ;
reg  PCB ;
reg  PCC ;
reg  PCD ;
reg  PCE ;
reg  PCF ;
reg  PDA ;
reg  PDB ;
reg  PDC ;
reg  PDD ;
reg  PDE ;
reg  PDF ;
reg  PEA ;
reg  PEB ;
reg  PEC ;
reg  PFA ;
reg  PFB ;
reg  PFC ;
reg  PGA ;
reg  PGB ;
reg  PGC ;
reg  qaa ;
reg  qab ;
reg  qac ;
reg  qad ;
reg  QAE ;
reg  QBA ;
reg  QBB ;
reg  QBC ;
reg  QBD ;
reg  QBE ;
reg  QCA ;
reg  QCB ;
reg  QCC ;
reg  QCD ;
reg  QCE ;
reg  QDA ;
reg  qdb ;
reg  QDC ;
reg  QDD ;
reg  QDE ;
reg  QDI ;
reg  QDJ ;
reg  QDK ;
reg  QDL ;
reg  QEB ;
reg  qec ;
reg  qed ;
reg  QFA ;
reg  qha ;
reg  qhb ;
reg  qhc ;
reg  qhd ;
reg  QJA ;
reg  QJB ;
reg  QJC ;
reg  QJD ;
reg  QJE ;
reg  QJF ;
reg  QJG ;
reg  QJH ;
reg  QJI ;
reg  QJJ ;
reg  QJK ;
reg  QJM ;
reg  QJN ;
reg  QJP ;
reg  QKA ;
reg  QKB ;
reg  qla ;
reg  qlb ;
reg  qlc ;
reg  QLD ;
reg  qle ;
reg  QLF ;
reg  QLG ;
reg  QLH ;
reg  QPA ;
reg  QPB ;
reg  QPC ;
reg  QPD ;
reg  QPE ;
reg  QQA ;
reg  QQB ;
reg  QQC ;
reg  QQD ;
reg  TAA ;
reg  TAB ;
reg  TAC ;
reg  TAD ;
reg  TAE ;
reg  TAF ;
reg  TAG ;
reg  TAH ;
reg  TBA ;
reg  TBB ;
reg  TBC ;
reg  TBD ;
reg  TBE ;
reg  TBF ;
reg  TBG ;
reg  TBH ;
reg  TCA ;
reg  TCB ;
reg  TCC ;
reg  TCD ;
reg  TCE ;
reg  TCF ;
reg  TCG ;
reg  TCH ;
reg  TDA ;
reg  TDB ;
reg  TDC ;
reg  TDD ;
reg  TDE ;
reg  TDF ;
reg  TDG ;
reg  TDH ;
reg  TEA ;
reg  TEB ;
reg  TEC ;
reg  TED ;
reg  TEE ;
reg  TEF ;
reg  TEG ;
reg  TEH ;
reg  TFA ;
reg  TFB ;
reg  TFC ;
reg  TFD ;
reg  tga ;
reg  tgb ;
reg  tgc ;
reg  tgd ;
reg  TJA ;
reg  TJB ;
reg  TJC ;
reg  TJD ;
reg  TMA ;
reg  UAA ;
reg  UAB ;
reg  UAC ;
reg  UAD ;
reg  UAE ;
reg  UAF ;
reg  UAG ;
reg  UAI ;
reg  UAJ ;
reg  UAK ;
reg  UAL ;
reg  UAM ;
reg  UAN ;
reg  UAO ;
reg  UBA ;
reg  UBB ;
reg  UBC ;
reg  UBD ;
reg  UBE ;
reg  UBF ;
reg  UBG ;
reg  UBI ;
reg  UBJ ;
reg  UBK ;
reg  UBL ;
reg  UBM ;
reg  UBN ;
reg  UBO ;
reg  UCA ;
reg  UCB ;
reg  UCC ;
reg  UCD ;
reg  UCE ;
reg  UCF ;
reg  UCG ;
reg  UCI ;
reg  UCJ ;
reg  UCK ;
reg  UCL ;
reg  UCM ;
reg  UCN ;
reg  UCO ;
reg  UDA ;
reg  UDB ;
reg  UDC ;
reg  UDD ;
reg  UDE ;
reg  UDF ;
reg  UDG ;
reg  UDI ;
reg  UDJ ;
reg  UDK ;
reg  UDL ;
reg  UDM ;
reg  UDN ;
reg  UDO ;
reg  UEA ;
reg  UEB ;
reg  UEC ;
reg  UED ;
reg  UEE ;
reg  UEF ;
reg  UEG ;
reg  UEI ;
reg  UEJ ;
reg  UEK ;
reg  UEL ;
reg  UEM ;
reg  UEN ;
reg  UEO ;
reg  UFA ;
reg  UFB ;
reg  UFC ;
reg  UFD ;
reg  UFE ;
reg  UFF ;
reg  UFG ;
reg  UFI ;
reg  UFJ ;
reg  UFK ;
reg  UFL ;
reg  UFM ;
reg  UFN ;
reg  UFO ;
reg  UGA ;
reg  UGB ;
reg  UGC ;
reg  UGD ;
reg  UGE ;
reg  UGF ;
reg  UGG ;
reg  UGI ;
reg  UGJ ;
reg  UGK ;
reg  UGL ;
reg  UGM ;
reg  UGN ;
reg  UGO ;
reg  UHA ;
reg  UHB ;
reg  UHC ;
reg  UHD ;
reg  UHE ;
reg  UHF ;
reg  UHG ;
reg  UHI ;
reg  UHJ ;
reg  UHK ;
reg  UHL ;
reg  UHM ;
reg  UHN ;
reg  UHO ;
reg  UIA ;
reg  UIB ;
reg  UIC ;
reg  UID ;
reg  UIE ;
reg  UIF ;
reg  UIG ;
reg  UII ;
reg  UIJ ;
reg  UIK ;
reg  UIL ;
reg  UIM ;
reg  UIN ;
reg  UIO ;
reg  UJA ;
reg  UJB ;
reg  UJC ;
reg  UJD ;
reg  UJE ;
reg  UJF ;
reg  UJG ;
reg  UJI ;
reg  UJJ ;
reg  UJK ;
reg  UJL ;
reg  UJM ;
reg  UJN ;
reg  UJO ;
reg  UKA ;
reg  UKB ;
reg  UKC ;
reg  UKD ;
reg  UKE ;
reg  UKF ;
reg  UKG ;
reg  UKI ;
reg  UKJ ;
reg  UKK ;
reg  UKL ;
reg  UKM ;
reg  UKN ;
reg  UKO ;
reg  ULA ;
reg  ULB ;
reg  ULC ;
reg  ULD ;
reg  ULE ;
reg  ULF ;
reg  ULG ;
reg  ULI ;
reg  ULJ ;
reg  ULK ;
reg  ULL ;
reg  ULM ;
reg  ULN ;
reg  ULO ;
reg  UMA ;
reg  UMB ;
reg  UMC ;
reg  UMD ;
reg  UME ;
reg  UMF ;
reg  UMG ;
reg  UMI ;
reg  UMJ ;
reg  UMK ;
reg  UML ;
reg  UMM ;
reg  UMN ;
reg  UMO ;
reg  UNA ;
reg  UNB ;
reg  UNC ;
reg  UND ;
reg  UNE ;
reg  UNF ;
reg  UNG ;
reg  UNI ;
reg  UNJ ;
reg  UNK ;
reg  UNL ;
reg  UNM ;
reg  UNN ;
reg  UNO ;
reg  UOA ;
reg  UOB ;
reg  UOC ;
reg  UOD ;
reg  UOE ;
reg  UOF ;
reg  UOG ;
reg  UOI ;
reg  UOJ ;
reg  UOK ;
reg  UOL ;
reg  UOM ;
reg  UON ;
reg  UOO ;
reg  UPA ;
reg  UPB ;
reg  UPC ;
reg  UPD ;
reg  UPE ;
reg  UPF ;
reg  UPG ;
reg  UPI ;
reg  UPJ ;
reg  UPK ;
reg  UPL ;
reg  UPM ;
reg  UPN ;
reg  UPO ;
reg  VAA ;
reg  VAB ;
reg  VAC ;
reg  VAD ;
reg  VAE ;
reg  VAF ;
reg  VAG ;
reg  VAH ;
reg  VAI ;
reg  VAJ ;
reg  VAK ;
reg  VAL ;
reg  VAM ;
reg  VAN ;
reg  VAO ;
reg  VAP ;
reg  VBA ;
reg  VBB ;
reg  VBC ;
reg  VBD ;
reg  VBE ;
reg  VBF ;
reg  VBG ;
reg  VBH ;
reg  VBI ;
reg  VBJ ;
reg  VBK ;
reg  VBL ;
reg  VBM ;
reg  VBN ;
reg  VBO ;
reg  VBP ;
reg  VCA ;
reg  VCB ;
reg  VCC ;
reg  VCD ;
reg  VCE ;
reg  VCF ;
reg  VCG ;
reg  VCH ;
reg  VCI ;
reg  VCJ ;
reg  VCK ;
reg  VCL ;
reg  VCM ;
reg  VCN ;
reg  VCO ;
reg  VCP ;
reg  VDA ;
reg  VDB ;
reg  VDC ;
reg  VDD ;
reg  VDE ;
reg  VDF ;
reg  VDG ;
reg  VDH ;
reg  VDI ;
reg  VDJ ;
reg  VDK ;
reg  VDL ;
reg  VDM ;
reg  VDN ;
reg  VDO ;
reg  VDP ;
reg  WAA ;
reg  WAB ;
reg  WAC ;
reg  WAD ;
reg  WAE ;
reg  WAF ;
reg  WAG ;
reg  WAH ;
reg  WAI ;
reg  WAJ ;
reg  WAK ;
reg  WAL ;
reg  WAM ;
reg  WAN ;
reg  WAO ;
reg  WAP ;
reg  WBA ;
reg  WBB ;
reg  WBC ;
reg  WBD ;
reg  WBE ;
reg  WBF ;
reg  WBG ;
reg  WBH ;
reg  WBI ;
reg  WBJ ;
reg  WBK ;
reg  WBL ;
reg  WBM ;
reg  WBN ;
reg  WBO ;
reg  WBP ;
reg  WCA ;
reg  WCB ;
reg  WCC ;
reg  WCD ;
reg  WCE ;
reg  WCF ;
reg  WCG ;
reg  WCH ;
reg  WCI ;
reg  WCJ ;
reg  WCK ;
reg  WCL ;
reg  WCM ;
reg  WCN ;
reg  WCO ;
reg  WCP ;
reg  WDA ;
reg  WDB ;
reg  WDC ;
reg  WDD ;
reg  WDE ;
reg  WDF ;
reg  WDG ;
reg  WDH ;
reg  WDI ;
reg  WDJ ;
reg  WDK ;
reg  WDL ;
reg  WDM ;
reg  WDN ;
reg  WDO ;
reg  WDP ;
reg  WEA ;
reg  WEB ;
reg  WEC ;
reg  WED ;
reg  WEE ;
reg  WEF ;
reg  WEG ;
reg  WEH ;
reg  WEI ;
reg  WEJ ;
reg  WEK ;
reg  WEL ;
reg  WEM ;
reg  WEN ;
reg  WEO ;
reg  WEP ;
reg  WFA ;
reg  WFB ;
reg  WFC ;
reg  WFD ;
reg  WFE ;
reg  WFF ;
reg  WFG ;
reg  WFH ;
reg  WFI ;
reg  WFJ ;
reg  WFK ;
reg  WFL ;
reg  WFM ;
reg  WFN ;
reg  WFO ;
reg  WFP ;
reg  WGA ;
reg  WGB ;
reg  WGC ;
reg  WGD ;
reg  WGE ;
reg  WGF ;
reg  WGG ;
reg  WGH ;
reg  WGI ;
reg  WGJ ;
reg  WGK ;
reg  WGL ;
reg  WGM ;
reg  WGN ;
reg  WGO ;
reg  WGP ;
reg  WHA ;
reg  WHB ;
reg  WHC ;
reg  WHD ;
reg  WHE ;
reg  WHF ;
reg  WHG ;
reg  WHH ;
reg  WHI ;
reg  WHJ ;
reg  WHK ;
reg  WHL ;
reg  WHM ;
reg  WHN ;
reg  WHO ;
reg  WHP ;
wire  aaa ;
wire  aab ;
wire  aac ;
wire  aad ;
wire  aae ;
wire  aaf ;
wire  aag ;
wire  aah ;
wire  aai ;
wire  aaj ;
wire  aak ;
wire  aal ;
wire  aam ;
wire  aan ;
wire  aao ;
wire  aap ;
wire  aaq ;
wire  aar ;
wire  aas ;
wire  aat ;
wire  aau ;
wire  aav ;
wire  aaw ;
wire  aax ;
wire  aba ;
wire  abb ;
wire  abc ;
wire  abd ;
wire  abe ;
wire  abf ;
wire  abg ;
wire  abh ;
wire  abi ;
wire  abj ;
wire  abk ;
wire  abl ;
wire  abm ;
wire  abn ;
wire  abo ;
wire  abp ;
wire  abq ;
wire  abr ;
wire  abs ;
wire  abt ;
wire  abu ;
wire  abv ;
wire  abw ;
wire  abx ;
wire  aca ;
wire  acb ;
wire  acc ;
wire  acd ;
wire  ace ;
wire  acf ;
wire  acg ;
wire  ach ;
wire  aci ;
wire  acj ;
wire  ack ;
wire  acl ;
wire  acm ;
wire  acn ;
wire  aco ;
wire  acp ;
wire  acq ;
wire  acr ;
wire  acs ;
wire  act ;
wire  acu ;
wire  acv ;
wire  acw ;
wire  acx ;
wire  ada ;
wire  adb ;
wire  adc ;
wire  add ;
wire  ade ;
wire  adf ;
wire  adg ;
wire  adh ;
wire  adi ;
wire  adj ;
wire  adk ;
wire  adl ;
wire  adm ;
wire  adn ;
wire  ado ;
wire  adp ;
wire  adq ;
wire  adr ;
wire  ads ;
wire  adt ;
wire  adu ;
wire  adv ;
wire  adw ;
wire  adx ;
wire  aea ;
wire  aeb ;
wire  aec ;
wire  aed ;
wire  aee ;
wire  aef ;
wire  aeg ;
wire  aeh ;
wire  aei ;
wire  aej ;
wire  aek ;
wire  ael ;
wire  aem ;
wire  aen ;
wire  aeo ;
wire  aep ;
wire  aeq ;
wire  aer ;
wire  aes ;
wire  aet ;
wire  aeu ;
wire  aev ;
wire  aew ;
wire  aex ;
wire  afa ;
wire  afb ;
wire  afc ;
wire  afd ;
wire  afe ;
wire  aff ;
wire  afg ;
wire  afh ;
wire  afi ;
wire  afj ;
wire  afk ;
wire  afl ;
wire  afm ;
wire  afn ;
wire  afo ;
wire  afp ;
wire  afq ;
wire  afr ;
wire  afs ;
wire  aft ;
wire  afu ;
wire  afv ;
wire  afw ;
wire  afx ;
wire  aga ;
wire  agb ;
wire  agc ;
wire  agd ;
wire  age ;
wire  agf ;
wire  agg ;
wire  agh ;
wire  agi ;
wire  agj ;
wire  agk ;
wire  agl ;
wire  agm ;
wire  agn ;
wire  ago ;
wire  agp ;
wire  agq ;
wire  agr ;
wire  ags ;
wire  agt ;
wire  agu ;
wire  agv ;
wire  agw ;
wire  agx ;
wire  aha ;
wire  ahb ;
wire  ahc ;
wire  ahd ;
wire  ahe ;
wire  ahf ;
wire  ahg ;
wire  ahh ;
wire  ahi ;
wire  ahj ;
wire  ahk ;
wire  ahl ;
wire  ahm ;
wire  ahn ;
wire  aho ;
wire  ahp ;
wire  ahq ;
wire  ahr ;
wire  ahs ;
wire  aht ;
wire  ahu ;
wire  ahv ;
wire  ahw ;
wire  ahx ;
wire  aia ;
wire  aib ;
wire  aic ;
wire  aid ;
wire  aie ;
wire  aif ;
wire  aig ;
wire  aih ;
wire  aii ;
wire  aij ;
wire  aik ;
wire  ail ;
wire  aim ;
wire  ain ;
wire  aio ;
wire  aip ;
wire  aiq ;
wire  air ;
wire  ais ;
wire  ait ;
wire  aiu ;
wire  aiv ;
wire  aiw ;
wire  aix ;
wire  baa ;
wire  BAA ;
wire  bab ;
wire  BAB ;
wire  bac ;
wire  BAC ;
wire  bad ;
wire  BAD ;
wire  bae ;
wire  BAE ;
wire  baf ;
wire  BAF ;
wire  bag ;
wire  BAG ;
wire  bah ;
wire  BAH ;
wire  bba ;
wire  BBA ;
wire  bbb ;
wire  BBB ;
wire  bbc ;
wire  BBC ;
wire  bbd ;
wire  BBD ;
wire  bbe ;
wire  BBE ;
wire  bbf ;
wire  BBF ;
wire  bbg ;
wire  BBG ;
wire  bbh ;
wire  BBH ;
wire  bca ;
wire  BCA ;
wire  bcb ;
wire  BCB ;
wire  bcc ;
wire  BCC ;
wire  bcd ;
wire  BCD ;
wire  bce ;
wire  BCE ;
wire  bcf ;
wire  BCF ;
wire  bcg ;
wire  BCG ;
wire  bch ;
wire  BCH ;
wire  bda ;
wire  BDA ;
wire  bdb ;
wire  BDB ;
wire  bdc ;
wire  BDC ;
wire  bdd ;
wire  BDD ;
wire  bde ;
wire  BDE ;
wire  bdf ;
wire  BDF ;
wire  bdg ;
wire  BDG ;
wire  bdh ;
wire  BDH ;
wire  caa ;
wire  cab ;
wire  cba ;
wire  cbb ;
wire  cca ;
wire  ccb ;
wire  cda ;
wire  cdb ;
wire  daa ;
wire  dab ;
wire  dac ;
wire  dad ;
wire  dae ;
wire  daf ;
wire  dag ;
wire  dah ;
wire  dai ;
wire  daj ;
wire  dak ;
wire  dal ;
wire  dba ;
wire  dbb ;
wire  dbc ;
wire  dbe ;
wire  dbf ;
wire  dbg ;
wire  dbi ;
wire  dbj ;
wire  dbk ;
wire  eaa ;
wire  eab ;
wire  eac ;
wire  ead ;
wire  EBA ;
wire  EBB ;
wire  EBC ;
wire  faa ;
wire  fab ;
wire  fac ;
wire  fad ;
wire  gaa ;
wire  gab ;
wire  gac ;
wire  haa ;
wire  hab ;
wire  hac ;
wire  hba ;
wire  hbb ;
wire  hbc ;
wire  hca ;
wire  hcb ;
wire  hcc ;
wire  hda ;
wire  hdb ;
wire  hdc ;
wire  hea ;
wire  heb ;
wire  hec ;
wire  hfa ;
wire  hfb ;
wire  hfc ;
wire  hga ;
wire  hgb ;
wire  hgc ;
wire  hha ;
wire  hhb ;
wire  hhc ;
wire  hia ;
wire  hib ;
wire  hic ;
wire  hid ;
wire  iaa ;
wire  iab ;
wire  iac ;
wire  iad ;
wire  iae ;
wire  iaf ;
wire  iag ;
wire  iah ;
wire  iai ;
wire  iaj ;
wire  iak ;
wire  ial ;
wire  iam ;
wire  ian ;
wire  iao ;
wire  iap ;
wire  iba ;
wire  ibb ;
wire  ibc ;
wire  ibd ;
wire  ibe ;
wire  ibf ;
wire  ibg ;
wire  ibh ;
wire  ibi ;
wire  ibj ;
wire  ibk ;
wire  ibl ;
wire  ibm ;
wire  ibn ;
wire  ibo ;
wire  ibp ;
wire  ica ;
wire  icb ;
wire  icc ;
wire  icd ;
wire  ice ;
wire  icf ;
wire  icg ;
wire  ich ;
wire  ici ;
wire  icj ;
wire  ick ;
wire  icl ;
wire  icm ;
wire  icn ;
wire  ico ;
wire  icp ;
wire  ida ;
wire  idb ;
wire  idc ;
wire  idd ;
wire  ide ;
wire  idf ;
wire  idg ;
wire  idh ;
wire  idi ;
wire  idj ;
wire  idk ;
wire  idl ;
wire  idm ;
wire  idn ;
wire  ido ;
wire  idp ;
wire  iea ;
wire  ieb ;
wire  iec ;
wire  ied ;
wire  iee ;
wire  ief ;
wire  ieg ;
wire  ieh ;
wire  iei ;
wire  iej ;
wire  iek ;
wire  iel ;
wire  iem ;
wire  ien ;
wire  ieo ;
wire  iep ;
wire  ieq ;
wire  ier ;
wire  ies ;
wire  iet ;
wire  ieu ;
wire  iev ;
wire  iew ;
wire  iex ;
wire  ifa ;
wire  ifb ;
wire  ifc ;
wire  ifd ;
wire  iga ;
wire  igb ;
wire  igc ;
wire  iha ;
wire  ihb ;
wire  ijb ;
wire  ijd ;
wire  ije ;
wire  ijf ;
wire  jaa ;
wire  JAA ;
wire  jab ;
wire  JAB ;
wire  jac ;
wire  JAC ;
wire  jba ;
wire  JBA ;
wire  jbb ;
wire  JBB ;
wire  jbc ;
wire  JBC ;
wire  jca ;
wire  JCA ;
wire  jcb ;
wire  JCB ;
wire  jcc ;
wire  JCC ;
wire  jda ;
wire  JDA ;
wire  jdb ;
wire  JDB ;
wire  jdc ;
wire  JDC ;
wire  jea ;
wire  JEA ;
wire  jeb ;
wire  JEB ;
wire  jec ;
wire  JEC ;
wire  jed ;
wire  JED ;
wire  jee ;
wire  JEE ;
wire  jfa ;
wire  JFA ;
wire  jfb ;
wire  JFB ;
wire  jga ;
wire  JGA ;
wire  jgb ;
wire  JGB ;
wire  jgc ;
wire  JGC ;
wire  jha ;
wire  JHA ;
wire  jhb ;
wire  JHB ;
wire  jia ;
wire  JIA ;
wire  jib ;
wire  JIB ;
wire  jic ;
wire  JIC ;
wire  jid ;
wire  JID ;
wire  jja ;
wire  JJA ;
wire  jjb ;
wire  JJB ;
wire  jjc ;
wire  JJC ;
wire  jjd ;
wire  JJD ;
wire  jka ;
wire  JKA ;
wire  jkb ;
wire  JKB ;
wire  jkc ;
wire  JKC ;
wire  jkd ;
wire  JKD ;
wire  jla ;
wire  JLA ;
wire  jlb ;
wire  JLB ;
wire  jlc ;
wire  JLC ;
wire  jld ;
wire  JLD ;
wire  jle ;
wire  JLE ;
wire  jma ;
wire  JMA ;
wire  jmb ;
wire  JMB ;
wire  jmc ;
wire  JMC ;
wire  jna ;
wire  JNA ;
wire  jnb ;
wire  JNB ;
wire  jnc ;
wire  JNC ;
wire  jnd ;
wire  JND ;
wire  joa ;
wire  JOA ;
wire  jpa ;
wire  JPA ;
wire  jpb ;
wire  JPB ;
wire  jpc ;
wire  JPC ;
wire  jpe ;
wire  JPE ;
wire  jpf ;
wire  JPF ;
wire  jqa ;
wire  JQA ;
wire  jqb ;
wire  JQB ;
wire  jra ;
wire  JRA ;
wire  kaa ;
wire  KAA ;
wire  kab ;
wire  KAB ;
wire  kac ;
wire  KAC ;
wire  kad ;
wire  KAD ;
wire  kae ;
wire  KAE ;
wire  kaf ;
wire  KAF ;
wire  kag ;
wire  KAG ;
wire  kah ;
wire  KAH ;
wire  kai ;
wire  KAI ;
wire  kaj ;
wire  KAJ ;
wire  kak ;
wire  KAK ;
wire  kal ;
wire  KAL ;
wire  kam ;
wire  KAM ;
wire  kan ;
wire  KAN ;
wire  kao ;
wire  KAO ;
wire  kap ;
wire  KAP ;
wire  kba ;
wire  KBA ;
wire  kbb ;
wire  KBB ;
wire  kbc ;
wire  KBC ;
wire  kbd ;
wire  KBD ;
wire  kbe ;
wire  KBE ;
wire  kbf ;
wire  KBF ;
wire  kbg ;
wire  KBG ;
wire  kbh ;
wire  KBH ;
wire  kbi ;
wire  KBI ;
wire  kbj ;
wire  KBJ ;
wire  kbk ;
wire  KBK ;
wire  kbl ;
wire  KBL ;
wire  kbm ;
wire  KBM ;
wire  kbn ;
wire  KBN ;
wire  kbo ;
wire  KBO ;
wire  kbp ;
wire  KBP ;
wire  kca ;
wire  KCA ;
wire  kcb ;
wire  KCB ;
wire  kcc ;
wire  KCC ;
wire  kcd ;
wire  KCD ;
wire  kce ;
wire  KCE ;
wire  kcf ;
wire  KCF ;
wire  kcg ;
wire  KCG ;
wire  kch ;
wire  KCH ;
wire  kci ;
wire  KCI ;
wire  kcj ;
wire  KCJ ;
wire  kck ;
wire  KCK ;
wire  kcl ;
wire  KCL ;
wire  kcm ;
wire  KCM ;
wire  kcn ;
wire  KCN ;
wire  kco ;
wire  KCO ;
wire  kcp ;
wire  KCP ;
wire  kda ;
wire  KDA ;
wire  kdb ;
wire  KDB ;
wire  kdc ;
wire  KDC ;
wire  kdd ;
wire  KDD ;
wire  kde ;
wire  kdf ;
wire  KDF ;
wire  kdg ;
wire  KDG ;
wire  kdh ;
wire  KDH ;
wire  kdi ;
wire  KDI ;
wire  kdj ;
wire  KDJ ;
wire  kdk ;
wire  KDK ;
wire  kdl ;
wire  KDL ;
wire  kdm ;
wire  KDM ;
wire  kdn ;
wire  KDN ;
wire  kdo ;
wire  KDO ;
wire  kdp ;
wire  KDP ;
wire  oaa ;
wire  oab ;
wire  oac ;
wire  oad ;
wire  oae ;
wire  oaf ;
wire  oag ;
wire  oah ;
wire  oai ;
wire  oaj ;
wire  oak ;
wire  oal ;
wire  oam ;
wire  oan ;
wire  oao ;
wire  oap ;
wire  oba ;
wire  obb ;
wire  obc ;
wire  obd ;
wire  obe ;
wire  obf ;
wire  obg ;
wire  obh ;
wire  obi ;
wire  obj ;
wire  obk ;
wire  obl ;
wire  obm ;
wire  obn ;
wire  obo ;
wire  obp ;
wire  oca ;
wire  ocb ;
wire  occ ;
wire  ocd ;
wire  oce ;
wire  ocf ;
wire  ocg ;
wire  och ;
wire  oci ;
wire  ocj ;
wire  ock ;
wire  ocl ;
wire  ocm ;
wire  ocn ;
wire  oco ;
wire  ocp ;
wire  oda ;
wire  odb ;
wire  odc ;
wire  odd ;
wire  ode ;
wire  odf ;
wire  odg ;
wire  odh ;
wire  odi ;
wire  odj ;
wire  odk ;
wire  odl ;
wire  odm ;
wire  odn ;
wire  odo ;
wire  odp ;
wire  OEA ;
wire  OEB ;
wire  OEC ;
wire  OED ;
wire  OEE ;
wire  OEF ;
wire  OEG ;
wire  OEH ;
wire  OEI ;
wire  OEJ ;
wire  OEK ;
wire  OEL ;
wire  OEM ;
wire  OEN ;
wire  OEO ;
wire  OEP ;
wire  OFA ;
wire  OFB ;
wire  OFC ;
wire  OFD ;
wire  OFE ;
wire  OFF ;
wire  OFG ;
wire  OFH ;
wire  OFI ;
wire  OFJ ;
wire  OFK ;
wire  OFL ;
wire  OFM ;
wire  OFN ;
wire  OFO ;
wire  OFP ;
wire  OGA ;
wire  OGB ;
wire  OGC ;
wire  OGD ;
wire  OGE ;
wire  OGF ;
wire  OGG ;
wire  OGH ;
wire  OGI ;
wire  OGJ ;
wire  OGK ;
wire  OGL ;
wire  OGM ;
wire  OGN ;
wire  OGO ;
wire  OGP ;
wire  OHA ;
wire  OHB ;
wire  OHC ;
wire  OHD ;
wire  OHE ;
wire  OHF ;
wire  OHG ;
wire  OHH ;
wire  OHI ;
wire  OHJ ;
wire  OHK ;
wire  OHL ;
wire  OHM ;
wire  OHN ;
wire  OHO ;
wire  OHP ;
wire  oja ;
wire  ojb ;
wire  ojc ;
wire  OJD ;
wire  OJE ;
wire  oka ;
wire  okb ;
wire  okc ;
wire  okd ;
wire  oke ;
wire  OKF ;
wire  okg ;
wire  okh ;
wire  OKI ;
wire  OKJ ;
wire  OKK ;
wire  OKL ;
wire  OKM ;
wire  OKN ;
wire  OKO ;
wire  OKP ;
wire  OKQ ;
wire  OKR ;
wire  OKS ;
wire  OKT ;
wire  OKU ;
wire  OKV ;
wire  OKW ;
wire  OKX ;
wire  paa ;
wire  pab ;
wire  pac ;
wire  pad ;
wire  pae ;
wire  paf ;
wire  pba ;
wire  pbb ;
wire  pbc ;
wire  pbd ;
wire  pbe ;
wire  pbf ;
wire  pca ;
wire  pcb ;
wire  pcc ;
wire  pcd ;
wire  pce ;
wire  pcf ;
wire  pda ;
wire  pdb ;
wire  pdc ;
wire  pdd ;
wire  pde ;
wire  pdf ;
wire  pea ;
wire  peb ;
wire  pec ;
wire  pfa ;
wire  pfb ;
wire  pfc ;
wire  pga ;
wire  pgb ;
wire  pgc ;
wire  QAA ;
wire  QAB ;
wire  QAC ;
wire  QAD ;
wire  qae ;
wire  qba ;
wire  qbb ;
wire  qbc ;
wire  qbd ;
wire  qbe ;
wire  qca ;
wire  qcb ;
wire  qcc ;
wire  qcd ;
wire  qce ;
wire  qda ;
wire  QDB ;
wire  qdc ;
wire  qdd ;
wire  qde ;
wire  qdi ;
wire  qdj ;
wire  qdk ;
wire  qdl ;
wire  qeb ;
wire  QEC ;
wire  QED ;
wire  qfa ;
wire  QHA ;
wire  QHB ;
wire  QHC ;
wire  QHD ;
wire  qja ;
wire  qjb ;
wire  qjc ;
wire  qjd ;
wire  qje ;
wire  qjf ;
wire  qjg ;
wire  qjh ;
wire  qji ;
wire  qjj ;
wire  qjk ;
wire  qjm ;
wire  qjn ;
wire  qjp ;
wire  qka ;
wire  qkb ;
wire  QLA ;
wire  QLB ;
wire  QLC ;
wire  qld ;
wire  QLE ;
wire  qlf ;
wire  qlg ;
wire  qlh ;
wire  qpa ;
wire  qpb ;
wire  qpc ;
wire  qpd ;
wire  qpe ;
wire  qqa ;
wire  qqb ;
wire  qqc ;
wire  qqd ;
wire  taa ;
wire  tab ;
wire  tac ;
wire  tad ;
wire  tae ;
wire  taf ;
wire  tag ;
wire  tah ;
wire  tba ;
wire  tbb ;
wire  tbc ;
wire  tbd ;
wire  tbe ;
wire  tbf ;
wire  tbg ;
wire  tbh ;
wire  tca ;
wire  tcb ;
wire  tcc ;
wire  tcd ;
wire  tce ;
wire  tcf ;
wire  tcg ;
wire  tch ;
wire  tda ;
wire  tdb ;
wire  tdc ;
wire  tdd ;
wire  tde ;
wire  tdf ;
wire  tdg ;
wire  tdh ;
wire  tea ;
wire  teb ;
wire  tec ;
wire  ted ;
wire  tee ;
wire  tef ;
wire  teg ;
wire  teh ;
wire  tfa ;
wire  tfb ;
wire  tfc ;
wire  tfd ;
wire  TGA ;
wire  TGB ;
wire  TGC ;
wire  TGD ;
wire  tja ;
wire  tjb ;
wire  tjc ;
wire  tjd ;
wire  tma ;
wire  uaa ;
wire  uab ;
wire  uac ;
wire  uad ;
wire  uae ;
wire  uaf ;
wire  uag ;
wire  uai ;
wire  uaj ;
wire  uak ;
wire  ual ;
wire  uam ;
wire  uan ;
wire  uao ;
wire  uba ;
wire  ubb ;
wire  ubc ;
wire  ubd ;
wire  ube ;
wire  ubf ;
wire  ubg ;
wire  ubi ;
wire  ubj ;
wire  ubk ;
wire  ubl ;
wire  ubm ;
wire  ubn ;
wire  ubo ;
wire  uca ;
wire  ucb ;
wire  ucc ;
wire  ucd ;
wire  uce ;
wire  ucf ;
wire  ucg ;
wire  uci ;
wire  ucj ;
wire  uck ;
wire  ucl ;
wire  ucm ;
wire  ucn ;
wire  uco ;
wire  uda ;
wire  udb ;
wire  udc ;
wire  udd ;
wire  ude ;
wire  udf ;
wire  udg ;
wire  udi ;
wire  udj ;
wire  udk ;
wire  udl ;
wire  udm ;
wire  udn ;
wire  udo ;
wire  uea ;
wire  ueb ;
wire  uec ;
wire  ued ;
wire  uee ;
wire  uef ;
wire  ueg ;
wire  uei ;
wire  uej ;
wire  uek ;
wire  uel ;
wire  uem ;
wire  uen ;
wire  ueo ;
wire  ufa ;
wire  ufb ;
wire  ufc ;
wire  ufd ;
wire  ufe ;
wire  uff ;
wire  ufg ;
wire  ufi ;
wire  ufj ;
wire  ufk ;
wire  ufl ;
wire  ufm ;
wire  ufn ;
wire  ufo ;
wire  uga ;
wire  ugb ;
wire  ugc ;
wire  ugd ;
wire  uge ;
wire  ugf ;
wire  ugg ;
wire  ugi ;
wire  ugj ;
wire  ugk ;
wire  ugl ;
wire  ugm ;
wire  ugn ;
wire  ugo ;
wire  uha ;
wire  uhb ;
wire  uhc ;
wire  uhd ;
wire  uhe ;
wire  uhf ;
wire  uhg ;
wire  uhi ;
wire  uhj ;
wire  uhk ;
wire  uhl ;
wire  uhm ;
wire  uhn ;
wire  uho ;
wire  uia ;
wire  uib ;
wire  uic ;
wire  uid ;
wire  uie ;
wire  uif ;
wire  uig ;
wire  uii ;
wire  uij ;
wire  uik ;
wire  uil ;
wire  uim ;
wire  uin ;
wire  uio ;
wire  uja ;
wire  ujb ;
wire  ujc ;
wire  ujd ;
wire  uje ;
wire  ujf ;
wire  ujg ;
wire  uji ;
wire  ujj ;
wire  ujk ;
wire  ujl ;
wire  ujm ;
wire  ujn ;
wire  ujo ;
wire  uka ;
wire  ukb ;
wire  ukc ;
wire  ukd ;
wire  uke ;
wire  ukf ;
wire  ukg ;
wire  uki ;
wire  ukj ;
wire  ukk ;
wire  ukl ;
wire  ukm ;
wire  ukn ;
wire  uko ;
wire  ula ;
wire  ulb ;
wire  ulc ;
wire  uld ;
wire  ule ;
wire  ulf ;
wire  ulg ;
wire  uli ;
wire  ulj ;
wire  ulk ;
wire  ull ;
wire  ulm ;
wire  uln ;
wire  ulo ;
wire  uma ;
wire  umb ;
wire  umc ;
wire  umd ;
wire  ume ;
wire  umf ;
wire  umg ;
wire  umi ;
wire  umj ;
wire  umk ;
wire  uml ;
wire  umm ;
wire  umn ;
wire  umo ;
wire  una ;
wire  unb ;
wire  unc ;
wire  und ;
wire  une ;
wire  unf ;
wire  ung ;
wire  uni ;
wire  unj ;
wire  unk ;
wire  unl ;
wire  unm ;
wire  unn ;
wire  uno ;
wire  uoa ;
wire  uob ;
wire  uoc ;
wire  uod ;
wire  uoe ;
wire  uof ;
wire  uog ;
wire  uoi ;
wire  uoj ;
wire  uok ;
wire  uol ;
wire  uom ;
wire  uon ;
wire  uoo ;
wire  upa ;
wire  upb ;
wire  upc ;
wire  upd ;
wire  upe ;
wire  upf ;
wire  upg ;
wire  upi ;
wire  upj ;
wire  upk ;
wire  upl ;
wire  upm ;
wire  upn ;
wire  upo ;
wire  vaa ;
wire  vab ;
wire  vac ;
wire  vad ;
wire  vae ;
wire  vaf ;
wire  vag ;
wire  vah ;
wire  vai ;
wire  vaj ;
wire  vak ;
wire  val ;
wire  vam ;
wire  van ;
wire  vao ;
wire  vap ;
wire  vba ;
wire  vbb ;
wire  vbc ;
wire  vbd ;
wire  vbe ;
wire  vbf ;
wire  vbg ;
wire  vbh ;
wire  vbi ;
wire  vbj ;
wire  vbk ;
wire  vbl ;
wire  vbm ;
wire  vbn ;
wire  vbo ;
wire  vbp ;
wire  vca ;
wire  vcb ;
wire  vcc ;
wire  vcd ;
wire  vce ;
wire  vcf ;
wire  vcg ;
wire  vch ;
wire  vci ;
wire  vcj ;
wire  vck ;
wire  vcl ;
wire  vcm ;
wire  vcn ;
wire  vco ;
wire  vcp ;
wire  vda ;
wire  vdb ;
wire  vdc ;
wire  vdd ;
wire  vde ;
wire  vdf ;
wire  vdg ;
wire  vdh ;
wire  vdi ;
wire  vdj ;
wire  vdk ;
wire  vdl ;
wire  vdm ;
wire  vdn ;
wire  vdo ;
wire  vdp ;
wire  waa ;
wire  wab ;
wire  wac ;
wire  wad ;
wire  wae ;
wire  waf ;
wire  wag ;
wire  wah ;
wire  wai ;
wire  waj ;
wire  wak ;
wire  wal ;
wire  wam ;
wire  wan ;
wire  wao ;
wire  wap ;
wire  wba ;
wire  wbb ;
wire  wbc ;
wire  wbd ;
wire  wbe ;
wire  wbf ;
wire  wbg ;
wire  wbh ;
wire  wbi ;
wire  wbj ;
wire  wbk ;
wire  wbl ;
wire  wbm ;
wire  wbn ;
wire  wbo ;
wire  wbp ;
wire  wca ;
wire  wcb ;
wire  wcc ;
wire  wcd ;
wire  wce ;
wire  wcf ;
wire  wcg ;
wire  wch ;
wire  wci ;
wire  wcj ;
wire  wck ;
wire  wcl ;
wire  wcm ;
wire  wcn ;
wire  wco ;
wire  wcp ;
wire  wda ;
wire  wdb ;
wire  wdc ;
wire  wdd ;
wire  wde ;
wire  wdf ;
wire  wdg ;
wire  wdh ;
wire  wdi ;
wire  wdj ;
wire  wdk ;
wire  wdl ;
wire  wdm ;
wire  wdn ;
wire  wdo ;
wire  wdp ;
wire  wea ;
wire  web ;
wire  wec ;
wire  wed ;
wire  wee ;
wire  wef ;
wire  weg ;
wire  weh ;
wire  wei ;
wire  wej ;
wire  wek ;
wire  wel ;
wire  wem ;
wire  wen ;
wire  weo ;
wire  wep ;
wire  wfa ;
wire  wfb ;
wire  wfc ;
wire  wfd ;
wire  wfe ;
wire  wff ;
wire  wfg ;
wire  wfh ;
wire  wfi ;
wire  wfj ;
wire  wfk ;
wire  wfl ;
wire  wfm ;
wire  wfn ;
wire  wfo ;
wire  wfp ;
wire  wga ;
wire  wgb ;
wire  wgc ;
wire  wgd ;
wire  wge ;
wire  wgf ;
wire  wgg ;
wire  wgh ;
wire  wgi ;
wire  wgj ;
wire  wgk ;
wire  wgl ;
wire  wgm ;
wire  wgn ;
wire  wgo ;
wire  wgp ;
wire  wha ;
wire  whb ;
wire  whc ;
wire  whd ;
wire  whe ;
wire  whf ;
wire  whg ;
wire  whh ;
wire  whi ;
wire  whj ;
wire  whk ;
wire  whl ;
wire  whm ;
wire  whn ;
wire  who ;
wire  whp ;
wire  ZZI ;
wire  ZZO ;
assign ZZI = 1'b1;
assign ZZO = 1'b0;
assign uaa = ~UAA;  //complement 
assign uba = ~UBA;  //complement 
assign uaf = ~UAF;  //complement 
assign uag = ~UAG;  //complement 
assign ubf = ~UBF;  //complement 
assign ubg = ~UBG;  //complement 
assign uab = ~UAB;  //complement 
assign ubb = ~UBB;  //complement 
assign uae = ~UAE;  //complement 
assign ube = ~UBE;  //complement 
assign uac = ~UAC;  //complement 
assign ubc = ~UBC;  //complement 
assign uad = ~UAD;  //complement 
assign ubd = ~UBD;  //complement 
assign uce = ~UCE;  //complement 
assign ude = ~UDE;  //complement 
assign uca = ~UCA;  //complement 
assign uda = ~UDA;  //complement 
assign ucf = ~UCF;  //complement 
assign ucg = ~UCG;  //complement 
assign ucb = ~UCB;  //complement 
assign udb = ~UDB;  //complement 
assign ucc = ~UCC;  //complement 
assign udc = ~UDC;  //complement 
assign udf = ~UDF;  //complement 
assign udg = ~UDG;  //complement 
assign ucd = ~UCD;  //complement 
assign udd = ~UDD;  //complement 
assign qda = ~QDA;  //complement 
assign tea = ~TEA;  //complement 
assign oaa = ~OAA;  //complement 
assign vaa = ~VAA;  //complement 
assign KAA =  WEA & TFA  |  VAA & TGA  ; 
assign kaa = ~KAA;  //complement 
assign KAI =  WEI & TFA  |  VAI & TGA  ; 
assign kai = ~KAI;  //complement 
assign oai = ~OAI;  //complement 
assign vai = ~VAI;  //complement 
assign waa = ~WAA;  //complement 
assign wai = ~WAI;  //complement 
assign wea = ~WEA;  //complement 
assign wei = ~WEI;  //complement 
assign oba = ~OBA;  //complement 
assign vba = ~VBA;  //complement 
assign KDA =  WHA & TFD  |  VDA & TGD  ; 
assign kda = ~KDA;  //complement 
assign KBA =  WFA & TFB  |  VBA & TGB  ; 
assign kba = ~KBA;  //complement 
assign KBI =  WFI & TFB  |  VBI & TGB  ; 
assign kbi = ~KBI;  //complement 
assign obi = ~OBI;  //complement 
assign vbi = ~VBI;  //complement 
assign wba = ~WBA;  //complement 
assign wbi = ~WBI;  //complement 
assign wfa = ~WFA;  //complement 
assign wfi = ~WFI;  //complement 
assign oca = ~OCA;  //complement 
assign vca = ~VCA;  //complement 
assign jac =  qba & qca  ; 
assign JAC = ~jac;  //complement 
assign KCA =  WGA & TFC  |  VCA & TGC  ; 
assign kca = ~KCA;  //complement 
assign KCI =  WGI & TFC  |  VCI & TGC  ; 
assign kci = ~KCI;  //complement 
assign qqa = ~QQA;  //complement 
assign oci = ~OCI;  //complement 
assign vci = ~VCI;  //complement 
assign wca = ~WCA;  //complement 
assign wci = ~WCI;  //complement 
assign wga = ~WGA;  //complement 
assign wgi = ~WGI;  //complement 
assign QHA = ~qha;  //complement 
assign oda = ~ODA;  //complement 
assign vda = ~VDA;  //complement 
assign KDI =  WHI & TFD  |  VDI & TGD  ; 
assign kdi = ~KDI;  //complement 
assign JIA =  daj & dai & QJM  ; 
assign jia = ~JIA;  //complement  
assign JNA =  daf & dae  ; 
assign jna = ~JNA;  //complement 
assign odi = ~ODI;  //complement 
assign vdi = ~VDI;  //complement 
assign wda = ~WDA;  //complement 
assign wdi = ~WDI;  //complement 
assign wha = ~WHA;  //complement 
assign whi = ~WHI;  //complement 
assign taa = ~TAA;  //complement 
assign tba = ~TBA;  //complement 
assign tca = ~TCA;  //complement 
assign tda = ~TDA;  //complement 
assign aga = ~AGA;  //complement 
assign agi = ~AGI;  //complement 
assign agq = ~AGQ;  //complement 
assign aea = ~AEA;  //complement 
assign aei = ~AEI;  //complement 
assign aeq = ~AEQ;  //complement 
assign aca = ~ACA;  //complement 
assign aci = ~ACI;  //complement 
assign OKJ = ~okj;  //complement 
assign acq = ~ACQ;  //complement 
assign aaa = ~AAA;  //complement 
assign aai = ~AAI;  //complement 
assign aaq = ~AAQ;  //complement 
assign aha = ~AHA;  //complement 
assign ahi = ~AHI;  //complement 
assign ahq = ~AHQ;  //complement 
assign afa = ~AFA;  //complement 
assign afi = ~AFI;  //complement 
assign afq = ~AFQ;  //complement 
assign aia = ~AIA;  //complement 
assign ada = ~ADA;  //complement 
assign adi = ~ADI;  //complement 
assign adq = ~ADQ;  //complement 
assign aii = ~AII;  //complement 
assign aba = ~ABA;  //complement 
assign abi = ~ABI;  //complement 
assign abq = ~ABQ;  //complement 
assign aiq = ~AIQ;  //complement 
assign BDA =  AIA & aha  |  aia & AHA  |  AII & ahi  |  aii & AHI  |  AIQ & ahq  |  aiq & AHQ  ;
assign bda = ~BDA;  //complement 
assign BCA =  AIA & afa  |  aia & AFA  |  AII & afi  |  aii & AFI  |  AIQ & afq  |  aiq & AFQ  ;
assign bca = ~BCA;  //complement 
assign BBA =  AIA & ada  |  aia & ADA  |  AII & adi  |  aii & ADI  |  AIQ & adq  |  aiq & ADQ  ;
assign bba = ~BBA;  //complement 
assign BAA =  AIA & aba  |  aia & ABA  |  AII & abi  |  aii & ABI  |  AIQ & abq  |  aiq & ABQ  ;
assign baa = ~BAA;  //complement 
assign qjk = ~QJK;  //complement 
assign OEA = ~oea;  //complement 
assign OEI = ~oei;  //complement 
assign OFA = ~ofa;  //complement 
assign OFI = ~ofi;  //complement 
assign JPA =  QQA & QQB & QQC & QQD & QJK  ; 
assign jpa = ~JPA;  //complement  
assign okb = ~OKB;  //complement 
assign qjh = ~QJH;  //complement 
assign OGA = ~oga;  //complement 
assign OGI = ~ogi;  //complement 
assign OHA = ~oha;  //complement 
assign OHI = ~ohi;  //complement 
assign qce = ~QCE;  //complement 
assign qde = ~QDE;  //complement 
assign qae = ~QAE;  //complement 
assign qbe = ~QBE;  //complement 
assign qba = ~QBA;  //complement 
assign qca = ~QCA;  //complement 
assign qdi = ~QDI;  //complement 
assign qpa = ~QPA;  //complement 
assign QAA = ~qaa;  //complement 
assign QAB = ~qab;  //complement 
assign QAC = ~qac;  //complement 
assign QAD = ~qad;  //complement 
assign paa = ~PAA;  //complement 
assign pac = ~PAC;  //complement 
assign pae = ~PAE;  //complement 
assign pab = ~PAB;  //complement 
assign pad = ~PAD;  //complement 
assign paf = ~PAF;  //complement 
assign JAA =  QPA  ; 
assign jaa = ~JAA;  //complement 
assign JAB =  QPA & PAA  ; 
assign jab = ~JAB;  //complement 
assign uea = ~UEA;  //complement 
assign ufa = ~UFA;  //complement 
assign uef = ~UEF;  //complement 
assign ueg = ~UEG;  //complement 
assign ueb = ~UEB;  //complement 
assign ufb = ~UFB;  //complement 
assign uee = ~UEE;  //complement 
assign ufe = ~UFE;  //complement 
assign uec = ~UEC;  //complement 
assign ufc = ~UFC;  //complement 
assign uff = ~UFF;  //complement 
assign ufg = ~UFG;  //complement 
assign ued = ~UED;  //complement 
assign ufd = ~UFD;  //complement 
assign uga = ~UGA;  //complement 
assign uha = ~UHA;  //complement 
assign ugf = ~UGF;  //complement 
assign ugg = ~UGG;  //complement 
assign ugb = ~UGB;  //complement 
assign uhb = ~UHB;  //complement 
assign uge = ~UGE;  //complement 
assign uhe = ~UHE;  //complement 
assign ugc = ~UGC;  //complement 
assign uhc = ~UHC;  //complement 
assign uhf = ~UHF;  //complement 
assign uhg = ~UHG;  //complement 
assign ugd = ~UGD;  //complement 
assign uhd = ~UHD;  //complement 
assign QDB = ~qdb;  //complement 
assign teb = ~TEB;  //complement 
assign oab = ~OAB;  //complement 
assign vab = ~VAB;  //complement 
assign aec = ~AEC;  //complement 
assign KAB =  WEB & TFA  |  VAB & TGA  ; 
assign kab = ~KAB;  //complement 
assign KAJ =  WEJ & TFA  |  VAJ & TGA  ; 
assign kaj = ~KAJ;  //complement 
assign oaj = ~OAJ;  //complement 
assign vaj = ~VAJ;  //complement 
assign afc = ~AFC;  //complement 
assign wab = ~WAB;  //complement 
assign waj = ~WAJ;  //complement 
assign web = ~WEB;  //complement 
assign wej = ~WEJ;  //complement 
assign obb = ~OBB;  //complement 
assign vbb = ~VBB;  //complement 
assign KDB =  WHB & TFD  |  VDB & TGD  ; 
assign kdb = ~KDB;  //complement 
assign KBB =  WFB & TFB  |  VBB & TGB  ; 
assign kbb = ~KBB;  //complement 
assign KBJ =  WFJ & TFB  |  VBJ & TGB  ; 
assign kbj = ~KBJ;  //complement 
assign wcj = ~WCJ;  //complement 
assign obj = ~OBJ;  //complement 
assign vbj = ~VBJ;  //complement 
assign wbb = ~WBB;  //complement 
assign wbj = ~WBJ;  //complement 
assign wfb = ~WFB;  //complement 
assign wfj = ~WFJ;  //complement 
assign OEC = ~oec;  //complement 
assign ocb = ~OCB;  //complement 
assign vcb = ~VCB;  //complement 
assign jbc =  qbb & qcb  ; 
assign JBC = ~jbc;  //complement 
assign KCB =  WGB & TFC  |  VCB & TGC  ; 
assign kcb = ~KCB;  //complement 
assign KCJ =  WGJ & TFC  |  VCJ & TGC  ; 
assign kcj = ~KCJ;  //complement 
assign qqb = ~QQB;  //complement 
assign ocj = ~OCJ;  //complement 
assign vcj = ~VCJ;  //complement 
assign wcb = ~WCB;  //complement 
assign wgb = ~WGB;  //complement 
assign wgj = ~WGJ;  //complement 
assign QHB = ~qhb;  //complement 
assign odb = ~ODB;  //complement 
assign vdb = ~VDB;  //complement 
assign KDJ =  WHJ & TFD  |  VDJ & TGD  ; 
assign kdj = ~KDJ;  //complement 
assign JIB =  daj & DAI & QJM  ; 
assign jib = ~JIB;  //complement  
assign JNB =  daf & DAE  ; 
assign jnb = ~JNB;  //complement 
assign odj = ~ODJ;  //complement 
assign vdj = ~VDJ;  //complement 
assign wdb = ~WDB;  //complement 
assign wdj = ~WDJ;  //complement 
assign whb = ~WHB;  //complement 
assign whj = ~WHJ;  //complement 
assign tab = ~TAB;  //complement 
assign tbb = ~TBB;  //complement 
assign tcb = ~TCB;  //complement 
assign tdb = ~TDB;  //complement 
assign agb = ~AGB;  //complement 
assign agj = ~AGJ;  //complement 
assign agr = ~AGR;  //complement 
assign aeb = ~AEB;  //complement 
assign aej = ~AEJ;  //complement 
assign aer = ~AER;  //complement 
assign acb = ~ACB;  //complement 
assign acj = ~ACJ;  //complement 
assign acr = ~ACR;  //complement 
assign aab = ~AAB;  //complement 
assign aaj = ~AAJ;  //complement 
assign aar = ~AAR;  //complement 
assign ahb = ~AHB;  //complement 
assign ahj = ~AHJ;  //complement 
assign ahr = ~AHR;  //complement 
assign afb = ~AFB;  //complement 
assign afj = ~AFJ;  //complement 
assign afr = ~AFR;  //complement 
assign aib = ~AIB;  //complement 
assign adb = ~ADB;  //complement 
assign adj = ~ADJ;  //complement 
assign adr = ~ADR;  //complement 
assign aij = ~AIJ;  //complement 
assign abb = ~ABB;  //complement 
assign abj = ~ABJ;  //complement 
assign abr = ~ABR;  //complement 
assign air = ~AIR;  //complement 
assign BDB =  AIB & ahb  |  aib & AHB  |  AIJ & ahj  |  aij & AHJ  |  AIR & ahr  |  air & AHR  ;
assign bdb = ~BDB;  //complement 
assign BCB =  AIB & afb  |  aib & AFB  |  AIJ & afj  |  aij & AFJ  |  AIR & afr  |  air & AFR  ;
assign bcb = ~BCB;  //complement 
assign BBB =  AIB & adb  |  aib & ADB  |  AIJ & adj  |  aij & ADJ  |  AIR & adr  |  air & ADR  ;
assign bbb = ~BBB;  //complement 
assign BAB =  AIB & abb  |  aib & ABB  |  AIJ & abj  |  aij & ABJ  |  AIR & abr  |  air & ABR  ;
assign bab = ~BAB;  //complement 
assign OEB = ~oeb;  //complement 
assign OEJ = ~oej;  //complement 
assign OFB = ~ofb;  //complement 
assign OFJ = ~ofj;  //complement 
assign OKK = ~okk;  //complement 
assign okc = ~OKC;  //complement 
assign qji = ~QJI;  //complement 
assign OGB = ~ogb;  //complement 
assign OGJ = ~ogj;  //complement 
assign OHB = ~ohb;  //complement 
assign OHJ = ~ohj;  //complement 
assign OKL = ~okl;  //complement 
assign qbb = ~QBB;  //complement 
assign qcb = ~QCB;  //complement 
assign qdj = ~QDJ;  //complement 
assign qpb = ~QPB;  //complement 
assign OKM = ~okm;  //complement 
assign OKN = ~okn;  //complement 
assign pba = ~PBA;  //complement 
assign pbc = ~PBC;  //complement 
assign pbe = ~PBE;  //complement 
assign pbb = ~PBB;  //complement 
assign pbd = ~PBD;  //complement 
assign pbf = ~PBF;  //complement 
assign JBA =  QPB  ; 
assign jba = ~JBA;  //complement 
assign JBB =  QPB & PBA  ; 
assign jbb = ~JBB;  //complement 
assign uia = ~UIA;  //complement 
assign uja = ~UJA;  //complement 
assign uif = ~UIF;  //complement 
assign uig = ~UIG;  //complement 
assign uib = ~UIB;  //complement 
assign ujb = ~UJB;  //complement 
assign uie = ~UIE;  //complement 
assign uje = ~UJE;  //complement 
assign ujc = ~UJC;  //complement 
assign uic = ~UIC;  //complement 
assign ujf = ~UJF;  //complement 
assign ujg = ~UJG;  //complement 
assign uid = ~UID;  //complement 
assign ujd = ~UJD;  //complement 
assign uka = ~UKA;  //complement 
assign ula = ~ULA;  //complement 
assign ukf = ~UKF;  //complement 
assign ukg = ~UKG;  //complement 
assign ukb = ~UKB;  //complement 
assign ulb = ~ULB;  //complement 
assign uke = ~UKE;  //complement 
assign ule = ~ULE;  //complement 
assign ukc = ~UKC;  //complement 
assign ulc = ~ULC;  //complement 
assign ulf = ~ULF;  //complement 
assign ulg = ~ULG;  //complement 
assign ukd = ~UKD;  //complement 
assign uld = ~ULD;  //complement 
assign qdc = ~QDC;  //complement 
assign tec = ~TEC;  //complement 
assign oac = ~OAC;  //complement 
assign vac = ~VAC;  //complement 
assign KAC =  WEC & TFA  |  VAC & TGA  ; 
assign kac = ~KAC;  //complement 
assign KAK =  WEK & TFA  |  VAK & TGA  ; 
assign kak = ~KAK;  //complement 
assign oak = ~OAK;  //complement 
assign vak = ~VAK;  //complement 
assign wac = ~WAC;  //complement 
assign wak = ~WAK;  //complement 
assign wec = ~WEC;  //complement 
assign wek = ~WEK;  //complement 
assign obc = ~OBC;  //complement 
assign vbc = ~VBC;  //complement 
assign KDC =  WHC & TFD  |  VDC & TGD  ; 
assign kdc = ~KDC;  //complement 
assign KBC =  WFC & TFB  |  VBC & TGB  ; 
assign kbc = ~KBC;  //complement 
assign KBK =  WFK & TFB  |  VBK & TGB  ; 
assign kbk = ~KBK;  //complement 
assign obk = ~OBK;  //complement 
assign vbk = ~VBK;  //complement 
assign wbc = ~WBC;  //complement 
assign wbk = ~WBK;  //complement 
assign wfc = ~WFC;  //complement 
assign wfk = ~WFK;  //complement 
assign occ = ~OCC;  //complement 
assign vcc = ~VCC;  //complement 
assign jcc =  qbc & qcc  ; 
assign JCC = ~jcc;  //complement 
assign KCC =  WGC & TFC  |  VCC & TGC  ; 
assign kcc = ~KCC;  //complement 
assign KCK =  WGK & TFC  |  VCK & TGC  ; 
assign kck = ~KCK;  //complement 
assign qqc = ~QQC;  //complement 
assign ock = ~OCK;  //complement 
assign vck = ~VCK;  //complement 
assign wcc = ~WCC;  //complement 
assign wgc = ~WGC;  //complement 
assign wgk = ~WGK;  //complement 
assign wck = ~WCK;  //complement 
assign QHC = ~qhc;  //complement 
assign odc = ~ODC;  //complement 
assign vdc = ~VDC;  //complement 
assign KDK =  WHK & TFD  |  VDK & TGD  ; 
assign kdk = ~KDK;  //complement 
assign JIC =  DAJ & dai & QJM  ; 
assign jic = ~JIC;  //complement  
assign JNC =  DAF & dae  ; 
assign jnc = ~JNC;  //complement 
assign odk = ~ODK;  //complement 
assign vdk = ~VDK;  //complement 
assign wdc = ~WDC;  //complement 
assign wdk = ~WDK;  //complement 
assign whc = ~WHC;  //complement 
assign whk = ~WHK;  //complement 
assign tac = ~TAC;  //complement 
assign tbc = ~TBC;  //complement 
assign tcc = ~TCC;  //complement 
assign tdc = ~TDC;  //complement 
assign agc = ~AGC;  //complement 
assign agk = ~AGK;  //complement 
assign ags = ~AGS;  //complement 
assign aek = ~AEK;  //complement 
assign aes = ~AES;  //complement 
assign acc = ~ACC;  //complement 
assign ack = ~ACK;  //complement 
assign acs = ~ACS;  //complement 
assign aac = ~AAC;  //complement 
assign aak = ~AAK;  //complement 
assign aas = ~AAS;  //complement 
assign ahc = ~AHC;  //complement 
assign ahk = ~AHK;  //complement 
assign ahs = ~AHS;  //complement 
assign afk = ~AFK;  //complement 
assign afs = ~AFS;  //complement 
assign aic = ~AIC;  //complement 
assign adc = ~ADC;  //complement 
assign adk = ~ADK;  //complement 
assign ads = ~ADS;  //complement 
assign aik = ~AIK;  //complement 
assign abc = ~ABC;  //complement 
assign abk = ~ABK;  //complement 
assign abs = ~ABS;  //complement 
assign ais = ~AIS;  //complement 
assign BDC =  AIC & ahc  |  aic & AHC  |  AIK & ahk  |  aik & AHK  |  AIS & ahs  |  ais & AHS  ;
assign bdc = ~BDC;  //complement 
assign BCC =  AIC & afc  |  aic & AFC  |  AIK & afk  |  aik & AFK  |  AIS & afs  |  ais & AFS  ;
assign bcc = ~BCC;  //complement 
assign BBC =  AIC & adc  |  aic & ADC  |  AIK & adk  |  aik & ADK  |  AIS & ads  |  ais & ADS  ;
assign bbc = ~BBC;  //complement 
assign BAC =  AIC & abc  |  aic & ABC  |  AIK & abk  |  aik & ABK  |  AIS & abs  |  ais & ABS  ;
assign bac = ~BAC;  //complement 
assign cca = ~CCA;  //complement 
assign caa = ~CAA;  //complement 
assign OEK = ~oek;  //complement 
assign OFK = ~ofk;  //complement 
assign OFC = ~ofc;  //complement 
assign okd = ~OKD;  //complement 
assign qjj = ~QJJ;  //complement 
assign OGC = ~ogc;  //complement 
assign OGK = ~ogk;  //complement 
assign OHC = ~ohc;  //complement 
assign qbc = ~QBC;  //complement 
assign qcc = ~QCC;  //complement 
assign qdk = ~QDK;  //complement 
assign qpc = ~QPC;  //complement 
assign OKO = ~oko;  //complement 
assign OKP = ~okp;  //complement 
assign OKQ = ~okq;  //complement 
assign pca = ~PCA;  //complement 
assign pcc = ~PCC;  //complement 
assign pce = ~PCE;  //complement 
assign pcb = ~PCB;  //complement 
assign pcd = ~PCD;  //complement 
assign pcf = ~PCF;  //complement 
assign JCA =  QPC  ; 
assign jca = ~JCA;  //complement 
assign JCB =  QPC & PCA  ; 
assign jcb = ~JCB;  //complement 
assign uma = ~UMA;  //complement 
assign una = ~UNA;  //complement 
assign umf = ~UMF;  //complement 
assign umg = ~UMG;  //complement 
assign umb = ~UMB;  //complement 
assign unb = ~UNB;  //complement 
assign ume = ~UME;  //complement 
assign une = ~UNE;  //complement 
assign umc = ~UMC;  //complement 
assign unc = ~UNC;  //complement 
assign unf = ~UNF;  //complement 
assign ung = ~UNG;  //complement 
assign umd = ~UMD;  //complement 
assign und = ~UND;  //complement 
assign uoa = ~UOA;  //complement 
assign upa = ~UPA;  //complement 
assign uof = ~UOF;  //complement 
assign uog = ~UOG;  //complement 
assign uob = ~UOB;  //complement 
assign upb = ~UPB;  //complement 
assign uoe = ~UOE;  //complement 
assign upe = ~UPE;  //complement 
assign uoc = ~UOC;  //complement 
assign upc = ~UPC;  //complement 
assign upf = ~UPF;  //complement 
assign upg = ~UPG;  //complement 
assign uod = ~UOD;  //complement 
assign upd = ~UPD;  //complement 
assign qdd = ~QDD;  //complement 
assign ted = ~TED;  //complement 
assign oad = ~OAD;  //complement 
assign vad = ~VAD;  //complement 
assign KAD =  WED & TFA  |  VAD & TGA  ; 
assign kad = ~KAD;  //complement 
assign KAL =  WEL & TFA  |  VAL & TGA  ; 
assign kal = ~KAL;  //complement 
assign oal = ~OAL;  //complement 
assign val = ~VAL;  //complement 
assign wad = ~WAD;  //complement 
assign wal = ~WAL;  //complement 
assign wed = ~WED;  //complement 
assign wel = ~WEL;  //complement 
assign obd = ~OBD;  //complement 
assign vbd = ~VBD;  //complement 
assign KDD =  WHD & TFD  |  VDD & TGD  ; 
assign kdd = ~KDD;  //complement 
assign KBD =  WFD & TFB  |  VBD & TGB  ; 
assign kbd = ~KBD;  //complement 
assign KBL =  WFL & TFB  |  VBL & TGB  ; 
assign kbl = ~KBL;  //complement 
assign wcl = ~WCL;  //complement 
assign obl = ~OBL;  //complement 
assign vbl = ~VBL;  //complement 
assign wbd = ~WBD;  //complement 
assign wbl = ~WBL;  //complement 
assign wfd = ~WFD;  //complement 
assign wfl = ~WFL;  //complement 
assign ocd = ~OCD;  //complement 
assign vcd = ~VCD;  //complement 
assign jdc =  qbd & qcd  ; 
assign JDC = ~jdc;  //complement 
assign KCD =  WGD & TFC  |  VCD & TGC  ; 
assign kcd = ~KCD;  //complement 
assign KCL =  WGL & TFC  |  VCL & TGC  ; 
assign kcl = ~KCL;  //complement 
assign qqd = ~QQD;  //complement 
assign ocl = ~OCL;  //complement 
assign vcl = ~VCL;  //complement 
assign wcd = ~WCD;  //complement 
assign wgd = ~WGD;  //complement 
assign wgl = ~WGL;  //complement 
assign QHD = ~qhd;  //complement 
assign odd = ~ODD;  //complement 
assign vdd = ~VDD;  //complement 
assign KDL =  WHL & TFD  |  VDL & TGD  ; 
assign kdl = ~KDL;  //complement 
assign JID =  DAJ & DAI & QJM  ; 
assign jid = ~JID;  //complement  
assign JND =  DAF & DAE  ; 
assign jnd = ~JND;  //complement 
assign odl = ~ODL;  //complement 
assign vdl = ~VDL;  //complement 
assign wdd = ~WDD;  //complement 
assign wdl = ~WDL;  //complement 
assign whd = ~WHD;  //complement 
assign whl = ~WHL;  //complement 
assign tad = ~TAD;  //complement 
assign tbd = ~TBD;  //complement 
assign tcd = ~TCD;  //complement 
assign tdd = ~TDD;  //complement 
assign agd = ~AGD;  //complement 
assign agl = ~AGL;  //complement 
assign agt = ~AGT;  //complement 
assign aed = ~AED;  //complement 
assign ael = ~AEL;  //complement 
assign aet = ~AET;  //complement 
assign acd = ~ACD;  //complement 
assign acl = ~ACL;  //complement 
assign act = ~ACT;  //complement 
assign aad = ~AAD;  //complement 
assign aal = ~AAL;  //complement 
assign aat = ~AAT;  //complement 
assign ahd = ~AHD;  //complement 
assign ahl = ~AHL;  //complement 
assign aht = ~AHT;  //complement 
assign afd = ~AFD;  //complement 
assign afl = ~AFL;  //complement 
assign aft = ~AFT;  //complement 
assign aid = ~AID;  //complement 
assign add = ~ADD;  //complement 
assign adt = ~ADT;  //complement 
assign ail = ~AIL;  //complement 
assign adl = ~ADL;  //complement 
assign abd = ~ABD;  //complement 
assign abl = ~ABL;  //complement 
assign abt = ~ABT;  //complement 
assign ait = ~AIT;  //complement 
assign BDD =  AID & ahd  |  aid & AHD  |  AIL & ahl  |  ail & AHL  |  AIT & aht  |  ait & AHR  ;
assign bdd = ~BDD;  //complement 
assign BCD =  AID & afd  |  aid & AFD  |  AIL & afl  |  ail & AFL  |  AIT & aft  |  ait & AFT  ;
assign bcd = ~BCD;  //complement 
assign BBD =  AID & add  |  aid & ADD  |  AIL & adl  |  ail & ADL  |  AIT & adt  |  ait & ADT  ;
assign bbd = ~BBD;  //complement 
assign BAD =  AID & abd  |  aid & ABD  |  AIL & abl  |  ail & ABL  |  AIT & abt  |  ait & ABT  ;
assign bad = ~BAD;  //complement 
assign cda = ~CDA;  //complement 
assign cba = ~CBA;  //complement 
assign OED = ~oed;  //complement 
assign OEL = ~oel;  //complement 
assign OFD = ~ofd;  //complement 
assign OFL = ~ofl;  //complement 
assign JJC =  cca & ccb  ; 
assign jjc = ~JJC;  //complement 
assign JJD =  cda & cdb  ; 
assign jjd = ~JJD;  //complement 
assign JJB =  cba & cbb  ; 
assign jjb = ~JJB;  //complement 
assign JJA =  caa & cab  ; 
assign jja = ~JJA;  //complement 
assign OGD = ~ogd;  //complement 
assign OGL = ~ogl;  //complement 
assign OHD = ~ohd;  //complement 
assign OHL = ~ohl;  //complement 
assign qeb = ~QEB;  //complement 
assign qbd = ~QBD;  //complement 
assign qcd = ~QCD;  //complement 
assign qdl = ~QDL;  //complement 
assign qpd = ~QPD;  //complement 
assign JDB =  QPD & PDA  ; 
assign jdb = ~JDB;  //complement 
assign OKR = ~okr;  //complement 
assign OKS = ~oks;  //complement 
assign OKT = ~okt;  //complement 
assign pda = ~PDA;  //complement 
assign pdc = ~PDC;  //complement 
assign pde = ~PDE;  //complement 
assign pdb = ~PDB;  //complement 
assign pdd = ~PDD;  //complement 
assign pdf = ~PDF;  //complement 
assign JDA =  QPD  ; 
assign jda = ~JDA;  //complement 
assign uai = ~UAI;  //complement 
assign ubi = ~UBI;  //complement 
assign uan = ~UAN;  //complement 
assign uao = ~UAO;  //complement 
assign ubn = ~UBN;  //complement 
assign ubo = ~UBO;  //complement 
assign uaj = ~UAJ;  //complement 
assign ubj = ~UBJ;  //complement 
assign uam = ~UAM;  //complement 
assign ubm = ~UBM;  //complement 
assign uak = ~UAK;  //complement 
assign ubk = ~UBK;  //complement 
assign obp = ~OBP;  //complement 
assign ual = ~UAL;  //complement 
assign ubl = ~UBL;  //complement 
assign uci = ~UCI;  //complement 
assign udi = ~UDI;  //complement 
assign ucn = ~UCN;  //complement 
assign uco = ~UCO;  //complement 
assign ucj = ~UCJ;  //complement 
assign udj = ~UDJ;  //complement 
assign ucm = ~UCM;  //complement 
assign udm = ~UDM;  //complement 
assign uck = ~UCK;  //complement 
assign udk = ~UDK;  //complement 
assign udn = ~UDN;  //complement 
assign udo = ~UDO;  //complement 
assign ucl = ~UCL;  //complement 
assign udl = ~UDL;  //complement 
assign tee = ~TEE;  //complement 
assign tde = ~TDE;  //complement 
assign oae = ~OAE;  //complement 
assign vae = ~VAE;  //complement 
assign KAE =  WEE & TFA  |  VAE & TGA  ; 
assign kae = ~KAE;  //complement 
assign KAM =  WEM & TFA  |  VAM & TGA  ; 
assign kam = ~KAM;  //complement 
assign oam = ~OAM;  //complement 
assign vam = ~VAM;  //complement 
assign wae = ~WAE;  //complement 
assign wam = ~WAM;  //complement 
assign wee = ~WEE;  //complement 
assign wem = ~WEM;  //complement 
assign obe = ~OBE;  //complement 
assign vbe = ~VBE;  //complement 
assign kde = ~KDE;  //complement 
assign KBE =  WFE & TFB  |  VBE & TGB  ; 
assign kbe = ~KBE;  //complement 
assign KBM =  WFM & TFB  |  VBM & TGB  ; 
assign kbm = ~KBM;  //complement 
assign obm = ~OBM;  //complement 
assign vbm = ~VBM;  //complement 
assign wbe = ~WBE;  //complement 
assign wbm = ~WBM;  //complement 
assign wfe = ~WFE;  //complement 
assign wfm = ~WFM;  //complement 
assign oce = ~OCE;  //complement 
assign vce = ~VCE;  //complement 
assign KCE =  WGE & TFC  |  VCE & TGC  ; 
assign kce = ~KCE;  //complement 
assign KCM =  WGM & TFC  |  VCM & TGC  ; 
assign kcm = ~KCM;  //complement 
assign ocm = ~OCM;  //complement 
assign vcm = ~VCM;  //complement 
assign wce = ~WCE;  //complement 
assign wcm = ~WCM;  //complement 
assign wge = ~WGE;  //complement 
assign wgm = ~WGM;  //complement 
assign hia = ~HIA;  //complement 
assign ode = ~ODE;  //complement 
assign vde = ~VDE;  //complement 
assign KDM =  WHM & TFD  |  VDM & TGD  ; 
assign kdm = ~KDM;  //complement 
assign jma =  daj & dai  ; 
assign JMA = ~jma;  //complement 
assign jmb =  daf  ; 
assign JMB = ~jmb;  //complement 
assign JMC =  DAJ & DAI  ; 
assign jmc = ~JMC;  //complement 
assign odm = ~ODM;  //complement 
assign vdm = ~VDM;  //complement 
assign wde = ~WDE;  //complement 
assign wdm = ~WDM;  //complement 
assign whe = ~WHE;  //complement 
assign whm = ~WHM;  //complement 
assign tae = ~TAE;  //complement 
assign tbe = ~TBE;  //complement 
assign tce = ~TCE;  //complement 
assign age = ~AGE;  //complement 
assign agm = ~AGM;  //complement 
assign agu = ~AGU;  //complement 
assign aee = ~AEE;  //complement 
assign aem = ~AEM;  //complement 
assign aeu = ~AEU;  //complement 
assign ace = ~ACE;  //complement 
assign acm = ~ACM;  //complement 
assign acu = ~ACU;  //complement 
assign aae = ~AAE;  //complement 
assign aam = ~AAM;  //complement 
assign aau = ~AAU;  //complement 
assign ahe = ~AHE;  //complement 
assign ahm = ~AHM;  //complement 
assign ahu = ~AHU;  //complement 
assign afe = ~AFE;  //complement 
assign afm = ~AFM;  //complement 
assign afu = ~AFU;  //complement 
assign aie = ~AIE;  //complement 
assign ade = ~ADE;  //complement 
assign adm = ~ADM;  //complement 
assign adu = ~ADU;  //complement 
assign aim = ~AIM;  //complement 
assign abe = ~ABE;  //complement 
assign abm = ~ABM;  //complement 
assign abu = ~ABU;  //complement 
assign aiu = ~AIU;  //complement 
assign BDE =  AIE & ahe  |  aie & AHE  |  AIM & ahm  |  aim & AHM  |  AIU & ahu  |  aiu & AHU  ;
assign bde = ~BDE;  //complement 
assign JHA =  DAC  ; 
assign jha = ~JHA;  //complement 
assign JHB =  DAD  ; 
assign jhb = ~JHB;  //complement 
assign BBE =  AIE & ade  |  aie & ADE  |  AIM & adm  |  aim & ADM  |  AIU & adu  |  aiu & ADU  ;
assign bbe = ~BBE;  //complement 
assign BAE =  AIE & abe  |  aie & ABE  |  AIM & abm  |  aim & ABM  |  AIU & abu  |  aiu & ABU  ;
assign bae = ~BAE;  //complement 
assign ccb = ~CCB;  //complement 
assign cab = ~CAB;  //complement 
assign OEE = ~oee;  //complement 
assign OEM = ~oem;  //complement 
assign OFE = ~ofe;  //complement 
assign OFM = ~ofm;  //complement 
assign eaa = ~EAA;  //complement 
assign eab = ~EAB;  //complement 
assign OGE = ~oge;  //complement 
assign OGM = ~ogm;  //complement 
assign OHE = ~ohe;  //complement 
assign OHM = ~ohm;  //complement 
assign JKA =  HIA & QFA  ; 
assign jka = ~JKA;  //complement 
assign eac = ~EAC;  //complement 
assign ead = ~EAD;  //complement 
assign JED =  qla & DAA & DAB & DAC  ; 
assign jed = ~JED;  //complement  
assign JEE =  DAA & DAB & DAC & DAD  ; 
assign jee = ~JEE;  //complement 
assign JEA =  qla  ; 
assign jea = ~JEA;  //complement 
assign JEC =  qla & DAA & DAB  ; 
assign jec = ~JEC;  //complement 
assign JEB =  qla & DAA & DAB  ; 
assign jeb = ~JEB;  //complement 
assign BCE =  AIE & afe  |  aie & AFE  |  AIM & afm  |  aim & AFM  |  AIU & afu  |  aiu & AFU  ;
assign bce = ~BCE;  //complement 
assign daa = ~DAA;  //complement 
assign dae = ~DAE;  //complement 
assign dai = ~DAI;  //complement 
assign dab = ~DAB;  //complement 
assign daf = ~DAF;  //complement 
assign daj = ~DAJ;  //complement 
assign dac = ~DAC;  //complement 
assign dag = ~DAG;  //complement 
assign dak = ~DAK;  //complement 
assign dad = ~DAD;  //complement 
assign dah = ~DAH;  //complement 
assign dal = ~DAL;  //complement 
assign uei = ~UEI;  //complement 
assign ufi = ~UFI;  //complement 
assign uen = ~UEN;  //complement 
assign ueo = ~UEO;  //complement 
assign uej = ~UEJ;  //complement 
assign ufj = ~UFJ;  //complement 
assign uem = ~UEM;  //complement 
assign ufm = ~UFM;  //complement 
assign ufk = ~UFK;  //complement 
assign uek = ~UEK;  //complement 
assign ufn = ~UFN;  //complement 
assign ufo = ~UFO;  //complement 
assign uel = ~UEL;  //complement 
assign ufl = ~UFL;  //complement 
assign ugi = ~UGI;  //complement 
assign uhi = ~UHI;  //complement 
assign ugn = ~UGN;  //complement 
assign ugo = ~UGO;  //complement 
assign ugj = ~UGJ;  //complement 
assign uhj = ~UHJ;  //complement 
assign ugm = ~UGM;  //complement 
assign uhm = ~UHM;  //complement 
assign ugk = ~UGK;  //complement 
assign uhk = ~UHK;  //complement 
assign uhn = ~UHN;  //complement 
assign uho = ~UHO;  //complement 
assign ugl = ~UGL;  //complement 
assign uhl = ~UHL;  //complement 
assign tef = ~TEF;  //complement 
assign oaf = ~OAF;  //complement 
assign vaf = ~VAF;  //complement 
assign KAF =  WEF & TFA  |  VAF & TGA  ; 
assign kaf = ~KAF;  //complement 
assign KAN =  WEN & TFA  |  VAN & TGA  ; 
assign kan = ~KAN;  //complement 
assign tfa = ~TFA;  //complement 
assign TGA = ~tga;  //complement 
assign oan = ~OAN;  //complement 
assign van = ~VAN;  //complement 
assign waf = ~WAF;  //complement 
assign wan = ~WAN;  //complement 
assign wef = ~WEF;  //complement 
assign wen = ~WEN;  //complement 
assign obf = ~OBF;  //complement 
assign vbf = ~VBF;  //complement 
assign KDF =  WHF & TFD  |  VDF & TGD  ; 
assign kdf = ~KDF;  //complement 
assign KBF =  WFF & TFB  |  VBF & TGB  ; 
assign kbf = ~KBF;  //complement 
assign KBN =  WFN & TFB  |  VBN & TGB  ; 
assign kbn = ~KBN;  //complement 
assign tfb = ~TFB;  //complement 
assign TGB = ~tgb;  //complement 
assign obn = ~OBN;  //complement 
assign vbn = ~VBN;  //complement 
assign wbf = ~WBF;  //complement 
assign wbn = ~WBN;  //complement 
assign wff = ~WFF;  //complement 
assign wfn = ~WFN;  //complement 
assign ocf = ~OCF;  //complement 
assign vcf = ~VCF;  //complement 
assign KCF =  WGF & TFC  |  VCF & TGC  ; 
assign kcf = ~KCF;  //complement 
assign KCN =  WGN & TFC  |  VCN & TGC  ; 
assign kcn = ~KCN;  //complement 
assign tfc = ~TFC;  //complement 
assign TGC = ~tgc;  //complement 
assign ocn = ~OCN;  //complement 
assign vcn = ~VCN;  //complement 
assign wcf = ~WCF;  //complement 
assign wcn = ~WCN;  //complement 
assign wgf = ~WGF;  //complement 
assign wgn = ~WGN;  //complement 
assign hib = ~HIB;  //complement 
assign odf = ~ODF;  //complement 
assign vdf = ~VDF;  //complement 
assign KDN =  WHN & TFD  |  VDN & TGD  ; 
assign kdn = ~KDN;  //complement 
assign tfd = ~TFD;  //complement 
assign TGD = ~tgd;  //complement 
assign odn = ~ODN;  //complement 
assign vdn = ~VDN;  //complement 
assign wdf = ~WDF;  //complement 
assign wdn = ~WDN;  //complement 
assign whf = ~WHF;  //complement 
assign whn = ~WHN;  //complement 
assign taf = ~TAF;  //complement 
assign tbf = ~TBF;  //complement 
assign tcf = ~TCF;  //complement 
assign tdf = ~TDF;  //complement 
assign agf = ~AGF;  //complement 
assign agn = ~AGN;  //complement 
assign agv = ~AGV;  //complement 
assign aef = ~AEF;  //complement 
assign aen = ~AEN;  //complement 
assign aev = ~AEV;  //complement 
assign OKI = ~oki;  //complement 
assign acf = ~ACF;  //complement 
assign acn = ~ACN;  //complement 
assign acv = ~ACV;  //complement 
assign aaf = ~AAF;  //complement 
assign aan = ~AAN;  //complement 
assign aav = ~AAV;  //complement 
assign ahf = ~AHF;  //complement 
assign ahn = ~AHN;  //complement 
assign ahv = ~AHV;  //complement 
assign aff = ~AFF;  //complement 
assign afn = ~AFN;  //complement 
assign afv = ~AFV;  //complement 
assign aif = ~AIF;  //complement 
assign adf = ~ADF;  //complement 
assign adn = ~ADN;  //complement 
assign adv = ~ADV;  //complement 
assign ain = ~AIN;  //complement 
assign abf = ~ABF;  //complement 
assign abn = ~ABN;  //complement 
assign abv = ~ABV;  //complement 
assign aiv = ~AIV;  //complement 
assign BCF =  AIF & aff  |  aif & AFF  |  AIN & afn  |  ain & AFN  |  AIV & afv  |  aiv & AFV  ;
assign bcf = ~BCF;  //complement 
assign EBC = ~ebc;  //complement 
assign BBF =  AIF & adf  |  aif & ADF  |  AIN & adn  |  ain & ADN  |  AIV & adv  |  aiv & ADV  ;
assign bbf = ~BBF;  //complement 
assign BAF =  AIF & abf  |  aif & ABF  |  AIN & abn  |  ain & ABN  |  AIV & abv  |  aiv & ABV  ;
assign baf = ~BAF;  //complement 
assign qjp = ~QJP;  //complement 
assign cdb = ~CDB;  //complement 
assign cbb = ~CBB;  //complement 
assign OEF = ~oef;  //complement 
assign OEN = ~oen;  //complement 
assign OFF = ~off;  //complement 
assign OFN = ~ofn;  //complement 
assign okh = ~OKH;  //complement 
assign qjd = ~QJD;  //complement 
assign QEC = ~qec;  //complement 
assign QED = ~qed;  //complement 
assign qjf = ~QJF;  //complement 
assign OGF = ~ogf;  //complement 
assign OGN = ~ogn;  //complement 
assign OHF = ~ohf;  //complement 
assign OHN = ~ohn;  //complement 
assign JKB =  HIB & QFA  ; 
assign jkb = ~JKB;  //complement 
assign JOA =  QJD & QJF  ; 
assign joa = ~JOA;  //complement 
assign JQA =  QJA  ; 
assign jqa = ~JQA;  //complement 
assign oka = ~OKA;  //complement 
assign qjm = ~QJM;  //complement 
assign qjn = ~QJN;  //complement 
assign oke = ~OKE;  //complement 
assign qjc = ~QJC;  //complement 
assign qje = ~QJE;  //complement 
assign qjg = ~QJG;  //complement 
assign EBA = ~eba;  //complement 
assign EBB = ~ebb;  //complement 
assign BDF =  AIF & ahf  |  aif & AHF  |  AIN & ahn  |  ain & AHN  |  AIV & ahv  |  aiv & AHV  ;
assign bdf = ~BDF;  //complement 
assign QLA = ~qla;  //complement 
assign QLB = ~qlb;  //complement 
assign dba = ~DBA;  //complement 
assign dbe = ~DBE;  //complement 
assign dbi = ~DBI;  //complement 
assign dbb = ~DBB;  //complement 
assign dbf = ~DBF;  //complement 
assign dbj = ~DBJ;  //complement 
assign dbc = ~DBC;  //complement 
assign dbg = ~DBG;  //complement 
assign dbk = ~DBK;  //complement 
assign QLC = ~qlc;  //complement 
assign QLE = ~qle;  //complement 
assign uii = ~UII;  //complement 
assign uji = ~UJI;  //complement 
assign uin = ~UIN;  //complement 
assign uio = ~UIO;  //complement 
assign uij = ~UIJ;  //complement 
assign ujj = ~UJJ;  //complement 
assign uim = ~UIM;  //complement 
assign ujm = ~UJM;  //complement 
assign uik = ~UIK;  //complement 
assign ujk = ~UJK;  //complement 
assign ujn = ~UJN;  //complement 
assign ujo = ~UJO;  //complement 
assign uil = ~UIL;  //complement 
assign ujl = ~UJL;  //complement 
assign uki = ~UKI;  //complement 
assign uli = ~ULI;  //complement 
assign ukn = ~UKN;  //complement 
assign uko = ~UKO;  //complement 
assign ukj = ~UKJ;  //complement 
assign ulj = ~ULJ;  //complement 
assign ukm = ~UKM;  //complement 
assign ulm = ~ULM;  //complement 
assign ukk = ~UKK;  //complement 
assign ulk = ~ULK;  //complement 
assign uln = ~ULN;  //complement 
assign ulo = ~ULO;  //complement 
assign ukl = ~UKL;  //complement 
assign ull = ~ULL;  //complement 
assign teg = ~TEG;  //complement 
assign oag = ~OAG;  //complement 
assign vag = ~VAG;  //complement 
assign KAG =  WEG & TFA  |  VAG & TGA  ; 
assign kag = ~KAG;  //complement 
assign KAO =  WEO & TFA  |  VAO & TGA  ; 
assign kao = ~KAO;  //complement 
assign faa = ~FAA;  //complement 
assign oao = ~OAO;  //complement 
assign vao = ~VAO;  //complement 
assign wag = ~WAG;  //complement 
assign wao = ~WAO;  //complement 
assign weg = ~WEG;  //complement 
assign weo = ~WEO;  //complement 
assign fab = ~FAB;  //complement 
assign obg = ~OBG;  //complement 
assign vbg = ~VBG;  //complement 
assign KDG =  WHG & TFD  |  VDG & TGD  ; 
assign kdg = ~KDG;  //complement 
assign KBG =  WFG & TFB  |  VBG & TGB  ; 
assign kbg = ~KBG;  //complement 
assign KBO =  WFO & TFB  |  VBO & TGB  ; 
assign kbo = ~KBO;  //complement 
assign fac = ~FAC;  //complement 
assign obo = ~OBO;  //complement 
assign vbo = ~VBO;  //complement 
assign wbg = ~WBG;  //complement 
assign wbo = ~WBO;  //complement 
assign wfg = ~WFG;  //complement 
assign wfo = ~WFO;  //complement 
assign fad = ~FAD;  //complement 
assign ocg = ~OCG;  //complement 
assign vcg = ~VCG;  //complement 
assign KCG =  WGG & TFC  |  VCG & TGC  ; 
assign kcg = ~KCG;  //complement 
assign KCO =  WGO & TFC  |  VCO & TGC  ; 
assign kco = ~KCO;  //complement 
assign OHK = ~ohk;  //complement 
assign oco = ~OCO;  //complement 
assign vco = ~VCO;  //complement 
assign wcg = ~WCG;  //complement 
assign wco = ~WCO;  //complement 
assign wgg = ~WGG;  //complement 
assign wgo = ~WGO;  //complement 
assign hic = ~HIC;  //complement 
assign odg = ~ODG;  //complement 
assign vdg = ~VDG;  //complement 
assign KDO =  WHO & TFD  |  VDO & TGD  ; 
assign kdo = ~KDO;  //complement 
assign qpe = ~QPE;  //complement 
assign odo = ~ODO;  //complement 
assign vdo = ~VDO;  //complement 
assign wdg = ~WDG;  //complement 
assign wdo = ~WDO;  //complement 
assign whg = ~WHG;  //complement 
assign who = ~WHO;  //complement 
assign tag = ~TAG;  //complement 
assign tbg = ~TBG;  //complement 
assign tcg = ~TCG;  //complement 
assign tdg = ~TDG;  //complement 
assign agg = ~AGG;  //complement 
assign ago = ~AGO;  //complement 
assign agw = ~AGW;  //complement 
assign aeg = ~AEG;  //complement 
assign aeo = ~AEO;  //complement 
assign aew = ~AEW;  //complement 
assign acg = ~ACG;  //complement 
assign aco = ~ACO;  //complement 
assign acw = ~ACW;  //complement 
assign aag = ~AAG;  //complement 
assign aao = ~AAO;  //complement 
assign aaw = ~AAW;  //complement 
assign ahg = ~AHG;  //complement 
assign aho = ~AHO;  //complement 
assign ahw = ~AHW;  //complement 
assign afg = ~AFG;  //complement 
assign afo = ~AFO;  //complement 
assign afw = ~AFW;  //complement 
assign aig = ~AIG;  //complement 
assign adg = ~ADG;  //complement 
assign ado = ~ADO;  //complement 
assign adw = ~ADW;  //complement 
assign aio = ~AIO;  //complement 
assign abg = ~ABG;  //complement 
assign abo = ~ABO;  //complement 
assign abw = ~ABW;  //complement 
assign aiw = ~AIW;  //complement 
assign BDG =  AIG & ahg  |  aig & AHG  |  AIO & aho  |  aio & AHO  |  AIW & ahw  |  aiw & AHW  ;
assign bdg = ~BDG;  //complement 
assign BCG =  AIG & afg  |  aig & AFG  |  AIO & afo  |  aio & AFO  |  AIW & afw  |  aiw & AFW  ;
assign bcg = ~BCG;  //complement 
assign BBG =  AIG & adg  |  aig & ADG  |  AIO & ado  |  aio & ADO  |  AIW & adw  |  aiw & ADW  ;
assign bbg = ~BBG;  //complement 
assign BAG =  AIG & abg  |  aig & ABG  |  AIO & abo  |  aio & ABO  |  AIW & abw  |  aiw & ABW  ;
assign bag = ~BAG;  //complement 
assign JLA =  QDE  ; 
assign jla = ~JLA;  //complement 
assign JLC =  QDE & FAA & FAB  ; 
assign jlc = ~JLC;  //complement 
assign JLB =  QDE & FAA & FAB  ; 
assign jlb = ~JLB;  //complement 
assign OEG = ~oeg;  //complement 
assign OEO = ~oeo;  //complement 
assign OFG = ~ofg;  //complement 
assign OFO = ~ofo;  //complement 
assign JLE =  QDE & FAA & FAB & FAC & FAD  ; 
assign jle = ~JLE;  //complement  
assign JLD =  QDE & FAA & FAB & FAC  ; 
assign jld = ~JLD;  //complement 
assign JPB =  QJF & qed & qja & qjd & qjn & qjp  ; 
assign jpb = ~JPB;  //complement  
assign JPC =  qha & qhb & qhc & qhd & qlh  ; 
assign jpc = ~JPC;  //complement  
assign OGG = ~ogg;  //complement 
assign OGO = ~ogo;  //complement 
assign OHG = ~ohg;  //complement 
assign OHO = ~oho;  //complement 
assign jpe =  qeb & qed  ; 
assign JPE = ~jpe;  //complement 
assign JQB =  QJA  ; 
assign jqb = ~JQB;  //complement 
assign JKC =  HIC & QFA  ; 
assign jkc = ~JKC;  //complement 
assign jpf =  qeb & qed  ; 
assign JPF = ~jpf;  //complement 
assign OKF = ~okf;  //complement 
assign okg = ~OKG;  //complement 
assign qja = ~QJA;  //complement 
assign qjb = ~QJB;  //complement 
assign oja = ~OJA;  //complement 
assign ojb = ~OJB;  //complement 
assign OJD = ~ojd;  //complement 
assign OJE = ~oje;  //complement 
assign jfb =  PEA & dba  |  pea & DBA  |  PEB & dbb  |  peb & DBB  |  PEC & dbc  |  pec & DBC  ;
assign JFB = ~jfb;  //complement 
assign jfa =  PEA & hea  |  pea & HEA  |  PEB & heb  |  peb & HEB  |  PEC & hec  |  pec & HEC  ;
assign JFA = ~jfa;  //complement 
assign JGA =  QPE  ; 
assign jga = ~JGA;  //complement 
assign JGC =  QPE & PEA & PEB  ; 
assign jgc = ~JGC;  //complement 
assign JGB =  QPE & PEA & PEB  ; 
assign jgb = ~JGB;  //complement 
assign qlg = ~QLG;  //complement 
assign qlh = ~QLH;  //complement 
assign pea = ~PEA;  //complement 
assign pfa = ~PFA;  //complement 
assign pga = ~PGA;  //complement 
assign peb = ~PEB;  //complement 
assign pfb = ~PFB;  //complement 
assign pgb = ~PGB;  //complement 
assign pec = ~PEC;  //complement 
assign pfc = ~PFC;  //complement 
assign pgc = ~PGC;  //complement 
assign qld = ~QLD;  //complement 
assign qlf = ~QLF;  //complement 
assign umi = ~UMI;  //complement 
assign uni = ~UNI;  //complement 
assign umn = ~UMN;  //complement 
assign umo = ~UMO;  //complement 
assign umj = ~UMJ;  //complement 
assign unj = ~UNJ;  //complement 
assign umm = ~UMM;  //complement 
assign unm = ~UNM;  //complement 
assign umk = ~UMK;  //complement 
assign unk = ~UNK;  //complement 
assign unn = ~UNN;  //complement 
assign uno = ~UNO;  //complement 
assign uml = ~UML;  //complement 
assign unl = ~UNL;  //complement 
assign gab = ~GAB;  //complement 
assign uoi = ~UOI;  //complement 
assign upi = ~UPI;  //complement 
assign uon = ~UON;  //complement 
assign uoo = ~UOO;  //complement 
assign uoj = ~UOJ;  //complement 
assign upj = ~UPJ;  //complement 
assign uom = ~UOM;  //complement 
assign upm = ~UPM;  //complement 
assign uok = ~UOK;  //complement 
assign upk = ~UPK;  //complement 
assign upn = ~UPN;  //complement 
assign upo = ~UPO;  //complement 
assign uol = ~UOL;  //complement 
assign upl = ~UPL;  //complement 
assign teh = ~TEH;  //complement 
assign oah = ~OAH;  //complement 
assign vah = ~VAH;  //complement 
assign KAH =  WEH & TFA  |  VAH & TGA  ; 
assign kah = ~KAH;  //complement 
assign KAP =  WEP & TFA  |  VAP & TGA  ; 
assign kap = ~KAP;  //complement 
assign JRA =  GAA & GAB  ; 
assign jra = ~JRA;  //complement 
assign oap = ~OAP;  //complement 
assign vap = ~VAP;  //complement 
assign wah = ~WAH;  //complement 
assign wap = ~WAP;  //complement 
assign weh = ~WEH;  //complement 
assign wep = ~WEP;  //complement 
assign gaa = ~GAA;  //complement 
assign obh = ~OBH;  //complement 
assign vbh = ~VBH;  //complement 
assign KDH =  WHH & TFD  |  VDH & TGD  ; 
assign kdh = ~KDH;  //complement 
assign KBH =  WFH & TFB  |  VBH & TGB  ; 
assign kbh = ~KBH;  //complement 
assign KBP =  WFP & TFB  |  VBP & TGB  ; 
assign kbp = ~KBP;  //complement 
assign vbp = ~VBP;  //complement 
assign wch = ~WCH;  //complement 
assign wbh = ~WBH;  //complement 
assign wbp = ~WBP;  //complement 
assign wfh = ~WFH;  //complement 
assign wfp = ~WFP;  //complement 
assign och = ~OCH;  //complement 
assign vch = ~VCH;  //complement 
assign KCH =  WGH & TFC  |  VCH & TGC  ; 
assign kch = ~KCH;  //complement 
assign KCP =  WGP & TFC  |  VCP & TGC  ; 
assign kcp = ~KCP;  //complement 
assign ocp = ~OCP;  //complement 
assign vcp = ~VCP;  //complement 
assign wgh = ~WGH;  //complement 
assign wgp = ~WGP;  //complement 
assign wcp = ~WCP;  //complement 
assign hid = ~HID;  //complement 
assign ojc = ~OJC;  //complement 
assign odh = ~ODH;  //complement 
assign vdh = ~VDH;  //complement 
assign gac = ~GAC;  //complement 
assign KDP =  WHP & TFD  |  VDP & TGD  ; 
assign kdp = ~KDP;  //complement 
assign tja = ~TJA;  //complement 
assign tjb = ~TJB;  //complement 
assign tjc = ~TJC;  //complement 
assign tjd = ~TJD;  //complement 
assign odp = ~ODP;  //complement 
assign vdp = ~VDP;  //complement 
assign wdh = ~WDH;  //complement 
assign wdp = ~WDP;  //complement 
assign whh = ~WHH;  //complement 
assign whp = ~WHP;  //complement 
assign tah = ~TAH;  //complement 
assign tbh = ~TBH;  //complement 
assign tch = ~TCH;  //complement 
assign tdh = ~TDH;  //complement 
assign agh = ~AGH;  //complement 
assign agp = ~AGP;  //complement 
assign agx = ~AGX;  //complement 
assign aeh = ~AEH;  //complement 
assign aep = ~AEP;  //complement 
assign aex = ~AEX;  //complement 
assign OKU = ~oku;  //complement 
assign ach = ~ACH;  //complement 
assign acp = ~ACP;  //complement 
assign acx = ~ACX;  //complement 
assign OKV = ~okv;  //complement 
assign aah = ~AAH;  //complement 
assign aap = ~AAP;  //complement 
assign aax = ~AAX;  //complement 
assign ahh = ~AHH;  //complement 
assign ahp = ~AHP;  //complement 
assign ahx = ~AHX;  //complement 
assign afh = ~AFH;  //complement 
assign afp = ~AFP;  //complement 
assign afx = ~AFX;  //complement 
assign aih = ~AIH;  //complement 
assign adh = ~ADH;  //complement 
assign adp = ~ADP;  //complement 
assign adx = ~ADX;  //complement 
assign aip = ~AIP;  //complement 
assign abh = ~ABH;  //complement 
assign abp = ~ABP;  //complement 
assign abx = ~ABX;  //complement 
assign aix = ~AIX;  //complement 
assign BDH =  AIH & ahh  |  aih & AHH  |  AIP & ahp  |  aip & AHP  |  AIX & ahx  |  aix & AHX  ;
assign bdh = ~BDH;  //complement 
assign BCH =  AIH & afh  |  aih & AFH  |  AIP & afp  |  aip & AFP  |  AIX & afx  |  aix & AFX  ;
assign bch = ~BCH;  //complement 
assign BBH =  AIH & adh  |  aih & ADH  |  AIP & adp  |  aip & ADP  |  AIX & adx  |  aix & ADX  ;
assign bbh = ~BBH;  //complement 
assign BAH =  AIH & abh  |  aih & ABH  |  AIP & abp  |  aip & ABP  |  AIX & abx  |  aix & ABX  ;
assign bah = ~BAH;  //complement 
assign haa = ~HAA;  //complement 
assign hba = ~HBA;  //complement 
assign hca = ~HCA;  //complement 
assign hda = ~HDA;  //complement 
assign hab = ~HAB;  //complement 
assign hbb = ~HBB;  //complement 
assign hcb = ~HCB;  //complement 
assign hdb = ~HDB;  //complement 
assign hac = ~HAC;  //complement 
assign hbc = ~HBC;  //complement 
assign hcc = ~HCC;  //complement 
assign hdc = ~HDC;  //complement 
assign OEH = ~oeh;  //complement 
assign OEP = ~oep;  //complement 
assign OFH = ~ofh;  //complement 
assign OFP = ~ofp;  //complement 
assign hea = ~HEA;  //complement 
assign hfa = ~HFA;  //complement 
assign hga = ~HGA;  //complement 
assign hha = ~HHA;  //complement 
assign heb = ~HEB;  //complement 
assign hfb = ~HFB;  //complement 
assign hgb = ~HGB;  //complement 
assign hhb = ~HHB;  //complement 
assign hec = ~HEC;  //complement 
assign hfc = ~HFC;  //complement 
assign hgc = ~HGC;  //complement 
assign hhc = ~HHC;  //complement 
assign OGH = ~ogh;  //complement 
assign OGP = ~ogp;  //complement 
assign OHH = ~ohh;  //complement 
assign OHP = ~ohp;  //complement 
assign JKD =  HID & QFA  ; 
assign jkd = ~JKD;  //complement 
assign qfa = ~QFA;  //complement 
assign tma = ~TMA;  //complement 
assign qkb = ~QKB;  //complement 
assign OKW = ~okw;  //complement 
assign OKX = ~okx;  //complement 
assign qka = ~QKA;  //complement 
assign iaa = ~IAA; //complement 
assign iab = ~IAB; //complement 
assign iac = ~IAC; //complement 
assign iad = ~IAD; //complement 
assign iae = ~IAE; //complement 
assign iaf = ~IAF; //complement 
assign iag = ~IAG; //complement 
assign iah = ~IAH; //complement 
assign iai = ~IAI; //complement 
assign iaj = ~IAJ; //complement 
assign iak = ~IAK; //complement 
assign ial = ~IAL; //complement 
assign iam = ~IAM; //complement 
assign ian = ~IAN; //complement 
assign iao = ~IAO; //complement 
assign iap = ~IAP; //complement 
assign iba = ~IBA; //complement 
assign ibb = ~IBB; //complement 
assign ibc = ~IBC; //complement 
assign ibd = ~IBD; //complement 
assign ibe = ~IBE; //complement 
assign ibf = ~IBF; //complement 
assign ibg = ~IBG; //complement 
assign ibh = ~IBH; //complement 
assign ibi = ~IBI; //complement 
assign ibj = ~IBJ; //complement 
assign ibk = ~IBK; //complement 
assign ibl = ~IBL; //complement 
assign ibm = ~IBM; //complement 
assign ibn = ~IBN; //complement 
assign ibo = ~IBO; //complement 
assign ibp = ~IBP; //complement 
assign ica = ~ICA; //complement 
assign icb = ~ICB; //complement 
assign icc = ~ICC; //complement 
assign icd = ~ICD; //complement 
assign ice = ~ICE; //complement 
assign icf = ~ICF; //complement 
assign icg = ~ICG; //complement 
assign ich = ~ICH; //complement 
assign ici = ~ICI; //complement 
assign icj = ~ICJ; //complement 
assign ick = ~ICK; //complement 
assign icl = ~ICL; //complement 
assign icm = ~ICM; //complement 
assign icn = ~ICN; //complement 
assign ico = ~ICO; //complement 
assign icp = ~ICP; //complement 
assign ida = ~IDA; //complement 
assign idb = ~IDB; //complement 
assign idc = ~IDC; //complement 
assign idd = ~IDD; //complement 
assign ide = ~IDE; //complement 
assign idf = ~IDF; //complement 
assign idg = ~IDG; //complement 
assign idh = ~IDH; //complement 
assign idi = ~IDI; //complement 
assign idj = ~IDJ; //complement 
assign idk = ~IDK; //complement 
assign idl = ~IDL; //complement 
assign idm = ~IDM; //complement 
assign idn = ~IDN; //complement 
assign ido = ~IDO; //complement 
assign idp = ~IDP; //complement 
assign iea = ~IEA; //complement 
assign ieb = ~IEB; //complement 
assign iec = ~IEC; //complement 
assign ied = ~IED; //complement 
assign iee = ~IEE; //complement 
assign ief = ~IEF; //complement 
assign ieg = ~IEG; //complement 
assign ieh = ~IEH; //complement 
assign iei = ~IEI; //complement 
assign iej = ~IEJ; //complement 
assign iek = ~IEK; //complement 
assign iel = ~IEL; //complement 
assign iem = ~IEM; //complement 
assign ien = ~IEN; //complement 
assign ieo = ~IEO; //complement 
assign iep = ~IEP; //complement 
assign ieq = ~IEQ; //complement 
assign ier = ~IER; //complement 
assign ies = ~IES; //complement 
assign iet = ~IET; //complement 
assign ieu = ~IEU; //complement 
assign iev = ~IEV; //complement 
assign iew = ~IEW; //complement 
assign iex = ~IEX; //complement 
assign ifa = ~IFA; //complement 
assign ifb = ~IFB; //complement 
assign ifc = ~IFC; //complement 
assign ifd = ~IFD; //complement 
assign iga = ~IGA; //complement 
assign igb = ~IGB; //complement 
assign igc = ~IGC; //complement 
assign iha = ~IHA; //complement 
assign ihb = ~IHB; //complement 
assign ijb = ~IJB; //complement 
assign ijd = ~IJD; //complement 
assign ije = ~IJE; //complement 
assign ijf = ~IJF; //complement 
always@(posedge IZZ )
   begin 
 UAA <=  PAC & TEA  |  DAG & tea  ; 
 UBA <=  PAC & TEA  |  DAG & tea  ; 
 UAF <= QDA ; 
 UAG <= QDA ; 
 UBF <= QDA ; 
 UBG <= QDA ; 
 UAB <=  PAD & TEA  |  DAH & tea  ; 
 UBB <=  PAD & TEA  |  DAH & tea  ; 
 UAE <=  PFC & TEA  |  DBG & tea  ; 
 UBE <=  PFC & TEA  |  DBG & tea  ; 
 UAC <=  PFA & TEA  |  DBE & tea  ; 
 UBC <=  PFA & TEA  |  DBE & tea  ; 
 UAD <=  PFB & TEA  |  DBF & tea  ; 
 UBD <=  PFB & TEA  |  DBF & tea  ; 
 UCE <=  PGC & TEA  |  DBK & tea  ; 
 UDE <=  PGC & TEA  |  DBK & tea  ; 
 UCA <=  PAC & TEA  |  DAK & tea  ; 
 UDA <=  PAC & TEA  |  DAK & tea  ; 
 UCF <= QDA ; 
 UCG <= QDA ; 
 UCB <=  PAD & TEA  |  DAL & tea  ; 
 UDB <=  PAD & TEA  |  DAL & tea  ; 
 UCC <=  PGA & TEA  |  DBI & tea  ; 
 UDC <=  PGA & TEA  |  DBI & tea  ; 
 UDF <= QDA ; 
 UDG <= QDA ; 
 UCD <=  PGB & TEA  |  DBJ & tea  ; 
 UDD <=  PGB & TEA  |  DBJ & tea  ; 
 QDA <= QCA ; 
 TEA <= JAC ; 
 OAA <=  RAA & TAA  |  REA & TBA  |  RIA & TCA  |  RMA & TDA  |  KAA  ; 
 VAA <=  RAA & TAA  |  REA & TBA  |  RIA & TCA  |  RMA & TDA  |  KAA  ; 
 OAI <=  RAI & TAB  |  REI & TBB  |  RII & TCB  |  RMI & TDB  |  KAI  ; 
 VAI <=  RAI & TAB  |  REI & TBB  |  RII & TCB  |  RMI & TDB  |  KAI  ; 
 WAA <= IAA ; 
 WAI <= IAI ; 
 WEA <= IAA ; 
 WEI <= IAI ; 
 OBA <=  RBA & TAC  |  RFA & TBC  |  RJA & TCC  |  RNA & TDC  |  KBA  ; 
 VBA <=  RBA & TAC  |  RFA & TBC  |  RJA & TCC  |  RNA & TDC  |  KBA  ; 
 OBI <=  RBI & TAD  |  RFI & TBD  |  RJI & TCD  |  RNI & TDD  |  KBI  ; 
 VBI <=  RBI & TAD  |  RFI & TBD  |  RJI & TCD  |  RNI & TDD  |  KBI  ; 
 WBA <= IBA ; 
 WBI <= IBI ; 
 WFA <= IBA ; 
 WFI <= IBI ; 
 OCA <=  RCA & TAE  |  RGA & TBE  |  RKA & TCE  |  ROA & TDE  |  KCA  ; 
 VCA <=  RCA & TAE  |  RGA & TBE  |  RKA & TCE  |  ROA & TDE  |  KCA  ; 
 QQA <=  QQA & jqb  |  QDI  ; 
 OCI <=  RCI & TAF  |  RGI & TBF  |  RKI & TCF  |  ROI & TDF  |  KCI  ; 
 VCI <=  RCI & TAF  |  RGI & TBF  |  RKI & TCF  |  ROI & TDF  |  KCI  ; 
 WCA <= ICA ; 
 WCI <= ICI ; 
 WGA <= ICA ; 
 WGI <= ICI ; 
 qha <=  qaa & qba & qca  |  jna  ; 
 ODA <=  RDA & TAG  |  RHA & TBG  |  RLA & TCG  |  RPA & TDG  |  KDA  ; 
 VDA <=  RDA & TAG  |  RHA & TBG  |  RLA & TCG  |  RPA & TDG  |  KDA  ; 
 ODI <=  RDI & TAH  |  RHI & TBH  |  RLI & TCH  |  RPI & TDH  |  KDI  ; 
 VDI <=  RDI & TAH  |  RHI & TBH  |  RLI & TCH  |  RPI & TDH  |  KDI  ; 
 WDA <= IDA ; 
 WDI <= IDI ; 
 WHA <= IDA ; 
 WHI <= IDI ; 
 TAA <= QED & JNA ; 
 TBA <= QED & JNB ; 
 TCA <= QED & JNC ; 
 TDA <= QED & JND ; 
 AGA <= AFA ; 
 AGI <= AFI ; 
 AGQ <= AFQ ; 
 AEA <= ADA ; 
 AEI <= ADI ; 
 AEQ <= ADQ ; 
 ACA <= ABA ; 
 ACI <= ABI ; 
 okj <= qjk ; 
 ACQ <= ABQ ; 
 AAA <= IEA & QKB |  AHA & qkb ; 
 AAI <= IEI & QKB |  AHI & qkb ; 
 AAQ <= IEQ & QKB |  AHQ & qkb ; 
 AHA <= AGA ; 
 AHI <= AGI ; 
 AHQ <= AGQ ; 
 AFA <= AEA ; 
 AFI <= AEI ; 
 AFQ <= AEQ ; 
 AIA <= IEA ; 
 ADA <= ACA ; 
 ADI <= ACI ; 
 ADQ <= ACQ ; 
 AII <= IEE ; 
 ABA <= AAA ; 
 ABI <= AAI ; 
 ABQ <= AAQ ; 
 AIQ <= IEQ ; 
 QJK <=  QJK & jqa & jpa  |  QJG  ; 
 oea <= iaa ; 
 oei <= iai ; 
 ofa <= iba ; 
 ofi <= ibi ; 
 OKB <=  QJH & jqa & qec  |  QJI  |  JPA  ; 
 QJH <=  QJH & jqa & qec  |  QJI  |  JPA  ; 
 oga <= ica ; 
 ogi <= ici ; 
 oha <= ida ; 
 ohi <= idi ; 
 QCE <= QBE ; 
 QDE <= QCE ; 
 QAE <= IGC ; 
 QBE <= QAE ; 
 QBA <= QAA ; 
 QCA <= QBA ; 
 QDI <= QCA ; 
 QPA <=  JMA & TJC  |  QCA  ; 
 qaa <=  igc  |  IGB  |  IGA  ; 
 qab <=  igc  |  IGB  |  iga  ; 
 qac <=  igc  |  igb  |  IGA  ; 
 qad <=  igc  |  igb  |  iga  ; 
 PAA <=  PAA & tja & jaa  |  JHA & TJA  |  paa & JAA  ; 
 PAC <=  PAA & tja & jaa  |  JHA & TJA  |  paa & JAA  ; 
 PAE <=  PAA & tja & jaa  |  JHA & TJA  |  paa & JAA  ; 
 PAB <=  PAA & tjb & jab  |  JHB & TJB  |  pab & JAB  ; 
 PAD <=  PAA & tjb & jab  |  JHB & TJB  |  pab & JAB  ; 
 PAF <=  PAA & tjb & jab  |  JHB & TJB  |  pab & JAB  ; 
 UEA <=  PBC & TEB  |  DAG & teb  ; 
 UFA <=  PBC & TEB  |  DAG & teb  ; 
 UEF <= QDB ; 
 UEG <= QDB ; 
 UEB <=  PBD & TEB  |  DAH & teb  ; 
 UFB <=  PBD & TEB  |  DAH & teb  ; 
 UEE <=  PFC & TEB  |  DBG & teb  ; 
 UFE <=  PFC & TEB  |  DBG & teb  ; 
 UEC <=  PFA & TEB  |  DBE & teb  ; 
 UFC <=  PFA & TEB  |  DBE & teb  ; 
 UFF <= QDB ; 
 UFG <= QDB ; 
 UED <=  PFB & TEB  |  DBF & teb  ; 
 UFD <=  PFB & TEB  |  DBF & teb  ; 
 UGA <=  PBC & TEB  |  DAK & teb  ; 
 UHA <=  PBC & TEB  |  DAK & teb  ; 
 UGF <= QDB ; 
 UGG <= QDB ; 
 UGB <=  PBD & TEB  |  DAL & teb  ; 
 UHB <=  PBD & TEB  |  DAL & teb  ; 
 UGE <=  PGC & TEB  |  DBK & teb  ; 
 UHE <=  PGC & TEB  |  DBK & teb  ; 
 UGC <=  PGA & TEB  |  DBI & teb  ; 
 UHC <=  PGA & TEB  |  DBI & teb  ; 
 UHF <= QDB ; 
 UHG <= QDB ; 
 UGD <=  PGB & TEB  |  DBJ & teb  ; 
 UHD <=  PGB & TEB  |  DBJ & teb  ; 
 qdb <= qcb ; 
 TEB <= JBC ; 
 OAB <=  RAB & TAA  |  REB & TBA  |  RIB & TCA  |  RMB & TDA  |  KAB  ; 
 VAB <=  RAB & TAA  |  REB & TBA  |  RIB & TCA  |  RMB & TDA  |  KAB  ; 
 AEC <= ADC ; 
 OAJ <=  RAJ & TAB  |  REJ & TBB  |  RIJ & TCB  |  RMJ & TDB  |  KAJ  ; 
 VAJ <=  RAJ & TAB  |  REJ & TBB  |  RIJ & TCB  |  RMJ & TDB  |  KAJ  ; 
 AFC <= AEC ; 
 WAB <= IAB ; 
 WAJ <= IAJ ; 
 WEB <= IAB ; 
 WEJ <= IAJ ; 
 OBB <=  RBB & TAC  |  RFB & TBC  |  RJB & TCC  |  RNB & TDC  |  KBB  ; 
 VBB <=  RBB & TAC  |  RFB & TBC  |  RJB & TCC  |  RNB & TDC  |  KBB  ; 
 WCJ <= TAD & ICJ ; 
 OBJ <= TAD & RBJ ; 
 VBJ <= TAD & RBJ ; 
 WBB <= IBB ; 
 WBJ <= IBJ ; 
 WFB <= IBB ; 
 WFJ <= IBJ ; 
 oec <= iac ; 
 OCB <=  RCB & TAE  |  RGB & TBE  |  RKB & TCE  |  ROB & TDE  |  KCB  ; 
 VCB <=  RCB & TAE  |  RGB & TBE  |  RKB & TCE  |  ROB & TDE  |  KCB  ; 
 QQB <=  QQB & jqb  |  QDJ  ; 
 OCJ <=  RCJ & TAF  |  RGJ & TBF  |  RKJ & TCF  |  ROJ & TDF  |  KCJ  ; 
 VCJ <=  RCJ & TAF  |  RGJ & TBF  |  RKJ & TCF  |  ROJ & TDF  |  KCJ  ; 
 WCB <= ICB ; 
 WGB <= ICB ; 
 WGJ <= ICJ ; 
 qhb <=  qab & qbb & qcb  |  jnb  ; 
 ODB <=  RDB & TAG  |  RHB & TBG  |  RLB & TCG  |  RPB & TDG  |  KDB  ; 
 VDB <=  RDB & TAG  |  RHB & TBG  |  RLB & TCG  |  RPB & TDG  |  KDB  ; 
 ODJ <=  RDJ & TAH  |  RHJ & TBH  |  RLJ & TCH  |  RPJ & TDH  |  KDJ  ; 
 VDJ <=  RDJ & TAH  |  RHJ & TBH  |  RLJ & TCH  |  RPJ & TDH  |  KDJ  ; 
 WDB <= IDB ; 
 WDJ <= IDJ ; 
 WHB <= IDB ; 
 WHJ <= IDJ ; 
 TAB <= QED & JMA ; 
 TBB <= QED & JNB ; 
 TCB <= QED & JNC ; 
 TDB <= QED & JND ; 
 AGB <= AFB ; 
 AGJ <= AFJ ; 
 AGR <= AFR ; 
 AEB <= ADB ; 
 AEJ <= ADJ ; 
 AER <= ADR ; 
 ACB <= ABB ; 
 ACJ <= ABJ ; 
 ACR <= ABR ; 
 AAB <= IEB & QKB |  AHB & qkb ; 
 AAJ <= IEJ & QKB |  AHJ & qkb ; 
 AAR <= IER & QKB |  AHR & qkb ; 
 AHB <= AGB ; 
 AHJ <= AGJ ; 
 AHR <= AGR ; 
 AFB <= AEB ; 
 AFJ <= AEJ ; 
 AFR <= AER ; 
 AIB <= IEB ; 
 ADB <= ACB ; 
 ADJ <= ACJ ; 
 ADR <= ACR ; 
 AIJ <= IEJ ; 
 ABB <= AAB ; 
 ABJ <= AAJ ; 
 ABR <= AAR ; 
 AIR <= IER ; 
 oeb <= iab ; 
 oej <= iaj ; 
 ofb <= ibb ; 
 ofj <= ibj ; 
 okk <= daa ; 
 OKC <=  QJI & jqa & qec  |  QJJ  |  JPA  ; 
 QJI <=  QJI & jqa & qec  |  QJJ  |  JPA  ; 
 ogb <= icb ; 
 ogj <= icj ; 
 ohb <= idb ; 
 ohj <= idj ; 
 okl <= daj ; 
 QBB <= QAB ; 
 QCB <= QBB ; 
 QDJ <= QCB ; 
 QPB <=  JMB & TJC  |  QCB  ; 
 okm <= dak ; 
 okn <= dal ; 
 PBA <=  PBA & tja & jba  |  JHA & TJA  |  pba & JBA  ; 
 PBC <=  PBA & tja & jba  |  JHA & TJA  |  pba & JBA  ; 
 PBE <=  PBA & tja & jba  |  JHA & TJA  |  pba & JBA  ; 
 PBB <=  PBB & tjb & jbb  |  JHB & TJB  |  pbb & JBB  ; 
 PBD <=  PBB & tjb & jbb  |  JHB & TJB  |  pbb & JBB  ; 
 PBF <=  PBB & tjb & jbb  |  JHB & TJB  |  pbb & JBB  ; 
 UIA <=  PCC & TEC  |  DAG & tec  ; 
 UJA <=  PCC & TEC  |  DAG & tec  ; 
 UIF <= QDC ; 
 UIG <= QDC ; 
 UIB <=  PCD & TEC  |  DAH & tec  ; 
 UJB <=  PCD & TEC  |  DAH & tec  ; 
 UIE <=  PFC & TEC  |  DBG & tec  ; 
 UJE <=  PFC & TEC  |  DBG & tec  ; 
 UJC <=  PFA & TEC  |  DBE & tec  ; 
 UIC <=  PFA & TEC  |  DBE & tec  ; 
 UJF <= QDC ; 
 UJG <= QDC ; 
 UID <=  PFB & TEC  |  DBF & tec  ; 
 UJD <=  PFB & TEC  |  DBF & tec  ; 
 UKA <=  PCC & TEC  |  DAK & tec  ; 
 ULA <=  PCC & TEC  |  DAK & tec  ; 
 UKF <= QDC ; 
 UKG <= QDC ; 
 UKB <=  PCD & TEC  |  DAL & tec  ; 
 ULB <=  PCD & TEC  |  DAL & tec  ; 
 UKE <=  PGC & TEC  |  DBK & tec  ; 
 ULE <=  PGC & TEC  |  DBK & tec  ; 
 UKC <=  PGA & TEC  |  DBI & tec  ; 
 ULC <=  PGA & TEC  |  DBI & tec  ; 
 ULF <= QDC ; 
 ULG <= QDC ; 
 UKD <=  PGB & TEC  |  DBJ & tec  ; 
 ULD <=  PGB & TEC  |  DBJ & tec  ; 
 QDC <= QCC ; 
 TEC <= JCC ; 
 OAC <=  RAC & TAA  |  REC & TBA  |  RIC & TCA  |  RMC & TDA  |  KAC  ; 
 VAC <=  RAC & TAA  |  REC & TBA  |  RIC & TCA  |  RMC & TDA  |  KAC  ; 
 OAK <=  RAK & TAB  |  REK & TBB  |  RIK & TCB  |  RMK & TDB  |  KAK  ; 
 VAK <=  RAK & TAB  |  REK & TBB  |  RIK & TCB  |  RMK & TDB  |  KAK  ; 
 WAC <= IAC ; 
 WAK <= IAK ; 
 WEC <= IAC ; 
 WEK <= IAK ; 
 OBC <=  RBC & TAC  |  RFC & TBC  |  RJC & TCC  |  RNC & TDC  |  KBC  ; 
 VBC <=  RBC & TAC  |  RFC & TBC  |  RJC & TCC  |  RNC & TDC  |  KBC  ; 
 OBK <=  RBK & TAD  |  RFK & TBD  |  RJK & TCD  |  RNK & TDD  |  KBK  ; 
 VBK <=  RBK & TAD  |  RFK & TBD  |  RJK & TCD  |  RNK & TDD  |  KBK  ; 
 WBC <= IBC ; 
 WBK <= IBK ; 
 WFC <= IBC ; 
 WFK <= IBK ; 
 OCC <=  RCC & TAE  |  RGC & TBE  |  RKC & TCE  |  ROC & TDE  |  KCC  ; 
 VCC <=  RCC & TAE  |  RGC & TBE  |  RKC & TCE  |  ROC & TDE  |  KCC  ; 
 QQC <=  QQC & jqb  |  QDK  ; 
 OCK <=  RCK & TAF  |  RGK & TBF  |  RKK & TCF  |  ROK & TDF  |  KCK  ; 
 VCK <=  RCK & TAF  |  RGK & TBF  |  RKK & TCF  |  ROK & TDF  |  KCK  ; 
 WCC <= ICC ; 
 WGC <= ICC ; 
 WGK <= ICK ; 
 WCK <= ICK ; 
 qhc <=  qac & qbc & qcc  |  jnc  ; 
 ODC <=  RDC & TAG  |  RHC & TBG  |  RLC & TCG  |  RPC & TDG  |  KDC  ; 
 VDC <=  RDC & TAG  |  RHC & TBG  |  RLC & TCG  |  RPC & TDG  |  KDC  ; 
 ODK <=  RDK & TAH  |  RHK & TBH  |  RLK & TCH  |  RPK & TDH  |  KDK  ; 
 VDK <=  RDK & TAH  |  RHK & TBH  |  RLK & TCH  |  RPK & TDH  |  KDK  ; 
 WDC <= IDC ; 
 WDK <= IDK ; 
 WHC <= IDC ; 
 WHK <= IDK ; 
 TAC <= QED & JNA ; 
 TBC <= QED & JNB ; 
 TCC <= QED & JMC ; 
 TDC <= QED & JND ; 
 AGC <= AFC ; 
 AGK <= AFK ; 
 AGS <= AFS ; 
 AEK <= ADK ; 
 AES <= ADS ; 
 ACC <= ABC ; 
 ACK <= ABK ; 
 ACS <= ABS ; 
 AAC <= IEC & QKB |  AHC & qkb ; 
 AAK <= IEK & QKB |  AHK & qkb ; 
 AAS <= IES & QKB |  AHS & qkb ; 
 AHC <= AGC ; 
 AHK <= AGK ; 
 AHS <= AGS ; 
 AFK <= AEK ; 
 AFS <= AES ; 
 AIC <= IEC ; 
 ADC <= ACC ; 
 ADK <= ACK ; 
 ADS <= ACS ; 
 AIK <= IEK ; 
 ABC <= AAC ; 
 ABK <= AAK ; 
 ABS <= AAS ; 
 AIS <= IES ; 
 CCA <=  BCA  |  BCB  |  BCC  |  BCD  ; 
 CAA <=  BAA  |  BAB  |  BAC  |  BAD  ; 
 oek <= iak ; 
 ofk <= ibk ; 
 ofc <= ibc ; 
 OKD <=  QJJ & jqa & qec  |  JPA  ; 
 QJJ <=  QJJ & jqa & qec  |  JPA  ; 
 ogc <= icc ; 
 ogk <= ick ; 
 ohc <= idc ; 
 QBC <= QAC ; 
 QCC <= QBC ; 
 QDK <= QCC ; 
 QPC <=  JMC & TJC  |  QCC  ; 
 oko <= dbi ; 
 okp <= dbj ; 
 okq <= dbk ; 
 PCA <=  PCA & tja & jca  |  JHA & TJA  |  pca & JCA  ; 
 PCC <=  PCA & tja & jca  |  JHA & TJA  |  pca & JCA  ; 
 PCE <=  PCA & tja & jca  |  JHA & TJA  |  pca & JCA  ; 
 PCB <=  PCB & tjb & jcb  |  JHB & TJB  |  pcb & JCB  ; 
 PCD <=  PCB & tjb & jcb  |  JHB & TJB  |  pcb & JCB  ; 
 PCF <=  PCB & tjb & jcb  |  JHB & TJB  |  pcb & JCB  ; 
 UMA <=  PDC & TED  |  DAG & ted  ; 
 UNA <=  PDC & TED  |  DAG & ted  ; 
 UMF <= QDD ; 
 UMG <= QDD ; 
 UMB <=  PDD & TED  |  DAH & ted  ; 
 UNB <=  PDD & TED  |  DAH & ted  ; 
 UME <=  PFC & TED  |  DBG & ted  ; 
 UNE <=  PFC & TED  |  DBG & ted  ; 
 UMC <=  PFA & TED  |  DBE & ted  ; 
 UNC <=  PFA & TED  |  DBE & ted  ; 
 UNF <= QDD ; 
 UNG <= QDD ; 
 UMD <=  PFB & TED  |  DBF & ted  ; 
 UND <=  PFB & TED  |  DBF & ted  ; 
 UOA <=  PDC & TED  |  DAK & ted  ; 
 UPA <=  PDC & TED  |  DAK & ted  ; 
 UOF <= QDD ; 
 UOG <= QDD ; 
 UOB <=  PDD & TED  |  DAL & ted  ; 
 UPB <=  PDD & TED  |  DAL & ted  ; 
 UOE <=  PGC & TED  |  DBK & ted  ; 
 UPE <=  PGC & TED  |  DBK & ted  ; 
 UOC <=  PGA & TED  |  DBI & ted  ; 
 UPC <=  PGA & TED  |  DBI & ted  ; 
 UPF <= QDD ; 
 UPG <= QDD ; 
 UOD <=  PGB & TED  |  DBJ & ted  ; 
 UPD <=  PGB & TED  |  DBJ & ted  ; 
 QDD <= QCD ; 
 TED <= JDC ; 
 OAD <=  RAD & TAA  |  RED & TBA  |  RID & TCA  |  RMD & TDA  |  KAD  ; 
 VAD <=  RAD & TAA  |  RED & TBA  |  RID & TCA  |  RMD & TDA  |  KAD  ; 
 OAL <=  RAL & TAB  |  REL & TBB  |  RIL & TCB  |  RML & TDB  |  KAL  ; 
 VAL <=  RAL & TAB  |  REL & TBB  |  RIL & TCB  |  RML & TDB  |  KAL  ; 
 WAD <= IAD ; 
 WAL <= IAL ; 
 WED <= IAD ; 
 WEL <= IAL ; 
 OBD <=  RBD & TAC  |  RFD & TBC  |  RJD & TCC  |  RND & TDC  |  KBD  ; 
 VBD <=  RBD & TAC  |  RFD & TBC  |  RJD & TCC  |  RND & TDC  |  KBD  ; 
 WCL <= TAD & ICL ; 
 OBL <= TAD & RBL ; 
 VBL <= TAD & RBL ; 
 WBD <= IBD ; 
 WBL <= IBL ; 
 WFD <= IBD ; 
 WFL <= IBL ; 
 OCD <=  RCD & TAE  |  RGD & TBE  |  RKD & TCE  |  ROD & TDE  |  KCD  ; 
 VCD <=  RCD & TAE  |  RGD & TBE  |  RKD & TCE  |  ROD & TDE  |  KCD  ; 
 QQD <=  QQD & jqb  |  QDL  ; 
 OCL <=  RCL & TAF  |  RGL & TBF  |  RKL & TCF  |  ROL & TDF  |  KCL  ; 
 VCL <=  RCL & TAF  |  RGL & TBF  |  RKL & TCF  |  ROL & TDF  |  KCL  ; 
 WCD <= ICD ; 
 WGD <= ICD ; 
 WGL <= ICL ; 
 qhd <=  qad & qbd & qcd  |  jnd  ; 
 ODD <=  RDD & TAG  |  RHD & TBG  |  RLD & TCG  |  RPD & TDG  |  KDD  ; 
 VDD <=  RDD & TAG  |  RHD & TBG  |  RLD & TCG  |  RPD & TDG  |  KDD  ; 
 ODL <=  RDL & TAH  |  RHL & TBH  |  RLL & TCH  |  RPL & TDH  |  KDL  ; 
 VDL <=  RDL & TAH  |  RHL & TBH  |  RLL & TCH  |  RPL & TDH  |  KDL  ; 
 WDD <= IDD ; 
 WDL <= IDL ; 
 WHD <= IDD ; 
 WHL <= IDL ; 
 TAD <= QED & JNA ; 
 TBD <= QED & JNB ; 
 TCD <= QED & JNC ; 
 TDD <= QED & JND ; 
 AGD <= AFD ; 
 AGL <= AFL ; 
 AGT <= AFT ; 
 AED <= ADD ; 
 AEL <= ADL ; 
 AET <= ADT ; 
 ACD <= ABD ; 
 ACL <= ABL ; 
 ACT <= ABT ; 
 AAD <= IED & QKB |  AHD & qkb ; 
 AAL <= IEL & QKB |  AHL & qkb ; 
 AAT <= IET & QKB |  AHT & qkb ; 
 AHD <= AGD ; 
 AHL <= AGL ; 
 AHT <= AGT ; 
 AFD <= AED ; 
 AFL <= AEL ; 
 AFT <= AET ; 
 AID <= IED ; 
 ADD <= ACD ; 
 ADT <= ACT ; 
 AIL <= IEL ; 
 ADL <= ACL ; 
 ABD <= AAD ; 
 ABL <= AAL ; 
 ABT <= AAT ; 
 AIT <= IET ; 
 CDA <=  BDA  |  BDB  |  BDC  |  BDD  ; 
 CBA <=  BBA  |  BBB  |  BBC  |  BBD  ; 
 oed <= iad ; 
 oel <= ial ; 
 ofd <= ibd ; 
 ofl <= ibl ; 
 ogd <= icd ; 
 ogl <= icl ; 
 ohd <= idd ; 
 ohl <= idl ; 
 QEB <=  QCA & JIA  |  QCB & JIB  |  QCC & JIC  |  QCD & JID  ; 
 QBD <= QAD ; 
 QCD <= QBD ; 
 QDL <= QCD ; 
 QPD <=  QCD  ; 
 okr <= pga ; 
 oks <= pgb ; 
 okt <= pgc ; 
 PDA <=  PDA & tja & jda  |  JHA & TJA  |  pda & JDA  ; 
 PDC <=  PDA & tja & jda  |  JHA & TJA  |  pda & JDA  ; 
 PDE <=  PDA & tja & jda  |  JHA & TJA  |  pda & JDA  ; 
 PDB <=  PDB & tjb & jdb  |  JHB & TJB  |  pdb & JDB  ; 
 PDD <=  PDB & tjb & jdb  |  JHB & TJB  |  pdb & JDB  ; 
 PDF <=  PDB & tjb & jdb  |  JHB & TJB  |  pdb & JDB  ; 
 UAI <=  PAE & TEE  |  DAG & tee  ; 
 UBI <=  PAE & TEE  |  DAG & tee  ; 
 UAN <= QDA ; 
 UAO <= QDA ; 
 UBN <= QDA ; 
 UBO <= QDA ; 
 UAJ <=  PAF & TEE  |  DAH & tee  ; 
 UBJ <=  PAF & TEE  |  DAH & tee  ; 
 UAM <=  PFC & TEE  |  DBG & tee  ; 
 UBM <=  PFC & TEE  |  DBG & tee  ; 
 UAK <=  PFA & TEE  |  DBE & tee  ; 
 UBK <=  PFA & TEE  |  DBE & tee  ; 
 OBP <=  RBP & TAD  |  RFP & TBD  |  RJP & TCD  |  RNP & TDD  |  KBP  ; 
 UAL <=  PFB & TEE  |  DBF & tee  ; 
 UBL <=  PFB & TEE  |  DBF & tee  ; 
 UCI <=  PAE & TEE  |  DAK & tee  ; 
 UDI <=  PAE & TEE  |  DAK & tee  ; 
 UCN <= QDA ; 
 UCO <= QDA ; 
 UCJ <=  PAF & TEE  |  DAL & tee  ; 
 UDJ <=  PAF & TEE  |  DAL & tee  ; 
 UCM <=  PGC & TEE  |  DBK & tee  ; 
 UDM <=  PGC & TEE  |  DBK & tee  ; 
 UCK <=  PGA & TEE  |  DBI & tee  ; 
 UDK <=  PGA & TEE  |  DBI & tee  ; 
 UDN <= QDA ; 
 UDO <= QDA ; 
 UCL <=  PGB & TEE  |  DBJ & tee  ; 
 UDL <=  PGB & TEE  |  DBJ & tee  ; 
 TEE <= QED & JAC ; 
 TDE <= QED & JND ; 
 OAE <=  RAE & TAA  |  REE & TBA  |  RIE & TCA  |  RME & TDA  |  KAE  ; 
 VAE <=  RAE & TAA  |  REE & TBA  |  RIE & TCA  |  RME & TDA  |  KAE  ; 
 OAM <=  RAM & TAB  |  REM & TBB  |  RIM & TCB  |  RMM & TDB  |  KAM  ; 
 VAM <=  RAM & TAB  |  REM & TBB  |  RIM & TCB  |  RMM & TDB  |  KAM  ; 
 WAE <= IAE ; 
 WAM <= IAM ; 
 WEE <= IAE ; 
 WEM <= IAM ; 
 OBE <=  RBE & TAC  |  RFE & TBC  |  RJE & TCC  |  RNE & TDC  |  KBE  ; 
 VBE <=  RBE & TAC  |  RFE & TBC  |  RJE & TCC  |  RNE & TDC  |  KBE  ; 
 KDE <=  WHE & TFD  |  VDE & TGD  ; 
 OBM <=  RBM & TAD  |  RFM & TBD  |  RJM & TCD  |  RNM & TDD  |  KBM  ; 
 VBM <=  RBM & TAD  |  RFM & TBD  |  RJM & TCD  |  RNM & TDD  |  KBM  ; 
 WBE <= IBE ; 
 WBM <= IBM ; 
 WFE <= IBE ; 
 WFM <= IBM ; 
 OCE <=  RCE & TAE  |  RGE & TBE  |  RKE & TCE  |  ROE & TDE  |  KCE  ; 
 VCE <=  RCE & TAE  |  RGE & TBE  |  RKE & TCE  |  ROE & TDE  |  KCE  ; 
 OCM <=  RCM & TAF  |  RGM & TBF  |  RKM & TCF  |  ROM & TDF  |  KCM  ; 
 VCM <=  RCM & TAF  |  RGM & TBF  |  RKM & TCF  |  ROM & TDF  |  KCM  ; 
 WCE <= ICE ; 
 WCM <= ICM ; 
 WGE <= ICE ; 
 WGM <= ICM ; 
 HIA <=  HBA & JJA  |  HDA & JJB  |  HFA & JJC  |  HHA & JJD  |  JKA  ; 
 ODE <=  RDE & TAG  |  RHE & TBG  |  RLE & TCG  |  RPE & TDG  |  KDE  ; 
 VDE <=  RDE & TAG  |  RHE & TBG  |  RLE & TCG  |  RPE & TDG  |  KDE  ; 
 ODM <=  RDM & TAH  |  RHM & TBH  |  RLM & TCH  |  RPM & TDH  |  KDM  ; 
 VDM <=  RDM & TAH  |  RHM & TBH  |  RLM & TCH  |  RPM & TDH  |  KDM  ; 
 WDE <= IDE ; 
 WDM <= IDM ; 
 WHE <= IDE ; 
 WHM <= IDM ; 
 TAE <= QED & JNA ; 
 TBE <= QED & JNB ; 
 TCE <= QED & JNC ; 
 AGE <= AFE ; 
 AGM <= AFM ; 
 AGU <= AFU ; 
 AEE <= ADE ; 
 AEM <= ADM ; 
 AEU <= ADU ; 
 ACE <= ABE ; 
 ACM <= ABM ; 
 ACU <= ABU ; 
 AAE <= IEE & QKB |  AHE & qkb ; 
 AAM <= IEM & QKB |  AHM & qkb ; 
 AAU <= IEU & QKB |  AHU & qkb ; 
 AHE <= AGE ; 
 AHM <= AGM ; 
 AHU <= AGU ; 
 AFE <= AEE ; 
 AFM <= AEM ; 
 AFU <= AEU ; 
 AIE <= IEE ; 
 ADE <= ACE ; 
 ADM <= ACM ; 
 ADU <= ACU ; 
 AIM <= IEM ; 
 ABE <= AAE ; 
 ABM <= AAM ; 
 ABU <= AAU ; 
 AIU <= IEU ; 
 CCB <=  BCE  |  BCF  |  BCG  |  BCH  ; 
 CAB <=  BAE  |  BAF  |  BAG  |  BAH  ; 
 oee <= iae ; 
 oem <= iam ; 
 ofe <= ibe ; 
 ofm <= ibm ; 
 EAA <=  DAA & qlb & jea  |  daa & JEA  |  EAA & QLB  ; 
 EAB <=  DAB & qlb & jeb  |  dab & JEB  |  EAB & QLB  ; 
 oge <= ice ; 
 ogm <= icm ; 
 ohe <= ide ; 
 ohm <= idm ; 
 EAC <=  DAC & qlb & jec  |  dac & JEC  |  EAC & QLB  ; 
 EAD <=  DAD & qlb & jed  |  dad & JED  |  EAD & QLB  ; 
 DAA <=  DAA & qlc & qld  |  IFA & QLC  |  EAA & QLD  ; 
 DAE <=  DAA & qlc & qld  |  IFA & QLC  |  EAA & QLD  ; 
 DAI <=  DAA & qlc & qld  |  IFA & QLC  |  EAA & QLD  ; 
 DAB <=  DAB & qlc & qld  |  IFB & QLC  |  EAB & QLD  ; 
 DAF <=  DAB & qlc & qld  |  IFB & QLC  |  EAB & QLD  ; 
 DAJ <=  DAB & qlc & qld  |  IFB & QLC  |  EAB & QLD  ; 
 DAC <=  DAC & qlc & qld  |  IFC & QLC  |  EAC & QLD  ; 
 DAG <=  DAC & qlc & qld  |  IFC & QLC  |  EAC & QLD  ; 
 DAK <=  DAC & qlc & qld  |  IFC & QLC  |  EAC & QLD  ; 
 DAD <=  DAD & qlc & qld  |  IFD & QLC  |  EAD & QLD  ; 
 DAH <=  DAD & qlc & qld  |  IFD & QLC  |  EAD & QLD  ; 
 DAL <=  DAD & qlc & qld  |  IFD & QLC  |  EAD & QLD  ; 
 UEI <=  PBE & TEF  |  DAG & tef  ; 
 UFI <=  PBE & TEF  |  DAG & tef  ; 
 UEN <= QDB ; 
 UEO <= QDB ; 
 UEJ <=  PBF & TEF  |  DAH & tef  ; 
 UFJ <=  PBF & TEF  |  DAH & tef  ; 
 UEM <=  PFC & TEF  |  DBG & tef  ; 
 UFM <=  PFC & TEF  |  DBG & tef  ; 
 UFK <=  PFA & TEF  |  DBE & tef  ; 
 UEK <=  PFA & TEF  |  DBE & tef  ; 
 UFN <= QDB ; 
 UFO <= QDB ; 
 UEL <=  PFB & TEF  |  DBF & tef  ; 
 UFL <=  PFB & TEF  |  DBF & tef  ; 
 UGI <=  PBE & TEF  |  DAK & tef  ; 
 UHI <=  PBE & TEF  |  DAK & tef  ; 
 UGN <= QDB ; 
 UGO <= QDB ; 
 UGJ <=  PBF & TEF  |  DAL & tef  ; 
 UHJ <=  PBF & TEF  |  DAL & tef  ; 
 UGM <=  PGC & TEF  |  DBK & tef  ; 
 UHM <=  PGC & TEF  |  DBK & tef  ; 
 UGK <=  PGA & TEF  |  DBI & tef  ; 
 UHK <=  PGA & TEF  |  DBI & tef  ; 
 UHN <= QDB ; 
 UHO <= QDB ; 
 UGL <=  PGB & TEF  |  DBJ & tef  ; 
 UHL <=  PGB & TEF  |  DBJ & tef  ; 
 TEF <= JBC ; 
 OAF <=  RAF & TAA  |  REFF  & TBA  |  RIF & TCA  |  RMF & TDA  |  KAF  ; 
 VAF <=  RAF & TAA  |  REFF  & TBA  |  RIF & TCA  |  RMF & TDA  |  KAF  ; 
 TFA <=  QEB  ; 
 tga <=  QEB  |  QEC  ; 
 OAN <=  RAN & TAB  |  REN & TBB  |  RIN & TCB  |  RMN & TDB  |  KAN  ; 
 VAN <=  RAN & TAB  |  REN & TBB  |  RIN & TCB  |  RMN & TDB  |  KAN  ; 
 WAF <= IAF ; 
 WAN <= IAN ; 
 WEF <= IAF ; 
 WEN <= IAN ; 
 OBF <=  RBF & TAC  |  RFF & TBC  |  RJF & TCC  |  RNF & TDC  |  KBF  ; 
 VBF <=  RBF & TAC  |  RFF & TBC  |  RJF & TCC  |  RNF & TDC  |  KBF  ; 
 TFB <=  QEB  ; 
 tgb <=  QEB  |  QEC  ; 
 OBN <=  RBN & TAD  |  RFN & TBD  |  RJN & TCD  |  RNN & TDD  |  KBN  ; 
 VBN <=  RBN & TAD  |  RFN & TBD  |  RJN & TCD  |  RNN & TDD  |  KBN  ; 
 WBF <= IBF ; 
 WBN <= IBN ; 
 WFF <= IBF ; 
 WFN <= IBN ; 
 OCF <=  RCF & TAE  |  RGF & TBE  |  RKF & TCE  |  ROF & TDE  |  KCF  ; 
 VCF <=  RCF & TAE  |  RGF & TBE  |  RKF & TCE  |  ROF & TDE  |  KCF  ; 
 TFC <=  QEB  ; 
 tgc <=  QEB  |  QEC  ; 
 OCN <=  RCN & TAF  |  RGN & TBF  |  RKN & TCF  |  RON & TDF  |  KCN  ; 
 VCN <=  RCN & TAF  |  RGN & TBF  |  RKN & TCF  |  RON & TDF  |  KCN  ; 
 WCF <= ICF ; 
 WCN <= ICN ; 
 WGF <= ICF ; 
 WGN <= ICN ; 
 HIB <=  HBB & JJA  |  HDB & JJB  |  HFB & JJC  |  HHB & JJD  |  JKB  ; 
 ODF <=  RDF & TAG  |  RHF & TBG  |  RLF & TCG  |  RPF & TDG  |  KDF  ; 
 VDF <=  RDF & TAG  |  RHF & TBG  |  RLF & TCG  |  RPF & TDG  |  KDF  ; 
 TFD <=  QEB  ; 
 tgd <=  QEB  |  QEC  ; 
 ODN <=  RDN & TAH  |  RHN & TBH  |  RLN & TCH  |  RPN & TDH  |  KDN  ; 
 VDN <=  RDN & TAH  |  RHN & TBH  |  RLN & TCH  |  RPN & TDH  |  KDN  ; 
 WDF <= IDF ; 
 WDN <= IDN ; 
 WHF <= IDF ; 
 WHN <= IDN ; 
 TAF <= QED & JNA ; 
 TBF <= QED & JNB ; 
 TCF <= QED & JNC ; 
 TDF <= QED & JND ; 
 AGF <= AFF ; 
 AGN <= AFN ; 
 AGV <= AFV ; 
 AEF <= ADF ; 
 AEN <= ADN ; 
 AEV <= ADV ; 
 oki <= qje ; 
 ACF <= ABF ; 
 ACN <= ABM ; 
 ACV <= ABV ; 
 AAF <= IEF & QKB |  AHF & qkb ; 
 AAN <= IEN & QKB |  AHN & qkb ; 
 AAV <= IEV & QKB |  AHV & qkb ; 
 AHF <= AGF ; 
 AHN <= AGN ; 
 AHV <= AGV ; 
 AFF <= AEF ; 
 AFN <= AEN ; 
 AFV <= AEV ; 
 AIF <= IEF ; 
 ADF <= ACF ; 
 ADN <= ACN ; 
 ADV <= ACV ; 
 AIN <= IEN ; 
 ABF <= AAF ; 
 ABN <= AAN ; 
 ABV <= AAV ; 
 AIV <= IEV ; 
 ebc <=  dbc & qlb & qle  |  ebc & QLB  |  pfc & QLE  ; 
 QJP <=  QJP & qlf  |  IJE  ; 
 CDB <=  BDE  |  BDF  |  BDG  |  BDH  ; 
 CBB <=  BBE  |  BBF  |  BBG  |  BBH  ; 
 oef <= iaf ; 
 oen <= ian ; 
 off <= ibf ; 
 ofn <= ibn ; 
 OKH <=  QJD & ijd & ije  |  JEE & JPF  ; 
 QJD <=  QJD & ijd & ije  |  JEE & JPF  ; 
 qec <=  QJE & JFB & qjh  |  ijd & jpc  |  jpb  ; 
 qed <=  QJE & JFB & qjh  |  ijd & jpc  |  jpb  ; 
 QJF <=  QJF & jpe  |  IHB  |  IJD  |  QJG  ; 
 ogf <= icf ; 
 ogn <= icn ; 
 ohf <= idf ; 
 ohn <= idn ; 
 OKA <=  QJM & qeb  |  IJE & qjd  ; 
 QJM <=  QJM & qeb  |  IJE & qjd  ; 
 QJN <=  QJM & qeb  |  IJE & qjd  ; 
 OKE <=  QJC & jfa  |  IJE  ; 
 QJC <=  QJC & jfa  |  IJE  ; 
 QJE <=  QJE & jle  |  IJE  ; 
 QJG <=  IJE & jle  ; 
 eba <=  dba & qlb & qle  |  eba & QLB  |  pfa & QLE  ; 
 ebb <=  dbb & qlb & qle  |  ebb & QLB  |  pfb & QLE  ; 
 qla <=  qja  |  qjb  |  IJD  ; 
 qlb <=  qja  |  qla  |  IJD  ; 
 DBA <=  DBA & qlc & qlf  |  HIA & QLC  |  EBA & QLF  ; 
 DBE <=  DBA & qlc & qlf  |  HIA & QLC  |  EBA & QLF  ; 
 DBI <=  DBA & qlc & qlf  |  HIA & QLC  |  EBA & QLF  ; 
 DBB <=  DBB & qlc & qlf  |  HIB & QLC  |  EBB & QLF  ; 
 DBF <=  DBB & qlc & qlf  |  HIB & QLC  |  EBB & QLF  ; 
 DBJ <=  DBB & qlc & qlf  |  HIB & QLC  |  EBB & QLF  ; 
 DBC <=  DBC & qlc & qlf  |  HIC & QLC  |  EBC & QLF  ; 
 DBG <=  DBC & qlc & qlf  |  HIC & QLC  |  EBC & QLF  ; 
 DBK <=  DBC & qlc & qlf  |  HIC & QLC  |  EBC & QLF  ; 
 qlc <=  qja  |  qfa  ; 
 qle <=  tjc  ; 
 UII <=  PCE & TEG  |  DAG & teg  ; 
 UJI <=  PCE & TEG  |  DAG & teg  ; 
 UIN <= QDC ; 
 UIO <= QDC ; 
 UIJ <=  PCF & TEG  |  DAH & teg  ; 
 UJJ <=  PCF & TEG  |  DAH & teg  ; 
 UIM <=  PFC & TEG  |  DBG & teg  ; 
 UJM <=  PFC & TEG  |  DBG & teg  ; 
 UIK <=  PFA & TEG  |  DBE & teg  ; 
 UJK <=  PFA & TEG  |  DBE & teg  ; 
 UJN <= QDC ; 
 UJO <= QDC ; 
 UIL <=  PFB & TEG  |  DBF & teg  ; 
 UJL <=  PFB & TEG  |  DBF & teg  ; 
 UKI <=  PCE & TEG  |  DAK & teg  ; 
 ULI <=  PCE & TEG  |  DAK & teg  ; 
 UKN <= QDC ; 
 UKO <= QDC ; 
 UKJ <=  PCF & TEG  |  DAL & teg  ; 
 ULJ <=  PCF & TEG  |  DAL & teg  ; 
 UKM <=  PGC & TEG  |  DBK & teg  ; 
 ULM <=  PGC & TEG  |  DBK & teg  ; 
 UKK <=  PGA & TEG  |  DBI & teg  ; 
 ULK <=  PGA & TEG  |  DBI & teg  ; 
 ULN <= QDC ; 
 ULO <= QDC ; 
 UKL <=  PGB & TEG  |  DBJ & teg  ; 
 ULL <=  PGB & TEG  |  DBJ & teg  ; 
 TEG <= JCC ; 
 OAG <=  RAG & TAA  |  REG & TBA  |  RIG & TCA  |  RMG & TDA  |  KAG  ; 
 VAG <=  RAG & TAA  |  REG & TBA  |  RIG & TCA  |  RMG & TDA  |  KAG  ; 
 FAA <=  FAA & tjd & jla  |  JLA & faa  ; 
 OAO <=  RAO & TAB  |  REO & TBB  |  RIO & TCB  |  RMO & TDB  |  KAO  ; 
 VAO <=  RAO & TAB  |  REO & TBB  |  RIO & TCB  |  RMO & TDB  |  KAO  ; 
 WAG <= IAG ; 
 WAO <= IAO ; 
 WEG <= IAG ; 
 WEO <= IAO ; 
 FAB <=  FAB & tjd & jlb  |  JLB & fab  ; 
 OBG <=  RBG & TAC  |  RFG & TBC  |  RJG & TCC  |  RNG & TDC  |  KBG  ; 
 VBG <=  RBG & TAC  |  RFG & TBC  |  RJG & TCC  |  RNG & TDC  |  KBG  ; 
 FAC <=  FAC & tjd & jlc  |  JLC & fac  ; 
 OBO <=  RBO & TAD  |  RFO & TBD  |  RJO & TCD  |  RNO & TDD  |  KBO  ; 
 VBO <=  RBO & TAD  |  RFO & TBD  |  RJO & TCD  |  RNO & TDD  |  KBO  ; 
 WBG <= IBG ; 
 WBO <= IBO ; 
 WFG <= IBG ; 
 WFO <= IBO ; 
 FAD <=  FAD & tjd & jld  |  JLD & fad  ; 
 OCG <=  RCG & TAE  |  RGG & TBE  |  RKG & TCE  |  ROG & TDE  |  KCG  ; 
 VCG <=  RCG & TAE  |  RGG & TBE  |  RKG & TCE  |  ROG & TDE  |  KCG  ; 
 ohk <= idk ; 
 OCO <=  RCO & TAF  |  RGO & TBF  |  RKO & TCF  |  ROO & TDF  |  KCO  ; 
 VCO <=  RCO & TAF  |  RGO & TBF  |  RKO & TCF  |  ROO & TDF  |  KCO  ; 
 WCG <= ICG ; 
 WCO <= ICO ; 
 WGG <= ICG ; 
 WGO <= ICO ; 
 HIC <=  HBC & JJA  |  HDC & JJB  |  HFC & JJC  |  HHC & JJD  |  JKC  ; 
 ODG <=  RDG & TAG  |  RHG & TBG  |  RLG & TCG  |  RPG & TDG  |  KDG  ; 
 VDG <=  RDG & TAG  |  RHG & TBG  |  RLG & TCG  |  RPG & TDG  |  KDG  ; 
 QPE <= JLE ; 
 ODO <=  RDO & TAH  |  RHO & TBH  |  RLO & TCH  |  RPO & TDH  |  KDO  ; 
 VDO <=  RDO & TAH  |  RHO & TBH  |  RLO & TCH  |  RPO & TDH  |  KDO  ; 
 WDG <= IDG ; 
 WDO <= IDO ; 
 WHG <= IDG ; 
 WHO <= IDO ; 
 TAG <= QED & JNA ; 
 TBG <= QED & JNB ; 
 TCG <= QED & JNC ; 
 TDG <= QED & JND ; 
 AGG <= AFG ; 
 AGO <= AFO ; 
 AGW <= AFW ; 
 AEG <= ADG ; 
 AEO <= ADO ; 
 AEW <= ADW ; 
 ACG <= ABG ; 
 ACO <= ABO ; 
 ACW <= ABW ; 
 AAG <= IEG & QKB |  AHG & qkb ; 
 AAO <= IEO & QKB |  AHO & qkb ; 
 AAW <= IEW & QKB |  AHV & qkb ; 
 AHG <= AGG ; 
 AHO <= AGO ; 
 AHW <= AGW ; 
 AFG <= AEG ; 
 AFO <= AEO ; 
 AFW <= AEW ; 
 AIG <= IEG ; 
 ADG <= ACG ; 
 ADO <= ACO ; 
 ADW <= ACW ; 
 AIO <= IEO ; 
 ABG <= AAG ; 
 ABO <= AAO ; 
 ABW <= AAW ; 
 AIW <= IEW ; 
 oeg <= iag ; 
 oeo <= iao ; 
 ofg <= ibg ; 
 ofo <= ibo ; 
 ogg <= icg ; 
 ogo <= ico ; 
 ohg <= idg ; 
 oho <= ido ; 
 okf <= jfb ; 
 OKG <= JPC ; 
 QJA <= IJB ; 
 QJB <= QJA ; 
 OJA <= JPE ; 
 OJB <= JOA ; 
 ojd <= jle ; 
 oje <= jfb ; 
 QLG <= IJF ; 
 QLH <= QLG ; 
 PEA <=  PEA & tma & jga  |  JGA & pea  ; 
 PFA <=  PEA & tma & jga  |  JGA & pea  ; 
 PGA <=  PEA & tma & jga  |  JGA & pea  ; 
 PEB <=  PEB & tma & jgb  |  JGB & peb  ; 
 PFB <=  PEB & tma & jgb  |  JGB & peb  ; 
 PGB <=  PEB & tma & jgb  |  JGB & peb  ; 
 PEC <=  PEC & tma & jgc  |  JGC & pec  ; 
 PFC <=  PEC & tma & jgc  |  JGC & pec  ; 
 PGC <=  PEC & tma & jgc  |  JGC & pec  ; 
 QLD <=  QPE  |  IJF  ; 
 QLF <=  IJF  |  QLE  ; 
 UMI <=  PDE & TEH  |  DAG & teh  ; 
 UNI <=  PDE & TEH  |  DAG & teh  ; 
 UMN <= QDD ; 
 UMO <= QDD ; 
 UMJ <=  PDF & TEH  |  DAH & teh  ; 
 UNJ <=  PDF & TEH  |  DAH & teh  ; 
 UMM <=  PFC & TEH  |  DBG & teh  ; 
 UNM <=  PFC & TEH  |  DBG & teh  ; 
 UMK <=  PFA & TEH  |  DBE & teh  ; 
 UNK <=  PFA & TEH  |  DBE & teh  ; 
 UNN <= QDD ; 
 UNO <= QDD ; 
 UML <=  PFB & TEH  |  DBF & teh  ; 
 UNL <=  PFB & TEH  |  DBF & teh  ; 
 GAB <=  GAB & gaa  |  TMA  |  gab & GAA  ; 
 UOI <=  PDE & TEH  |  DAK & teh  ; 
 UPI <=  PDE & TEH  |  DAK & teh  ; 
 UON <= QDD ; 
 UOO <= QDD ; 
 UOJ <=  PDF & TEH  |  DAL & teh  ; 
 UPJ <=  PDF & TEH  |  DAL & teh  ; 
 UOM <=  PGC & TEH  |  DBK & teh  ; 
 UPM <=  PGC & TEH  |  DBK & teh  ; 
 UOK <=  PGA & TEH  |  DBI & teh  ; 
 UPK <=  PGA & TEH  |  DBI & teh  ; 
 UPN <= QDD ; 
 UPO <= QDD ; 
 UOL <=  PGB & TEH  |  DBJ & teh  ; 
 UPL <=  PGB & TEH  |  DBJ & teh  ; 
 TEH <= JDC ; 
 OAH <=  RAH & TAA  |  REH & TBA  |  RIH & TCA  |  RMH & TDA  |  KAH  ; 
 VAH <=  RAH & TAA  |  REH & TBA  |  RIH & TCA  |  RMH & TDA  |  KAH  ; 
 OAP <=  RAP & TAB  |  REP & TBB  |  RIP & TCB  |  RMP & TDB  |  KAP  ; 
 VAP <=  RAP & TAB  |  REP & TBB  |  RIP & TCB  |  RMP & TDB  |  KAP  ; 
 WAH <= IAH ; 
 WAP <= IAP ; 
 WEH <= IAH ; 
 WEP <= IAP ; 
 GAA <=  gaa  |  TMA  ; 
 OBH <=  RBH & TAC  |  RFH & TBC  |  RJH & TCC  |  RNH & TDC  |  KBH  ; 
 VBH <=  RBH & TAC  |  RFH & TBC  |  RJH & TCC  |  RNH & TDC  |  KBH  ; 
 VBP <=  RBP & TAD  |  RFP & TBD  |  RJP & TCD  |  RNP & TDD  |  KBP  ; 
 WCH <= ICH ; 
 WBH <= IBH ; 
 WBP <= IBP ; 
 WFH <= IBH ; 
 WFP <= IBP ; 
 OCH <=  RCH & TAE  |  RGH & TBE  |  RKH & TCE  |  ROH & TDE  |  KCH  ; 
 VCH <=  RCH & TAE  |  RGH & TBE  |  RKH & TCE  |  ROH & TDE  |  KCH  ; 
 OCP <=  RCP & TAF  |  RGP & TBF  |  RKP & TCF  |  ROP & TDF  |  KCP  ; 
 VCP <=  RCP & TAF  |  RGP & TBF  |  RKP & TCF  |  ROP & TDF  |  KCP  ; 
 WGH <= ICH ; 
 WGP <= ICP ; 
 WCP <= ICP ; 
 HID <=  JJA  |  JJB  |  JJC  |  JJD  |  JKD  ; 
 OJC <=  JJA  |  JJB  |  JJC  |  JJD  |  JKD  ; 
 ODH <=  RDH & TAG  |  RHH & TBG  |  RLH & TCG  |  RPH & TDG  |  KDH  ; 
 VDH <=  RDH & TAG  |  RHH & TBG  |  RLH & TCG  |  RPH & TDG  |  KDH  ; 
 GAC <=  GAC & jra  |  gac & JRA  |  TMA  ; 
 TJA <= QKA ; 
 TJB <= QKA ; 
 TJC <= QKA ; 
 TJD <= QKA ; 
 ODP <=  RDP & TAH  |  RHP & TBH  |  RLP & TCH  |  RPP & TDH  |  KDP  ; 
 VDP <=  RDP & TAH  |  RHP & TBH  |  RLP & TCH  |  RPP & TDH  |  KDP  ; 
 WDH <= IDH ; 
 WDP <= IDP ; 
 WHH <= IDH ; 
 WHP <= IDP ; 
 TAH <= QED & JNA ; 
 TBH <= QED & JNB ; 
 TCH <= QED & JNC ; 
 TDH <= QED & JND ; 
 AGH <= AFH ; 
 AGP <= AFP ; 
 AGX <= AFX ; 
 AEH <= ADH ; 
 AEP <= ADP ; 
 AEX <= ADX ; 
 oku <= faa ; 
 ACH <= ABH ; 
 ACP <= ABP ; 
 ACX <= ABX ; 
 okv <= fab ; 
 AAH <= IEH & QKB |  AHH & qkb ; 
 AAP <= IEP & QKB |  AHP & qkb ; 
 AAX <= IEX & QKB |  AHX & qkb ; 
 AHH <= AGH ; 
 AHP <= AGP ; 
 AHX <= AGX ; 
 AFH <= AEH ; 
 AFP <= AEP ; 
 AFX <= AEX ; 
 AIH <= IEH ; 
 ADH <= ACH ; 
 ADP <= ACP ; 
 ADX <= ACX ; 
 AIP <= IEP ; 
 ABH <= AAH ; 
 ABP <= AAP ; 
 ABX <= AAX ; 
 AIX <= IEX ; 
 HAA <= GAA ; 
 HBA <= HAA ; 
 HCA <= HBA ; 
 HDA <= HCA ; 
 HAB <= GAB ; 
 HBB <= HAB ; 
 HCB <= HBB ; 
 HDB <= HCB ; 
 HAC <= GAC ; 
 HBC <= HAC ; 
 HCC <= HBC ; 
 HDC <= HCC ; 
 oeh <= iah ; 
 oep <= iap ; 
 ofh <= ibh ; 
 ofp <= ibp ; 
 HEA <= HDA ; 
 HFA <= HEA ; 
 HGA <= HFA ; 
 HHA <= HGA ; 
 HEB <= HDB ; 
 HFB <= HEB ; 
 HGB <= HFB ; 
 HHB <= HGB ; 
 HEC <= HDC ; 
 HFC <= HEC ; 
 HGC <= HFC ; 
 HHC <= HGC ; 
 ogh <= ich ; 
 ogp <= icp ; 
 ohh <= idh ; 
 ohp <= idp ; 
 QFA <= TJA ; 
 TMA <= IHA ; 
 QKB <=  QKA  |  TMA  ; 
 okw <= fac ; 
 okx <= fad ; 
 QKA <=  QJC & JFA  ; 
end
ram_16x4 rinst_0({&RAA,&RAB,&RAC,&RAD},{WAA,WAB,WAC,VAD},{uaa,uab,uac,uad}, uae, UAF, IZZ); 
ram_16x4 rinst_1({&RAA,&RAB,&RAC,&RAD},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_2({&RAI,&RAJ,&RAK,&RAL},{WAI,WAJ,WAK,WAL},{uaa,uab,uac,uad}, uae, UAG, IZZ); 
ram_16x4 rinst_3({&RAI,&RAJ,&RAK,&RAL},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_4({&RDA,&RDB,&RDC,&RDD},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_5({&RBA,&RBB,&RBC,&RBD},{WBA,WBB,WBC,WBD},{uba,ubb,ubc,ubd}, ube, UBF, IZZ); 
ram_16x4 rinst_6({&RBA,&RBB,&RBC,&RBD},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_7({&RBI,&RBJ,&RBK,&RBL},{WBI,WBJ,WBK,WBL},{uba,ubb,ubc,ubd}, ube, UBG, IZZ); 
ram_16x4 rinst_8({&RBI,&RBJ,&RBK,&RBL},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_9({&RCA,&RCB,&RCC,&RCD},{WCA,WCB,WCC,WCD},{uca,ucb,ucc,ucd}, uce, UCF, IZZ); 
ram_16x4 rinst_10({&RCA,&RCB,&RCC,&RCD},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_11({&RCI,&RCJ,&RCK,&RCL},{WCI,WCJ,WCK,WCL},{uca,ucb,ucc,ucd}, uce, UCG, IZZ); 
ram_16x4 rinst_12({&RCI,&RCJ,&RCK,&RCL},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_13({&RDA,&RDB,&RDC,&RDD},{WDA,WDB,WDC,WDD},{uda,udb,udc,udd}, ude, UDF, IZZ); 
ram_16x4 rinst_14({&RDI,&RDJ,&RDK,&RDL},{WDI,WDJ,WDK,WDL},{uda,udb,udc,udd}, ude, UDG, IZZ); 
ram_16x4 rinst_15({&RDI,&RDJ,&RDK,&RDL},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_16({&REA,&REB,&REC,&RED},{WAA,WAB,WAC,WAD},{uea,ueb,uec,ued}, uee, UEF, IZZ); 
ram_16x4 rinst_17({&REA,&REB,&REC,&RED},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_18({&REI,&REJ,&REK,&REL},{WAI,WAJ,WAK,WAL},{uea,ueb,uec,ued}, uee, UEG, IZZ); 
ram_16x4 rinst_19({&REI,&REJ,&REK,&REL},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_20({&RFA,&RFB,&RFC,&RFD},{WBA,WBB,WBC,WBD},{ufa,ufb,ufc,ufd}, ufe, UFF, IZZ); 
ram_16x4 rinst_21({&RFA,&RFB,&RFC,&RFD},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_22({&RFI,&RFJ,&RFK,&RFL},{WBI,WBJ,WBK,WBL},{ufa,ufb,ufc,ufd}, ufe, UFG, IZZ); 
ram_16x4 rinst_23({&RFI,&RFJ,&RFK,&RFL},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_24({&RGA,&RGB,&RGC,&RGD},{WCA,WCB,WCC,VCD},{uga,ugb,ugc,ugd}, uge, UGF, IZZ); 
ram_16x4 rinst_25({&RGA,&RGB,&RGC,&RGD},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_26({&RGI,&RGJ,&RGK,&RGL},{WCI,WCJ,WCK,WCL},{uga,ugb,ugc,ugd}, uge, UGG, IZZ); 
ram_16x4 rinst_27({&RGI,&RGJ,&RGK,&RGL},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_28({&RHA,&RHB,&RHC,&RHD},{WDA,WDB,WDC,WDD},{uha,uhb,uhc,uhd}, uhe, UHF, IZZ); 
ram_16x4 rinst_29({&RHA,&RHB,&RHC,&RHD},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_30({&RHI,&RHJ,&RHK,&RHL},{WDI,WDJ,WDK,WDL},{uha,uhb,uhc,uhd}, uhe, UHG, IZZ); 
ram_16x4 rinst_31({&RHI,&RHJ,&RHK,&RHL},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_32({&RIA,&RIB,&RIC,&RID},{WAA,WAB,WAC,WAD},{uia,uib,uic,uid}, uie, UIF, IZZ); 
ram_16x4 rinst_33({&RIA,&RIB,&RIC,&RID},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_34({&RII,&RIJ,&RIK,&RIL},{WAI,WAJ,WAK,WAL},{uia,uib,uic,uid}, uie, UIG, IZZ); 
ram_16x4 rinst_35({&RII,&RIJ,&RIK,&RIL},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_36({&RJA,&RJB,&RJC,&RJD},{WBA,WBB,WBC,WBD},{uja,ujb,ujc,ufd}, uje, UJF, IZZ); 
ram_16x4 rinst_37({&RJA,&RJB,&RJC,&RJD},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_38({&RJI,&RJJ,&RJK,&RJL},{WBI,WBJ,WBK,WBL},{uja,ujb,ujc,ujd}, uje, UJG, IZZ); 
ram_16x4 rinst_39({&RJI,&RJJ,&RJK,&RJL},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_40({&RKA,&RKB,&RKC,&RKD},{WCA,WCB,WCC,VCD},{uka,ukb,ukc,ukd}, uke, UKF, IZZ); 
ram_16x4 rinst_41({&RKA,&RKB,&RKC,&RKD},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_42({&RKI,&RKJ,&RKK,&RKL},{WCI,WCJ,WCK,WCL},{uka,ukb,ukc,ukd}, uke, UKG, IZZ); 
ram_16x4 rinst_43({&RKI,&RKJ,&RKK,&RKL},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_44({&RLA,&RLB,&RLC,&RLD},{WDA,WDB,WDC,WDD},{ula,ulb,ulc,uld}, ule, ULF, IZZ); 
ram_16x4 rinst_45({&RLA,&RLB,&RLC,&RLD},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_46({&RLI,&RLJ,&RLK,&RLL},{WDI,WDJ,WDK,WDL},{ula,ulb,ulc,uld}, ule, ULG, IZZ); 
ram_16x4 rinst_47({&RLI,&RLJ,&RLK,&RLL},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_48({&RMA,&RMB,&RMC,&RMD},{WAA,WAB,WAC,WAD},{uma,umb,umc,umd}, ume, UMF, IZZ); 
ram_16x4 rinst_49({&RMA,&RMB,&RMC,&RMD},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_50({&RMI,&RMJ,&RMK,&RML},{WAI,WAJ,WAK,WAL},{uma,umb,umc,umd}, ume, UMG, IZZ); 
ram_16x4 rinst_51({&RMI,&RMJ,&RMK,&RML},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_52({&RNA,&RNB,&RNC,&RND},{WBA,WBB,WBC,WBD},{una,unb,unc,ufd}, une, UNF, IZZ); 
ram_16x4 rinst_53({&RNA,&RNB,&RNC,&RND},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_54({&RNI,&RNJ,&RNK,&RNL},{WBI,WBJ,WBK,WBL},{una,unb,unc,und}, une, UNG, IZZ); 
ram_16x4 rinst_55({&RNI,&RNJ,&RNK,&RNL},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_56({&ROA,&ROB,&ROC,&ROD},{WCA,WCB,WCC,VCD},{uoa,uob,uoc,uod}, uoe, UOF, IZZ); 
ram_16x4 rinst_57({&ROA,&ROB,&ROC,&ROD},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_58({&ROI,&ROJ,&ROK,&ROL},{WCI,WCJ,WCK,WCL},{uoa,uob,uoc,uod}, uoe, UOG, IZZ); 
ram_16x4 rinst_59({&ROI,&ROJ,&ROK,&ROL},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_60({&RPA,&RPB,&RPC,&RPD},{WDA,WDB,WDC,WDD},{upa,upb,upc,upd}, upe, UPF, IZZ); 
ram_16x4 rinst_61({&RPA,&RPB,&RPC,&RPD},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_62({&RPI,&RPJ,&RPK,&RPL},{WDI,WDJ,WDK,WDL},{upa,upb,upc,upd}, upe, UPG, IZZ); 
ram_16x4 rinst_63({&RPI,&RPJ,&RPK,&RPL},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_64({&RAE,&RAF,&RAG,&RAH},{WAE,WAF,WAG,WAH},{uai,uaj,uak,ual}, uam, UAN, IZZ); 
ram_16x4 rinst_65({&RAE,&RAF,&RAG,&RAH},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_66({&RAM,&RAN,&RAO,&RAP},{WAM,WAN,WAO,WAP},{uai,uaj,uak,ual}, uam, UAO, IZZ); 
ram_16x4 rinst_67({&RAM,&RAN,&RAO,&RAP},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_68({&RDE,&RDF,&RDG,&RDH},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_69({&RBE,&RBF,&RBG,&RBH},{WBE,WBF,WBG,WBH},{ubi,ubj,ubk,ubl}, ubm, UBN, IZZ); 
ram_16x4 rinst_70({&RBE,&RBF,&RBG,&RBH},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_71({&RBM,&RBN,&RBO,&RBP},{WBM,WBN,WBO,WBP},{ubi,ubj,ubk,ubl}, ubm, UBO, IZZ); 
ram_16x4 rinst_72({&RBM,&RBN,&RBO,&RBP},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_73({&RCE,&RCF,&RCG,&RCH},{WCE,WCF,WCG,WCH},{uci,ucj,uck,ucl}, ucm, UCN, IZZ); 
ram_16x4 rinst_74({&RCE,&RCF,&RCG,&RCH},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_75({&RCM,&RCN,&RCO,&RCP},{WCM,WCN,WCO,WCP},{uci,ucj,uck,ucl}, ucm, UCO, IZZ); 
ram_16x4 rinst_76({&RCM,&RCN,&RCO,&RCP},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_77({&RDE,&RDF,&RDG,&RDH},{WDE,WDF,WDG,WDH},{udi,udj,udk,udl}, udm, UDN, IZZ); 
ram_16x4 rinst_78({&RDM,&RDN,&RDO,&RDP},{WDM,WDN,WDO,WDP},{udi,udj,udk,udl}, udm, UDO, IZZ); 
ram_16x4 rinst_79({&RDM,&RDN,&RDO,&RDP},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_80({&REE,&REFF ,&REG,&REH},{WAE,WAF,WAG,WAH},{uei,uei,uek,uel}, uem, UEN, IZZ); 
ram_16x4 rinst_81({&REE,&REFF ,&REG,&REH},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_82({&REM,&REN,&REO,&REP},{WAM,WAN,WAO,WAP},{uei,uej,uek,uel}, uem, UEO, IZZ); 
ram_16x4 rinst_83({&REM,&REN,&REO,&REP},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_84({&RFE,&RFF,&RFG,&RFH},{WBE,WBF,WBG,WBH},{ufi,ufj,ufk,ufl}, ufm, UFN, IZZ); 
ram_16x4 rinst_85({&RFE,&RFF,&RFG,&RFH},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_86({&RFM,&RFN,&RFO,&RFP},{WBM,WBN,WBO,WBP},{ufi,ufj,ufk,ufl}, ufm, UFO, IZZ); 
ram_16x4 rinst_87({&RFM,&RFN,&RFO,&RFP},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_88({&RGE,&RGF,&RGG,&RGH},{WCE,WCF,WCG,WCH},{ugi,ugj,ugk,ugl}, ugm, UGN, IZZ); 
ram_16x4 rinst_89({&RGE,&RGF,&RGG,&RGH},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_90({&RGM,&RGN,&RGO,&RGP},{WCM,WCN,WCO,WCP},{ugi,ugj,ugk,ugl}, ugm, UGO, IZZ); 
ram_16x4 rinst_91({&RGM,&RGN,&RGO,&RGP},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_92({&RHE,&RHF,&RHG,&RHH},{WDE,WDF,WDG,WDH},{uhi,uhj,uhk,uhl}, uhm, UHN, IZZ); 
ram_16x4 rinst_93({&RHE,&RHF,&RHG,&RHH},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_94({&RHM,&RHN,&RHO,&RHP},{WDM,WDN,WDO,WDP},{uhi,uhj,uhk,uhl}, uhm, UHO, IZZ); 
ram_16x4 rinst_95({&RHM,&RHN,&RHO,&RHP},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_96({&RIE,&RIF,&RIG,&RIH},{WAE,WAF,WAG,WAH},{uii,uii,uik,uil}, uim, UIN, IZZ); 
ram_16x4 rinst_97({&RIE,&RIF,&RIG,&RIH},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_98({&RIM,&RIN,&RIO,&RIP},{WAM,WAN,WAO,WAP},{uii,uij,uik,uil}, uim, UIO, IZZ); 
ram_16x4 rinst_99({&RIM,&RIN,&RIO,&RIP},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_100({&RJE,&RJF,&RJG,&RJH},{WBE,WBF,WBG,WBH},{uji,ujj,ujk,ujl}, ujm, UJN, IZZ); 
ram_16x4 rinst_101({&RJE,&RJF,&RJG,&RJH},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_102({&RJM,&RJN,&RJO,&RJP},{WBM,WBN,WBO,WBP},{uji,ujj,ujk,ujl}, ujm, UJO, IZZ); 
ram_16x4 rinst_103({&RJM,&RJN,&RJO,&RJP},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_104({&RKE,&RKF,&RKG,&RKH},{WCE,WCF,WCG,WCH},{uki,ukj,ukk,ukl}, ukm, UKN, IZZ); 
ram_16x4 rinst_105({&RKE,&RKF,&RKG,&RKH},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_106({&RKM,&RKN,&RKO,&RKP},{WCM,WCN,WCO,WCP},{uki,ukj,ukk,ukl}, ukm, UKO, IZZ); 
ram_16x4 rinst_107({&RKM,&RKN,&RKO,&RKP},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_108({&RLE,&RLF,&RLG,&RLH},{WDE,WDF,WDG,WDH},{uli,ulj,ulk,ull}, ulm, ULN, IZZ); 
ram_16x4 rinst_109({&RLE,&RLF,&RLG,&RLH},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_110({&RLM,&RLN,&RLO,&RLP},{WDM,WDN,WDO,WDP},{uli,ulj,ulk,ull}, ulm, ULO, IZZ); 
ram_16x4 rinst_111({&RLM,&RLN,&RLO,&RLP},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_112({&RME,&RMF,&RMG,&RMH},{WAE,WAF,WAG,WAH},{umi,umi,umk,uml}, umm, UMN, IZZ); 
ram_16x4 rinst_113({&RME,&RMF,&RMG,&RMH},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_114({&RMM,&RMN,&RMO,&RMP},{WAM,WAN,WAO,WAP},{umi,umj,umk,uml}, umm, UMO, IZZ); 
ram_16x4 rinst_115({&RMM,&RMN,&RMO,&RMP},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_116({&RNE,&RNF,&RNG,&RNH},{WBE,WBF,WBG,WBH},{uni,unj,unk,unl}, unm, UNN, IZZ); 
ram_16x4 rinst_117({&RNE,&RNF,&RNG,&RNH},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_118({&RNM,&RNN,&RNO,&RNP},{WBM,WBN,WBO,WBP},{uni,unj,unk,unl}, unm, UNO, IZZ); 
ram_16x4 rinst_119({&RNM,&RNN,&RNO,&RNP},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_120({&ROE,&ROF,&ROG,&ROH},{WCE,WCF,WCG,WCH},{uoi,uoj,uok,uol}, uom, UON, IZZ); 
ram_16x4 rinst_121({&ROE,&ROF,&ROG,&ROH},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_122({&ROM,&RON,&ROO,&ROP},{WCM,WCN,WCO,WCP},{uoi,uoj,uok,uol}, uom, UOO, IZZ); 
ram_16x4 rinst_123({&ROM,&RON,&ROO,&ROP},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_124({&RPE,&RPF,&RPG,&RPH},{WDE,WDF,WDG,WDH},{upi,upj,upk,upl}, upm, UPN, IZZ); 
ram_16x4 rinst_125({&RPE,&RPF,&RPG,&RPH},{,,,},{,,,}, , , IZZ); 
ram_16x4 rinst_126({&RPM,&RPN,&RPO,&RPP},{WDM,WDN,WDO,WDP},{upi,upj,upk,upl}, upm, UPO, IZZ); 
ram_16x4 rinst_127({&RPM,&RPN,&RPO,&RPP},{,,,},{,,,}, , , IZZ); 
endmodule;
