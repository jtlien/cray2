module vr( IZZ,
 IAA, 
 IAB, 
 IAC, 
 IAD, 
 IAE, 
 IAF, 
 IAG, 
 IAH, 
 IBA, 
 IBB, 
 IBC, 
 IBD, 
 IBE, 
 IBF, 
 IBG, 
 IBH, 
 ICA, 
 ICB, 
 ICC, 
 ICD, 
 ICE, 
 ICF, 
 ICG, 
 ICH, 
 IDA, 
 IDB, 
 IDC, 
 IDD, 
 IDE, 
 IDF, 
 IDG, 
 IDH, 
 IEA, 
 IEB, 
 IEC, 
 IED, 
 IEE, 
 IEF, 
 IEG, 
 IEH, 
 IFA, 
 IFB, 
 IFC, 
 IFD, 
 IFE, 
 IFFF , 
 IFG, 
 IFH, 
 IGA, 
 IGB, 
 IGC, 
 IGD, 
 IGE, 
 IGF, 
 IGG, 
 IGH, 
 IHA, 
 IHB, 
 IHC, 
 IHD, 
 IHE, 
 IHF, 
 IHG, 
 IHH, 
 IIA, 
 IIB, 
 IIC, 
 IID, 
 IIE, 
 IIF, 
 IIG, 
 IIH, 
 IJA, 
 IJB, 
 IJC, 
 IJD, 
 IJE, 
 IJF, 
 IJG, 
 IJH, 
 IKA, 
 IKB, 
 IKC, 
 IKD, 
 IKE, 
 IKF, 
 IKG, 
 IKH, 
 IMA, 
 IMB, 
 IMC, 
 IMD, 
 IME, 
 IMF, 
 IMG, 
 IMH, 
 INA, 
 INB, 
 INC, 
 IND, 
 INE, 
 INF, 
 ING, 
 INH, 
 IOA, 
 IOB, 
 IOC, 
 IOD, 
 IOE, 
 IOF, 
 IOG, 
 IOH, 
 IPA, 
 IPB, 
 IPC, 
 IPD, 
 IPE, 
 IPF, 
 IPG, 
 IPH, 
 IQA, 
 IQB, 
 IQC, 
 IQD, 
 IQE, 
 IQF, 
 IQG, 
 IQH, 
 IRA, 
 IRB, 
 IRC, 
 IRD, 
 IRE, 
 IRF, 
 IRG, 
 IRH, 
 ISA, 
 ISB, 
 ISC, 
 ISD, 
 ISE, 
 ISF, 
 ISG, 
 ITA, 
 ITB, 
 ITC, 
 ITD, 
 ITE, 
 ITF, 
 OAA, 
 OAB, 
 OAC, 
 OAD, 
 OAE, 
 OAF, 
 OAG, 
 OAH, 
 OBA, 
 OBB, 
 OBC, 
 OBD, 
 OBE, 
 OBF, 
 OBG, 
 OBH, 
 OCA, 
 OCB, 
 OCC, 
 OCD, 
 OCE, 
 OCF, 
 OCG, 
 OCH, 
 ODA, 
 ODB, 
 ODC, 
 ODD, 
 ODE, 
 ODF, 
 ODG, 
 ODH, 
 OEA, 
 OEB, 
 OEC, 
 OED, 
 OEE, 
 OEF, 
 OEG, 
 OEH, 
 OFA, 
 OFB, 
 OFC, 
 OFD, 
 OFE, 
 OFF, 
 OFG, 
 OFH, 
 OGA, 
 OGB, 
 OGC, 
 OGD, 
 OGE, 
 OGF, 
 OGG, 
 OGH, 
 OHA, 
 OHB, 
 OHC, 
 OHD, 
 OHE, 
 OHF, 
 OHG, 
 OHH, 
 OIA, 
 OIB, 
 OIC, 
 OID, 
 OIE, 
 OIF, 
 OIG, 
 OIH, 
 OJA, 
 OJB, 
 OJC, 
 OJD, 
 OJE, 
 OJF, 
 OJG, 
 OJH, 
 OKA, 
 OKB, 
 OKC, 
 OKD, 
 OKE, 
 OKF, 
 OKG, 
 OKH, 
 OLA, 
 OLB, 
 OLC, 
 OLD, 
 OLE, 
 OLF, 
 OLG, 
 OLH, 
 OMA, 
 OMB, 
 OMC, 
 OMD, 
 OME, 
 OMF, 
 OMG, 
 OMH, 
 ONA, 
 ONB, 
 ONC, 
 OND, 
 ONE, 
 ONF, 
 ONG, 
 ONH, 
 OOA, 
 OOB, 
 OOC, 
 OOD, 
 OOE, 
 OOF, 
 OOG, 
 OOH, 
 OQA, 
 OQB, 
ORA ); 
    
 input IZZ; 
 input IAA; 
 input IAB; 
 input IAC; 
 input IAD; 
 input IAE; 
 input IAF; 
 input IAG; 
 input IAH; 
 input IBA; 
 input IBB; 
 input IBC; 
 input IBD; 
 input IBE; 
 input IBF; 
 input IBG; 
 input IBH; 
 input ICA; 
 input ICB; 
 input ICC; 
 input ICD; 
 input ICE; 
 input ICF; 
 input ICG; 
 input ICH; 
 input IDA; 
 input IDB; 
 input IDC; 
 input IDD; 
 input IDE; 
 input IDF; 
 input IDG; 
 input IDH; 
 input IEA; 
 input IEB; 
 input IEC; 
 input IED; 
 input IEE; 
 input IEF; 
 input IEG; 
 input IEH; 
 input IFA; 
 input IFB; 
 input IFC; 
 input IFD; 
 input IFE; 
 input IFFF ; 
 input IFG; 
 input IFH; 
 input IGA; 
 input IGB; 
 input IGC; 
 input IGD; 
 input IGE; 
 input IGF; 
 input IGG; 
 input IGH; 
 input IHA; 
 input IHB; 
 input IHC; 
 input IHD; 
 input IHE; 
 input IHF; 
 input IHG; 
 input IHH; 
 input IIA; 
 input IIB; 
 input IIC; 
 input IID; 
 input IIE; 
 input IIF; 
 input IIG; 
 input IIH; 
 input IJA; 
 input IJB; 
 input IJC; 
 input IJD; 
 input IJE; 
 input IJF; 
 input IJG; 
 input IJH; 
 input IKA; 
 input IKB; 
 input IKC; 
 input IKD; 
 input IKE; 
 input IKF; 
 input IKG; 
 input IKH; 
 input IMA; 
 input IMB; 
 input IMC; 
 input IMD; 
 input IME; 
 input IMF; 
 input IMG; 
 input IMH; 
 input INA; 
 input INB; 
 input INC; 
 input IND; 
 input INE; 
 input INF; 
 input ING; 
 input INH; 
 input IOA; 
 input IOB; 
 input IOC; 
 input IOD; 
 input IOE; 
 input IOF; 
 input IOG; 
 input IOH; 
 input IPA; 
 input IPB; 
 input IPC; 
 input IPD; 
 input IPE; 
 input IPF; 
 input IPG; 
 input IPH; 
 input IQA; 
 input IQB; 
 input IQC; 
 input IQD; 
 input IQE; 
 input IQF; 
 input IQG; 
 input IQH; 
 input IRA; 
 input IRB; 
 input IRC; 
 input IRD; 
 input IRE; 
 input IRF; 
 input IRG; 
 input IRH; 
 input ISA; 
 input ISB; 
 input ISC; 
 input ISD; 
 input ISE; 
 input ISF; 
 input ISG; 
 input ITA; 
 input ITB; 
 input ITC; 
 input ITD; 
 input ITE; 
 input ITF; 
 output OAA; 
 output OAB; 
 output OAC; 
 output OAD; 
 output OAE; 
 output OAF; 
 output OAG; 
 output OAH; 
 output OBA; 
 output OBB; 
 output OBC; 
 output OBD; 
 output OBE; 
 output OBF; 
 output OBG; 
 output OBH; 
 output OCA; 
 output OCB; 
 output OCC; 
 output OCD; 
 output OCE; 
 output OCF; 
 output OCG; 
 output OCH; 
 output ODA; 
 output ODB; 
 output ODC; 
 output ODD; 
 output ODE; 
 output ODF; 
 output ODG; 
 output ODH; 
 output OEA; 
 output OEB; 
 output OEC; 
 output OED; 
 output OEE; 
 output OEF; 
 output OEG; 
 output OEH; 
 output OFA; 
 output OFB; 
 output OFC; 
 output OFD; 
 output OFE; 
 output OFF; 
 output OFG; 
 output OFH; 
 output OGA; 
 output OGB; 
 output OGC; 
 output OGD; 
 output OGE; 
 output OGF; 
 output OGG; 
 output OGH; 
 output OHA; 
 output OHB; 
 output OHC; 
 output OHD; 
 output OHE; 
 output OHF; 
 output OHG; 
 output OHH; 
 output OIA; 
 output OIB; 
 output OIC; 
 output OID; 
 output OIE; 
 output OIF; 
 output OIG; 
 output OIH; 
 output OJA; 
 output OJB; 
 output OJC; 
 output OJD; 
 output OJE; 
 output OJF; 
 output OJG; 
 output OJH; 
 output OKA; 
 output OKB; 
 output OKC; 
 output OKD; 
 output OKE; 
 output OKF; 
 output OKG; 
 output OKH; 
 output OLA; 
 output OLB; 
 output OLC; 
 output OLD; 
 output OLE; 
 output OLF; 
 output OLG; 
 output OLH; 
 output OMA; 
 output OMB; 
 output OMC; 
 output OMD; 
 output OME; 
 output OMF; 
 output OMG; 
 output OMH; 
 output ONA; 
 output ONB; 
 output ONC; 
 output OND; 
 output ONE; 
 output ONF; 
 output ONG; 
 output ONH; 
 output OOA; 
 output OOB; 
 output OOC; 
 output OOD; 
 output OOE; 
 output OOF; 
 output OOG; 
 output OOH; 
 output OQA; 
 output OQB; 
 output ORA; 
  
  
reg  AAA ;
reg  AAB ;
reg  AAC ;
reg  AAD ;
reg  AAE ;
reg  AAF ;
reg  AAG ;
reg  aba ;
reg  abb ;
reg  abc ;
reg  BAD ;
reg  BAE ;
reg  BAF ;
reg  BAJ ;
reg  BAK ;
reg  BAL ;
reg  BAM ;
reg  BAN ;
reg  BAO ;
reg  BAP ;
reg  BBA ;
reg  BBB ;
reg  BBC ;
reg  CAA ;
reg  CAB ;
reg  CAC ;
reg  CAD ;
reg  cae ;
reg  caf ;
reg  cag ;
reg  cah ;
reg  cai ;
reg  caj ;
reg  DAC ;
reg  DAD ;
reg  DAE ;
reg  DAF ;
reg  DAG ;
reg  dai ;
reg  daj ;
reg  dak ;
reg  dal ;
reg  DAM ;
reg  DAN ;
reg  DAO ;
reg  DAP ;
reg  DBC ;
reg  DBD ;
reg  DBE ;
reg  DBF ;
reg  DBG ;
reg  dbi ;
reg  dbj ;
reg  dbk ;
reg  dbl ;
reg  DBM ;
reg  DBN ;
reg  DBO ;
reg  DBP ;
reg  DCC ;
reg  DCD ;
reg  DCE ;
reg  DCF ;
reg  DCG ;
reg  dci ;
reg  dcj ;
reg  dck ;
reg  dcl ;
reg  DCM ;
reg  DCN ;
reg  DCO ;
reg  DCP ;
reg  DDC ;
reg  DDD ;
reg  DDE ;
reg  DDF ;
reg  DDG ;
reg  ddi ;
reg  ddj ;
reg  ddk ;
reg  ddl ;
reg  DDM ;
reg  DDN ;
reg  DDO ;
reg  DDP ;
reg  DEC ;
reg  DED ;
reg  DEE ;
reg  DEF ;
reg  DEG ;
reg  dei ;
reg  dej ;
reg  dek ;
reg  del ;
reg  DEM ;
reg  DEN ;
reg  DEO ;
reg  DEP ;
reg  DFC ;
reg  DFD ;
reg  DFE ;
reg  DFF ;
reg  DFG ;
reg  dfi ;
reg  dfj ;
reg  dfk ;
reg  dfl ;
reg  DFM ;
reg  DFN ;
reg  DFO ;
reg  DFP ;
reg  DGC ;
reg  DGD ;
reg  DGE ;
reg  DGF ;
reg  DGG ;
reg  dgi ;
reg  dgj ;
reg  dgk ;
reg  dgl ;
reg  DGM ;
reg  DGN ;
reg  DGO ;
reg  DGP ;
reg  DHC ;
reg  DHD ;
reg  DHE ;
reg  DHF ;
reg  DHG ;
reg  dhi ;
reg  dhj ;
reg  dhk ;
reg  dhl ;
reg  DHM ;
reg  DHN ;
reg  DHO ;
reg  DHP ;
reg  GAA ;
reg  GAB ;
reg  GAC ;
reg  GAD ;
reg  GAE ;
reg  GAF ;
reg  GAG ;
reg  GAH ;
reg  GAI ;
reg  GAJ ;
reg  GAK ;
reg  GAL ;
reg  GAM ;
reg  GAN ;
reg  GAO ;
reg  GAP ;
reg  GBA ;
reg  GBB ;
reg  GBC ;
reg  GBD ;
reg  GBE ;
reg  GBF ;
reg  GBG ;
reg  GBH ;
reg  GBI ;
reg  GBJ ;
reg  GBK ;
reg  GBL ;
reg  GBM ;
reg  GBN ;
reg  GBO ;
reg  GBP ;
reg  kaa ;
reg  kab ;
reg  kac ;
reg  kad ;
reg  kae ;
reg  kaf ;
reg  kag ;
reg  kah ;
reg  kba ;
reg  kbb ;
reg  kbc ;
reg  kbd ;
reg  kbe ;
reg  kbf ;
reg  kbg ;
reg  kbh ;
reg  kca ;
reg  kcb ;
reg  kcc ;
reg  kcd ;
reg  kce ;
reg  kcf ;
reg  kcg ;
reg  kch ;
reg  kda ;
reg  kdb ;
reg  kdc ;
reg  kdd ;
reg  kde ;
reg  kdf ;
reg  kdg ;
reg  kdh ;
reg  kea ;
reg  keb ;
reg  kec ;
reg  ked ;
reg  kee ;
reg  kef ;
reg  keg ;
reg  keh ;
reg  kfa ;
reg  kfb ;
reg  kfc ;
reg  kfd ;
reg  kfe ;
reg  kff ;
reg  kfg ;
reg  kfh ;
reg  LAA ;
reg  LAB ;
reg  LAC ;
reg  LBA ;
reg  LBB ;
reg  LBC ;
reg  LCA ;
reg  LCB ;
reg  LCC ;
reg  LDA ;
reg  LDB ;
reg  LDC ;
reg  LEA ;
reg  LEB ;
reg  LEC ;
reg  LFA ;
reg  LFB ;
reg  LFC ;
reg  LGA ;
reg  LGB ;
reg  LGC ;
reg  LHA ;
reg  LHB ;
reg  LHC ;
reg  LIA ;
reg  LIB ;
reg  LIC ;
reg  LJA ;
reg  LJB ;
reg  LJC ;
reg  LKA ;
reg  LKB ;
reg  LKC ;
reg  LLA ;
reg  LLB ;
reg  LLC ;
reg  LMA ;
reg  LMB ;
reg  LMC ;
reg  LNA ;
reg  LNB ;
reg  LNC ;
reg  LOA ;
reg  LOB ;
reg  LOC ;
reg  LPA ;
reg  LPB ;
reg  LPC ;
reg  LQA ;
reg  LQB ;
reg  LQC ;
reg  LRA ;
reg  LRB ;
reg  LRC ;
reg  LSA ;
reg  LSB ;
reg  LSC ;
reg  LTA ;
reg  LTB ;
reg  LTC ;
reg  NAA ;
reg  NAB ;
reg  NAC ;
reg  NAD ;
reg  NBA ;
reg  NBB ;
reg  NBC ;
reg  NBD ;
reg  NCA ;
reg  NCB ;
reg  NCC ;
reg  NCD ;
reg  NDA ;
reg  NDB ;
reg  NDC ;
reg  NDD ;
reg  NEA ;
reg  NEB ;
reg  NEC ;
reg  NED ;
reg  NFA ;
reg  NFB ;
reg  NFC ;
reg  NFD ;
reg  NGA ;
reg  NGB ;
reg  NGC ;
reg  NGD ;
reg  NHA ;
reg  NHB ;
reg  NHC ;
reg  NHD ;
reg  oaa ;
reg  oab ;
reg  oac ;
reg  oad ;
reg  oae ;
reg  oaf ;
reg  oag ;
reg  oah ;
reg  oba ;
reg  obb ;
reg  obc ;
reg  obd ;
reg  obe ;
reg  obf ;
reg  obg ;
reg  obh ;
reg  oca ;
reg  ocb ;
reg  occ ;
reg  ocd ;
reg  oce ;
reg  ocf ;
reg  ocg ;
reg  och ;
reg  ODA ;
reg  ODB ;
reg  ODC ;
reg  ODD ;
reg  ODE ;
reg  ODF ;
reg  ODG ;
reg  ODH ;
reg  OEA ;
reg  OEB ;
reg  OEC ;
reg  OED ;
reg  OEE ;
reg  OEF ;
reg  OEG ;
reg  OEH ;
reg  OFA ;
reg  OFB ;
reg  OFC ;
reg  OFD ;
reg  OFE ;
reg  OFF ;
reg  OFG ;
reg  OFH ;
reg  OGA ;
reg  OGB ;
reg  OGC ;
reg  OGD ;
reg  OGE ;
reg  OGF ;
reg  OGG ;
reg  OGH ;
reg  OHA ;
reg  OHB ;
reg  OHC ;
reg  OHD ;
reg  OHE ;
reg  OHF ;
reg  OHG ;
reg  OHH ;
reg  OIA ;
reg  OIB ;
reg  OIC ;
reg  OID ;
reg  OIE ;
reg  OIF ;
reg  OIG ;
reg  OIH ;
reg  OJA ;
reg  OJB ;
reg  OJC ;
reg  OJD ;
reg  OJE ;
reg  OJF ;
reg  OJG ;
reg  OJH ;
reg  OKA ;
reg  OKB ;
reg  OKC ;
reg  OKD ;
reg  OKE ;
reg  OKF ;
reg  OKG ;
reg  OKH ;
reg  OLA ;
reg  OLB ;
reg  OLC ;
reg  OLD ;
reg  OLE ;
reg  OLF ;
reg  OLG ;
reg  OLH ;
reg  OMA ;
reg  OMB ;
reg  OMC ;
reg  OMD ;
reg  OME ;
reg  OMF ;
reg  OMG ;
reg  OMH ;
reg  ONA ;
reg  ONB ;
reg  ONC ;
reg  OND ;
reg  ONE ;
reg  ONF ;
reg  ONG ;
reg  ONH ;
reg  OOA ;
reg  OOB ;
reg  OOC ;
reg  OOD ;
reg  OOE ;
reg  OOF ;
reg  OOG ;
reg  OOH ;
reg  oqa ;
reg  OQB ;
reg  ORA ;
reg  QAA ;
reg  QAB ;
reg  QAC ;
reg  QBA ;
reg  qca ;
reg  qcb ;
reg  qcc ;
reg  QDA ;
reg  QDB ;
reg  QDC ;
reg  QEA ;
reg  QEB ;
reg  QEC ;
reg  SAA ;
reg  SAB ;
reg  SAC ;
reg  SAD ;
reg  SAE ;
reg  SAF ;
reg  SAG ;
reg  SAH ;
reg  SBA ;
reg  SBB ;
reg  SBC ;
reg  SBD ;
reg  SBE ;
reg  SBF ;
reg  SBG ;
reg  SBH ;
reg  SCA ;
reg  SCB ;
reg  SCC ;
reg  SCD ;
reg  SCE ;
reg  SCF ;
reg  SCG ;
reg  SCH ;
reg  SDA ;
reg  SDB ;
reg  SDC ;
reg  SDD ;
reg  SDE ;
reg  SDF ;
reg  SDG ;
reg  SDH ;
reg  SEA ;
reg  SEB ;
reg  SEC ;
reg  SED ;
reg  SEE ;
reg  SEF ;
reg  SEG ;
reg  SEH ;
reg  SFA ;
reg  SFB ;
reg  SFC ;
reg  SFD ;
reg  SFE ;
reg  SFF ;
reg  SFG ;
reg  SFH ;
reg  SGA ;
reg  SGB ;
reg  SGC ;
reg  SGD ;
reg  SGE ;
reg  SGF ;
reg  SGG ;
reg  SGH ;
reg  SHA ;
reg  SHB ;
reg  SHC ;
reg  SHD ;
reg  SHE ;
reg  SHF ;
reg  SHG ;
reg  SHH ;
reg  SJA ;
reg  SJB ;
reg  SJC ;
reg  SJD ;
reg  SJE ;
reg  SJF ;
reg  SJG ;
reg  SJH ;
reg  ska ;
reg  skb ;
reg  skc ;
reg  skd ;
reg  ske ;
reg  skf ;
reg  skg ;
reg  skh ;
reg  TAA ;
reg  TAB ;
reg  TAC ;
reg  TAD ;
reg  TBA ;
reg  TBB ;
reg  TBC ;
reg  TBD ;
reg  TCA ;
reg  TCB ;
reg  TCC ;
reg  TCD ;
reg  TDA ;
reg  TDB ;
reg  TDC ;
reg  TDD ;
reg  TEA ;
reg  TEB ;
reg  TEC ;
reg  TED ;
reg  TFA ;
reg  TFB ;
reg  TFC ;
reg  TFD ;
reg  TGA ;
reg  TGB ;
reg  TGC ;
reg  TGD ;
reg  THA ;
reg  THB ;
reg  THC ;
reg  THD ;
reg  TIB ;
reg  TIC ;
reg  TID ;
reg  TIE ;
reg  TIF ;
reg  TIG ;
reg  TJB ;
reg  TJC ;
reg  TJD ;
reg  TJE ;
reg  TJF ;
reg  TJG ;
reg  TKB ;
reg  TKC ;
reg  TKD ;
reg  TKE ;
reg  TKF ;
reg  TKG ;
reg  TSA ;
reg  TSB ;
reg  TSC ;
reg  TSD ;
reg  TSE ;
reg  TSF ;
reg  TSG ;
reg  TSH ;
reg  UAA ;
reg  UAB ;
reg  UAC ;
reg  UAD ;
reg  UAE ;
reg  UAF ;
reg  UAG ;
reg  UAH ;
reg  UAI ;
reg  UAJ ;
reg  UAK ;
reg  UAL ;
reg  UAM ;
reg  UAN ;
reg  UAO ;
reg  UAP ;
reg  UAQ ;
reg  UAR ;
reg  UAS ;
reg  UAT ;
reg  UAU ;
reg  UAV ;
reg  UAW ;
reg  UAX ;
reg  UBA ;
reg  UBB ;
reg  UBC ;
reg  UBD ;
reg  UBE ;
reg  UBF ;
reg  UBG ;
reg  UBH ;
reg  UBI ;
reg  UBJ ;
reg  UBK ;
reg  UBL ;
reg  UBM ;
reg  UBN ;
reg  UBO ;
reg  UBP ;
reg  UBQ ;
reg  UBR ;
reg  UBS ;
reg  UBT ;
reg  UBU ;
reg  UBV ;
reg  UBW ;
reg  UBX ;
reg  UCA ;
reg  UCB ;
reg  UCC ;
reg  UCD ;
reg  UCE ;
reg  UCF ;
reg  UCG ;
reg  UCH ;
reg  UCI ;
reg  UCJ ;
reg  UCK ;
reg  UCL ;
reg  UCM ;
reg  UCN ;
reg  UCO ;
reg  UCP ;
reg  UCQ ;
reg  UCR ;
reg  UCS ;
reg  UCT ;
reg  UCU ;
reg  UCV ;
reg  UCW ;
reg  UCX ;
reg  UDA ;
reg  UDB ;
reg  UDC ;
reg  UDD ;
reg  UDE ;
reg  UDF ;
reg  UDG ;
reg  UDH ;
reg  UDI ;
reg  UDJ ;
reg  UDK ;
reg  UDL ;
reg  UDM ;
reg  UDN ;
reg  UDO ;
reg  UDP ;
reg  UDQ ;
reg  UDR ;
reg  UDS ;
reg  UDT ;
reg  UDU ;
reg  UDV ;
reg  UDW ;
reg  UDX ;
reg  UEA ;
reg  UEB ;
reg  UEC ;
reg  UED ;
reg  UEE ;
reg  UEF ;
reg  UEG ;
reg  UEH ;
reg  UEI ;
reg  UEJ ;
reg  UEK ;
reg  UEL ;
reg  UEM ;
reg  UEN ;
reg  UEO ;
reg  UEP ;
reg  UEQ ;
reg  UER ;
reg  UES ;
reg  UET ;
reg  UEU ;
reg  UEV ;
reg  UEW ;
reg  UEX ;
reg  UFA ;
reg  UFB ;
reg  UFC ;
reg  UFD ;
reg  UFE ;
reg  UFF ;
reg  UFG ;
reg  UFH ;
reg  UFI ;
reg  UFJ ;
reg  UFK ;
reg  UFL ;
reg  UFM ;
reg  UFN ;
reg  UFO ;
reg  UFP ;
reg  UFQ ;
reg  UFR ;
reg  UFS ;
reg  UFT ;
reg  UFU ;
reg  UFV ;
reg  UFW ;
reg  UFX ;
reg  UGA ;
reg  UGB ;
reg  UGC ;
reg  UGD ;
reg  UGE ;
reg  UGF ;
reg  UGG ;
reg  UGH ;
reg  UGI ;
reg  UGJ ;
reg  UGK ;
reg  UGL ;
reg  UGM ;
reg  UGN ;
reg  UGO ;
reg  UGP ;
reg  UGQ ;
reg  UGR ;
reg  UGS ;
reg  UGT ;
reg  UGU ;
reg  UGV ;
reg  UGW ;
reg  UGX ;
reg  UHA ;
reg  UHB ;
reg  UHC ;
reg  UHD ;
reg  UHE ;
reg  UHF ;
reg  UHG ;
reg  UHH ;
reg  UHI ;
reg  UHJ ;
reg  UHK ;
reg  UHL ;
reg  UHM ;
reg  UHN ;
reg  UHO ;
reg  UHP ;
reg  UHQ ;
reg  UHR ;
reg  UHS ;
reg  UHT ;
reg  UHU ;
reg  UHV ;
reg  UHW ;
reg  UHX ;
reg  VAA ;
reg  VAB ;
reg  VAC ;
reg  VAD ;
reg  VAE ;
reg  VAF ;
reg  VAG ;
reg  VAH ;
reg  VAI ;
reg  VAJ ;
reg  VAK ;
reg  VAL ;
reg  VAM ;
reg  VAN ;
reg  VAO ;
reg  VAP ;
reg  VBA ;
reg  VBB ;
reg  VBC ;
reg  VBD ;
reg  VBE ;
reg  VBF ;
reg  VBG ;
reg  VBH ;
reg  VBI ;
reg  VBJ ;
reg  VBK ;
reg  VBL ;
reg  VBM ;
reg  VBN ;
reg  VBO ;
reg  VBP ;
reg  VCA ;
reg  VCB ;
reg  VCC ;
reg  VCD ;
reg  VCE ;
reg  VCF ;
reg  VCG ;
reg  VCH ;
reg  VCI ;
reg  VCJ ;
reg  VCK ;
reg  VCL ;
reg  VCM ;
reg  VCN ;
reg  VCO ;
reg  VCP ;
reg  VDA ;
reg  VDB ;
reg  VDC ;
reg  VDD ;
reg  VDE ;
reg  VDF ;
reg  VDG ;
reg  VDH ;
reg  VDI ;
reg  VDJ ;
reg  VDK ;
reg  VDL ;
reg  VDM ;
reg  VDN ;
reg  VDO ;
reg  VDP ;
reg  VEA ;
reg  VEB ;
reg  VEC ;
reg  VED ;
reg  VEE ;
reg  VEF ;
reg  VEG ;
reg  VEH ;
reg  VEI ;
reg  VEJ ;
reg  VEK ;
reg  VEL ;
reg  VEM ;
reg  VEN ;
reg  VEO ;
reg  VEP ;
reg  VFA ;
reg  VFB ;
reg  VFC ;
reg  VFD ;
reg  VFE ;
reg  VFF ;
reg  VFG ;
reg  VFH ;
reg  VFI ;
reg  VFJ ;
reg  VFK ;
reg  VFL ;
reg  VFM ;
reg  VFN ;
reg  VFO ;
reg  VFP ;
reg  VGA ;
reg  VGB ;
reg  VGC ;
reg  VGD ;
reg  VGE ;
reg  VGF ;
reg  VGG ;
reg  VGH ;
reg  VGI ;
reg  VGJ ;
reg  VGK ;
reg  VGL ;
reg  VGM ;
reg  VGN ;
reg  VGO ;
reg  VGP ;
reg  VHA ;
reg  VHB ;
reg  VHC ;
reg  VHD ;
reg  VHE ;
reg  VHF ;
reg  VHG ;
reg  VHH ;
reg  VHI ;
reg  VHJ ;
reg  VHK ;
reg  VHL ;
reg  VHM ;
reg  VHN ;
reg  VHO ;
reg  VHP ;

reg  WAA ;
reg  WAB ;
reg  WAC ;
reg  WAD ;
reg  WAE ;
reg  WAF ;
reg  WAG ;
reg  WAH ;
reg  WBA ;
reg  WBB ;
reg  WBC ;
reg  WBD ;
reg  WBE ;
reg  WBF ;
reg  WBG ;
reg  WBH ;
reg  WCA ;
reg  WCB ;
reg  WCC ;
reg  WCD ;
reg  WCE ;
reg  WCF ;
reg  WCG ;
reg  WCH ;
reg  WDA ;
reg  WDB ;
reg  WDC ;
reg  WDD ;
reg  WDE ;
reg  WDF ;
reg  WDG ;
reg  WDH ;
reg  WEA ;
reg  WEB ;
reg  WEC ;
reg  WED ;
reg  WEE ;
reg  WEF ;
reg  WEG ;
reg  WEH ;
reg  WFA ;
reg  WFB ;
reg  WFC ;
reg  WFD ;
reg  WFE ;
reg  WFF ;
reg  WFG ;
reg  WFH ;
reg  WGA ;
reg  WGB ;
reg  WGC ;
reg  WGD ;
reg  WGE ;
reg  WGF ;
reg  WGG ;
reg  WGH ;
reg  WHA ;
reg  WHB ;
reg  WHC ;
reg  WHD ;
reg  WHE ;
reg  WHF ;
reg  WHG ;
reg  WHH ;
wire  aaa ;
wire  aab ;
wire  aac ;
wire  aad ;
wire  aae ;
wire  aaf ;
wire  aag ;
wire  ABA ;
wire  ABB ;
wire  ABC ;
wire  bad ;
wire  bae ;
wire  baf ;
wire  baj ;
wire  bak ;
wire  bal ;
wire  bam ;
wire  ban ;
wire  bao ;
wire  bap ;
wire  bba ;
wire  bbb ;
wire  bbc ;
wire  caa ;
wire  cab ;
wire  cac ;
wire  cad ;
wire  CAE ;
wire  CAF ;
wire  CAG ;
wire  CAH ;
wire  CAI ;
wire  CAJ ;
wire  dac ;
wire  dad ;
wire  dae ;
wire  daf ;
wire  dag ;
wire  DAI ;
wire  DAJ ;
wire  DAK ;
wire  DAL ;
wire  dam ;
wire  dan ;
wire  dao ;
wire  dap ;
wire  dbc ;
wire  dbd ;
wire  dbe ;
wire  dbf ;
wire  dbg ;
wire  DBI ;
wire  DBJ ;
wire  DBK ;
wire  DBL ;
wire  dbm ;
wire  dbn ;
wire  dbo ;
wire  dbp ;
wire  dcc ;
wire  dcd ;
wire  dce ;
wire  dcf ;
wire  dcg ;
wire  DCI ;
wire  DCJ ;
wire  DCK ;
wire  DCL ;
wire  dcm ;
wire  dcn ;
wire  dco ;
wire  dcp ;
wire  ddc ;
wire  ddd ;
wire  dde ;
wire  ddf ;
wire  ddg ;
wire  DDI ;
wire  DDJ ;
wire  DDK ;
wire  DDL ;
wire  ddm ;
wire  ddn ;
wire  ddo ;
wire  ddp ;
wire  dec ;
wire  ded ;
wire  dee ;
wire  def ;
wire  deg ;
wire  DEI ;
wire  DEJ ;
wire  DEK ;
wire  DEL ;
wire  dem ;
wire  den ;
wire  deo ;
wire  dep ;
wire  dfc ;
wire  dfd ;
wire  dfe ;
wire  dff ;
wire  dfg ;
wire  DFI ;
wire  DFJ ;
wire  DFK ;
wire  DFL ;
wire  dfm ;
wire  dfn ;
wire  dfo ;
wire  dfp ;
wire  dgc ;
wire  dgd ;
wire  dge ;
wire  dgf ;
wire  dgg ;
wire  DGI ;
wire  DGJ ;
wire  DGK ;
wire  DGL ;
wire  dgm ;
wire  dgn ;
wire  dgo ;
wire  dgp ;
wire  dhc ;
wire  dhd ;
wire  dhe ;
wire  dhf ;
wire  dhg ;
wire  DHI ;
wire  DHJ ;
wire  DHK ;
wire  DHL ;
wire  dhm ;
wire  dhn ;
wire  dho ;
wire  dhp ;
wire  eaa ;
wire  EAA ;
wire  eab ;
wire  EAB ;
wire  eac ;
wire  EAC ;
wire  ead ;
wire  EAD ;
wire  eae ;
wire  EAE ;
wire  FAA ;
wire  FAB ;
wire  FAC ;
wire  FAD ;
wire  FAE ;
wire  FAF ;
wire  FAG ;
wire  FAH ;
wire  FAI ;
wire  FBA ;
wire  FBB ;
wire  FBC ;
wire  FBD ;
wire  FBE ;
wire  FBF ;
wire  FBG ;
wire  FBH ;
wire  FBI ;
wire  FCA ;
wire  FCB ;
wire  FCC ;
wire  FCD ;
wire  FCE ;
wire  FCF ;
wire  FCG ;
wire  FCH ;
wire  FCI ;
wire  FDA ;
wire  FDB ;
wire  FDC ;
wire  FDD ;
wire  FDE ;
wire  FDF ;
wire  FDG ;
wire  FDH ;
wire  FDI ;
wire  FEA ;
wire  FEB ;
wire  FEC ;
wire  FED ;
wire  FEE ;
wire  FEF ;
wire  FEG ;
wire  FEH ;
wire  FEI ;
wire fda;
wire fdb;
wire fdc;
wire fdd;
wire fde;
wire fdf;
wire fdg;
wire fdh;
   
wire  gaa ;
wire  gab ;
wire  gac ;
wire  gad ;
wire  gae ;
wire  gaf ;
wire  gag ;
wire  gah ;
wire  gai ;
wire  gaj ;
wire  gak ;
wire  gal ;
wire  gam ;
wire  gan ;
wire  gao ;
wire  gap ;
wire  gba ;
wire  gbb ;
wire  gbc ;
wire  gbd ;
wire  gbe ;
wire  gbf ;
wire  gbg ;
wire  gbh ;
wire  gbi ;
wire  gbj ;
wire  gbk ;
wire  gbl ;
wire  gbm ;
wire  gbn ;
wire  gbo ;
wire  gbp ;
wire  haa ;
wire  HAA ;
wire  hab ;
wire  HAB ;
wire  hac ;
wire  HAC ;
wire  had ;
wire  HAD ;
wire  hae ;
wire  HAE ;
wire  haf ;
wire  HAF ;
wire  hag ;
wire  HAG ;
wire  hah ;
wire  HAH ;
wire  hai ;
wire  HAI ;
wire  haj ;
wire  HAJ ;
wire  hak ;
wire  HAK ;
wire  hal ;
wire  HAL ;
wire  ham ;
wire  HAM ;
wire  han ;
wire  HAN ;
wire  hao ;
wire  HAO ;
wire  hap ;
wire  HAP ;
wire  hba ;
wire  HBA ;
wire  hbb ;
wire  HBB ;
wire  hbc ;
wire  HBC ;
wire  hbd ;
wire  HBD ;
wire  hbe ;
wire  HBE ;
wire  hbf ;
wire  HBF ;
wire  hbg ;
wire  HBG ;
wire  hbh ;
wire  HBH ;
wire  hbi ;
wire  HBI ;
wire  hbj ;
wire  HBJ ;
wire  hbk ;
wire  HBK ;
wire  hbl ;
wire  HBL ;
wire  hbm ;
wire  HBM ;
wire  hbn ;
wire  HBN ;
wire  hbo ;
wire  HBO ;
wire  hbp ;
wire  HBP ;
wire  hca ;
wire  HCA ;
wire  hcb ;
wire  HCB ;
wire  hcc ;
wire  HCC ;
wire  hcd ;
wire  HCD ;
wire  hce ;
wire  HCE ;
wire  hcf ;
wire  HCF ;
wire  hcg ;
wire  HCG ;
wire  hch ;
wire  HCH ;
wire  hci ;
wire  HCI ;
wire  hcj ;
wire  HCJ ;
wire  hck ;
wire  HCK ;
wire  hcl ;
wire  HCL ;
wire  hcm ;
wire  HCM ;
wire  hcn ;
wire  HCN ;
wire  hco ;
wire  HCO ;
wire  hcp ;
wire  HCP ;
wire  hda ;
wire  HDA ;
wire  hdb ;
wire  HDB ;
wire  hdc ;
wire  HDC ;
wire  hdd ;
wire  HDD ;
wire  hde ;
wire  HDE ;
wire  hdf ;
wire  HDF ;
wire  hdg ;
wire  HDG ;
wire  hdh ;
wire  HDH ;
wire  hdi ;
wire  HDI ;
wire  hdj ;
wire  HDJ ;
wire  hdk ;
wire  HDK ;
wire  hdl ;
wire  HDL ;
wire  hdm ;
wire  HDM ;
wire  hdn ;
wire  HDN ;
wire  hdo ;
wire  HDO ;
wire  hdp ;
wire  HDP ;
wire  hea ;
wire  HEA ;
wire  heb ;
wire  HEB ;
wire  hec ;
wire  HEC ;
wire  hed ;
wire  HED ;
wire  hee ;
wire  HEE ;
wire  hef ;
wire  HEF ;
wire  heg ;
wire  HEG ;
wire  heh ;
wire  HEH ;
wire  hei ;
wire  HEI ;
wire  hej ;
wire  HEJ ;
wire  hek ;
wire  HEK ;
wire  hel ;
wire  HEL ;
wire  hem ;
wire  HEM ;
wire  hen ;
wire  HEN ;
wire  heo ;
wire  HEO ;
wire  hep ;
wire  HEP ;
wire  hfa ;
wire  HFA ;
wire  hfb ;
wire  HFB ;
wire  hfc ;
wire  HFC ;
wire  hfd ;
wire  HFD ;
wire  hfe ;
wire  HFE ;
wire  hff ;
wire  HFF ;
wire  hfg ;
wire  HFG ;
wire  hfh ;
wire  HFH ;
wire  hfi ;
wire  HFI ;
wire  hfj ;
wire  HFJ ;
wire  hfk ;
wire  HFK ;
wire  hfl ;
wire  HFL ;
wire  hfm ;
wire  HFM ;
wire  hfn ;
wire  HFN ;
wire  hfo ;
wire  HFO ;
wire  hfp ;
wire  HFP ;
wire  hga ;
wire  HGA ;
wire  hgb ;
wire  HGB ;
wire  hgc ;
wire  HGC ;
wire  hgd ;
wire  HGD ;
wire  hge ;
wire  HGE ;
wire  hgf ;
wire  HGF ;
wire  hgg ;
wire  HGG ;
wire  hgh ;
wire  HGH ;
wire  hgi ;
wire  HGI ;
wire  hgj ;
wire  HGJ ;
wire  hgk ;
wire  HGK ;
wire  hgl ;
wire  HGL ;
wire  hgm ;
wire  HGM ;
wire  hgn ;
wire  HGN ;
wire  hgo ;
wire  HGO ;
wire  hgp ;
wire  HGP ;
wire  hha ;
wire  HHA ;
wire  hhb ;
wire  HHB ;
wire  hhc ;
wire  HHC ;
wire  hhd ;
wire  HHD ;
wire  hhe ;
wire  HHE ;
wire  hhf ;
wire  HHF ;
wire  hhg ;
wire  HHG ;
wire  hhh ;
wire  HHH ;
wire  hhi ;
wire  HHI ;
wire  hhj ;
wire  HHJ ;
wire  hhk ;
wire  HHK ;
wire  hhl ;
wire  HHL ;
wire  hhm ;
wire  HHM ;
wire  hhn ;
wire  HHN ;
wire  hho ;
wire  HHO ;
wire  hhp ;
wire  HHP ;
wire  hia ;
wire  HIA ;
wire  hib ;
wire  HIB ;
wire  hic ;
wire  HIC ;
wire  hid ;
wire  HID ;
wire  hie ;
wire  HIE ;
wire  hif ;
wire  HIF ;
wire  hig ;
wire  HIG ;
wire  hih ;
wire  HIH ;
wire  hii ;
wire  HII ;
wire  hij ;
wire  HIJ ;
wire  hik ;
wire  HIK ;
wire  hil ;
wire  HIL ;
wire  him ;
wire  HIM ;
wire  hin ;
wire  HIN ;
wire  hio ;
wire  HIO ;
wire  hip ;
wire  HIP ;
wire  hja ;
wire  HJA ;
wire  hjb ;
wire  HJB ;
wire  hjc ;
wire  HJC ;
wire  hjd ;
wire  HJD ;
wire  hje ;
wire  HJE ;
wire  hjf ;
wire  HJF ;
wire  hjg ;
wire  HJG ;
wire  hjh ;
wire  HJH ;
wire  hji ;
wire  HJI ;
wire  hjj ;
wire  HJJ ;
wire  hjk ;
wire  HJK ;
wire  hjl ;
wire  HJL ;
wire  hjm ;
wire  HJM ;
wire  hjn ;
wire  HJN ;
wire  hjo ;
wire  HJO ;
wire  hjp ;
wire  HJP ;
wire  hka ;
wire  HKA ;
wire  hkb ;
wire  HKB ;
wire  hkc ;
wire  HKC ;
wire  hkd ;
wire  HKD ;
wire  hke ;
wire  HKE ;
wire  hkf ;
wire  HKF ;
wire  hkg ;
wire  HKG ;
wire  hkh ;
wire  HKH ;
wire  hki ;
wire  HKI ;
wire  hkj ;
wire  HKJ ;
wire  hkk ;
wire  HKK ;
wire  hkl ;
wire  HKL ;
wire  hkm ;
wire  HKM ;
wire  hkn ;
wire  HKN ;
wire  hko ;
wire  HKO ;
wire  hkp ;
wire  HKP ;
wire  hla ;
wire  HLA ;
wire  hlb ;
wire  HLB ;
wire  hlc ;
wire  HLC ;
wire  hld ;
wire  HLD ;
wire  hle ;
wire  HLE ;
wire  hlf ;
wire  HLF ;
wire  hlg ;
wire  HLG ;
wire  hlh ;
wire  HLH ;
wire  hli ;
wire  HLI ;
wire  hlj ;
wire  HLJ ;
wire  hlk ;
wire  HLK ;
wire  hll ;
wire  HLL ;
wire  hlm ;
wire  HLM ;
wire  hln ;
wire  HLN ;
wire  hlo ;
wire  HLO ;
wire  hlp ;
wire  HLP ;
wire  hma ;
wire  HMA ;
wire  hmb ;
wire  HMB ;
wire  hmc ;
wire  HMC ;
wire  hmd ;
wire  HMD ;
wire  hme ;
wire  HME ;
wire  hmf ;
wire  HMF ;
wire  hmg ;
wire  HMG ;
wire  hmh ;
wire  HMH ;
wire  hmi ;
wire  HMI ;
wire  hmj ;
wire  HMJ ;
wire  hmk ;
wire  HMK ;
wire  hml ;
wire  HML ;
wire  hmm ;
wire  HMM ;
wire  hmn ;
wire  HMN ;
wire  hmo ;
wire  HMO ;
wire  hmp ;
wire  HMP ;
wire  hna ;
wire  HNA ;
wire  hnb ;
wire  HNB ;
wire  hnc ;
wire  HNC ;
wire  hnd ;
wire  HND ;
wire  hne ;
wire  HNE ;
wire  hnf ;
wire  HNF ;
wire  hng ;
wire  HNG ;
wire  hnh ;
wire  HNH ;
wire  hni ;
wire  HNI ;
wire  hnj ;
wire  HNJ ;
wire  hnk ;
wire  HNK ;
wire  hnl ;
wire  HNL ;
wire  hnm ;
wire  HNM ;
wire  hnn ;
wire  HNN ;
wire  hno ;
wire  HNO ;
wire  hnp ;
wire  HNP ;
wire  hoa ;
wire  HOA ;
wire  hob ;
wire  HOB ;
wire  hoc ;
wire  HOC ;
wire  hod ;
wire  HOD ;
wire  hoe ;
wire  HOE ;
wire  hof ;
wire  HOF ;
wire  hog ;
wire  HOG ;
wire  hoh ;
wire  HOH ;
wire  hoi ;
wire  HOI ;
wire  hoj ;
wire  HOJ ;
wire  hok ;
wire  HOK ;
wire  hol ;
wire  HOL ;
wire  hom ;
wire  HOM ;
wire  hon ;
wire  HON ;
wire  hoo ;
wire  HOO ;
wire  hop ;
wire  HOP ;
wire  hpa ;
wire  HPA ;
wire  hpb ;
wire  HPB ;
wire  hpc ;
wire  HPC ;
wire  hpd ;
wire  HPD ;
wire  hpe ;
wire  HPE ;
wire  hpf ;
wire  HPF ;
wire  hpg ;
wire  HPG ;
wire  hph ;
wire  HPH ;
wire  hpi ;
wire  HPI ;
wire  hpj ;
wire  HPJ ;
wire  hpk ;
wire  HPK ;
wire  hpl ;
wire  HPL ;
wire  hpm ;
wire  HPM ;
wire  hpn ;
wire  HPN ;
wire  hpo ;
wire  HPO ;
wire  hpp ;
wire  HPP ;
wire  hqa ;
wire  HQA ;
wire  hqb ;
wire  HQB ;
wire  hqc ;
wire  HQC ;
wire  hqd ;
wire  HQD ;
wire  hqe ;
wire  HQE ;
wire  hqf ;
wire  HQF ;
wire  hqg ;
wire  HQG ;
wire  hqh ;
wire  HQH ;
wire  hqi ;
wire  HQI ;
wire  hqj ;
wire  HQJ ;
wire  hqk ;
wire  HQK ;
wire  hql ;
wire  HQL ;
wire  hqm ;
wire  HQM ;
wire  hqn ;
wire  HQN ;
wire  hqo ;
wire  HQO ;
wire  hqp ;
wire  HQP ;
wire  hra ;
wire  HRA ;
wire  hrb ;
wire  HRB ;
wire  hrc ;
wire  HRC ;
wire  hrd ;
wire  HRD ;
wire  hre ;
wire  HRE ;
wire  hrf ;
wire  HRF ;
wire  hrg ;
wire  HRG ;
wire  hrh ;
wire  HRH ;
wire  hri ;
wire  HRI ;
wire  hrj ;
wire  HRJ ;
wire  hrk ;
wire  HRK ;
wire  hrl ;
wire  HRL ;
wire  hrm ;
wire  HRM ;
wire  hrn ;
wire  HRN ;
wire  hro ;
wire  HRO ;
wire  hrp ;
wire  HRP ;
wire  hsa ;
wire  HSA ;
wire  hsb ;
wire  HSB ;
wire  hsc ;
wire  HSC ;
wire  hsd ;
wire  HSD ;
wire  hse ;
wire  HSE ;
wire  hsf ;
wire  HSF ;
wire  hsg ;
wire  HSG ;
wire  hsh ;
wire  HSH ;
wire  hsi ;
wire  HSI ;
wire  hsj ;
wire  HSJ ;
wire  hsk ;
wire  HSK ;
wire  hsl ;
wire  HSL ;
wire  hsm ;
wire  HSM ;
wire  hsn ;
wire  HSN ;
wire  hso ;
wire  HSO ;
wire  hsp ;
wire  HSP ;
wire  hta ;
wire  HTA ;
wire  htb ;
wire  HTB ;
wire  htc ;
wire  HTC ;
wire  htd ;
wire  HTD ;
wire  hte ;
wire  HTE ;
wire  htf ;
wire  HTF ;
wire  htg ;
wire  HTG ;
wire  hth ;
wire  HTH ;
wire  hti ;
wire  HTI ;
wire  htj ;
wire  HTJ ;
wire  htk ;
wire  HTK ;
wire  htl ;
wire  HTL ;
wire  htm ;
wire  HTM ;
wire  htn ;
wire  HTN ;
wire  hto ;
wire  HTO ;
wire  htp ;
wire  HTP ;
wire  iaa ;
wire  iab ;
wire  iac ;
wire  iad ;
wire  iae ;
wire  iaf ;
wire  iag ;
wire  iah ;
wire  iba ;
wire  ibb ;
wire  ibc ;
wire  ibd ;
wire  ibe ;
wire  ibf ;
wire  ibg ;
wire  ibh ;
wire  ica ;
wire  icb ;
wire  icc ;
wire  icd ;
wire  ice ;
wire  icf ;
wire  icg ;
wire  ich ;
wire  ida ;
wire  idb ;
wire  idc ;
wire  idd ;
wire  ide ;
wire  idf ;
wire  idg ;
wire  idh ;
wire  iea ;
wire  ieb ;
wire  iec ;
wire  ied ;
wire  iee ;
wire  ief ;
wire  ieg ;
wire  ieh ;
wire  ifa ;
wire  ifb ;
wire  ifc ;
wire  ifd ;
wire  ife ;
wire  ifff  ;
wire  ifg ;
wire  ifh ;
wire  iga ;
wire  igb ;
wire  igc ;
wire  igd ;
wire  ige ;
wire  igf ;
wire  igg ;
wire  igh ;
wire  iha ;
wire  ihb ;
wire  ihc ;
wire  ihd ;
wire  ihe ;
wire  ihf ;
wire  ihg ;
wire  ihh ;
wire  iia ;
wire  iib ;
wire  iic ;
wire  iid ;
wire  iie ;
wire  iif ;
wire  iig ;
wire  iih ;
wire  ija ;
wire  ijb ;
wire  ijc ;
wire  ijd ;
wire  ije ;
wire  ijf ;
wire  ijg ;
wire  ijh ;
wire  ika ;
wire  ikb ;
wire  ikc ;
wire  ikd ;
wire  ike ;
wire  ikf ;
wire  ikg ;
wire  ikh ;
wire  ima ;
wire  imb ;
wire  imc ;
wire  imd ;
wire  ime ;
wire  imf ;
wire  img ;
wire  imh ;
wire  ina ;
wire  inb ;
wire  inc ;
wire  ind ;
wire  ine ;
wire  inf ;
wire  ing ;
wire  inh ;
wire  ioa ;
wire  iob ;
wire  ioc ;
wire  iod ;
wire  ioe ;
wire  iof ;
wire  iog ;
wire  ioh ;
wire  ipa ;
wire  ipb ;
wire  ipc ;
wire  ipd ;
wire  ipe ;
wire  ipf ;
wire  ipg ;
wire  iph ;
wire  iqa ;
wire  iqb ;
wire  iqc ;
wire  iqd ;
wire  iqe ;
wire  iqf ;
wire  iqg ;
wire  iqh ;
wire  ira ;
wire  irb ;
wire  irc ;
wire  ird ;
wire  ire ;
wire  irf ;
wire  irg ;
wire  irh ;
wire  isa ;
wire  isb ;
wire  isc ;
wire  isd ;
wire  ise ;
wire  isf ;
wire  isg ;
wire  ita ;
wire  itb ;
wire  itc ;
wire  itd ;
wire  ite ;
wire  itf ;
wire  jaa ;
wire  JAA ;
wire  jab ;
wire  JAB ;
wire  jac ;
wire  JAC ;
wire  jad ;
wire  JAD ;
wire  jae ;
wire  JAE ;
wire  jaf ;
wire  JAF ;
wire  jag ;
wire  JAG ;
wire  jah ;
wire  JAH ;
wire  jai ;
wire  JAI ;
wire  jaj ;
wire  JAJ ;
wire  jak ;
wire  JAK ;
wire  jal ;
wire  JAL ;
wire  jam ;
wire  JAM ;
wire  jan ;
wire  JAN ;
wire  jao ;
wire  JAO ;
wire  jap ;
wire  JAP ;
wire  jba ;
wire  JBA ;
wire  jbb ;
wire  JBB ;
wire  jbc ;
wire  JBC ;
wire  jbd ;
wire  JBD ;
wire  jbe ;
wire  JBE ;
wire  jbf ;
wire  JBF ;
wire  jbg ;
wire  JBG ;
wire  jbh ;
wire  JBH ;
wire  jbi ;
wire  JBI ;
wire  jbj ;
wire  JBJ ;
wire  jbk ;
wire  JBK ;
wire  jbl ;
wire  JBL ;
wire  jbm ;
wire  JBM ;
wire  jbn ;
wire  JBN ;
wire  jbo ;
wire  JBO ;
wire  jbp ;
wire  JBP ;
wire  jea ;
wire  JEA ;
wire  jeb ;
wire  JEB ;
wire  jec ;
wire  JEC ;
wire  jed ;
wire  JED ;
wire  jee ;
wire  JEE ;
wire  jef ;
wire  JEF ;
wire  jeg ;
wire  JEG ;
wire  jeh ;
wire  JEH ;
wire  KAA ;
wire  KAB ;
wire  KAC ;
wire  KAD ;
wire  KAE ;
wire  KAF ;
wire  KAG ;
wire  KAH ;
wire  KBA ;
wire  KBB ;
wire  KBC ;
wire  KBD ;
wire  KBE ;
wire  KBF ;
wire  KBG ;
wire  KBH ;
wire  KCA ;
wire  KCB ;
wire  KCC ;
wire  KCD ;
wire  KCE ;
wire  KCF ;
wire  KCG ;
wire  KCH ;
wire  KDA ;
wire  KDB ;
wire  KDC ;
wire  KDD ;
wire  KDE ;
wire  KDF ;
wire  KDG ;
wire  KDH ;
wire  KEA ;
wire  KEB ;
wire  KEC ;
wire  KED ;
wire  KEE ;
wire  KEF ;
wire  KEG ;
wire  KEH ;
wire  KFA ;
wire  KFB ;
wire  KFC ;
wire  KFD ;
wire  KFE ;
wire  KFF ;
wire  KFG ;
wire  KFH ;
wire  laa ;
wire  lab ;
wire  lac ;
wire  lba ;
wire  lbb ;
wire  lbc ;
wire  lca ;
wire  lcb ;
wire  lcc ;
wire  lda ;
wire  ldb ;
wire  ldc ;
wire  lea ;
wire  leb ;
wire  lec ;
wire  lfa ;
wire  lfb ;
wire  lfc ;
wire  lga ;
wire  lgb ;
wire  lgc ;
wire  lha ;
wire  lhb ;
wire  lhc ;
wire  lia ;
wire  lib ;
wire  lic ;
wire  lja ;
wire  ljb ;
wire  ljc ;
wire  lka ;
wire  lkb ;
wire  lkc ;
wire  lla ;
wire  llb ;
wire  llc ;
wire  lma ;
wire  lmb ;
wire  lmc ;
wire  lna ;
wire  lnb ;
wire  lnc ;
wire  loa ;
wire  lob ;
wire  loc ;
wire  lpa ;
wire  lpb ;
wire  lpc ;
wire  lqa ;
wire  lqb ;
wire  lqc ;
wire  lra ;
wire  lrb ;
wire  lrc ;
wire  lsa ;
wire  lsb ;
wire  lsc ;
wire  lta ;
wire  ltb ;
wire  ltc ;
wire  maa ;
wire  MAA ;
wire  mab ;
wire  MAB ;
wire  mac ;
wire  MAC ;
wire  mad ;
wire  MAD ;
wire  mae ;
wire  MAE ;
wire  maf ;
wire  MAF ;
wire  mag ;
wire  MAG ;
wire  mah ;
wire  MAH ;
wire  naa ;
wire  nab ;
wire  nac ;
wire  nad ;
wire  nba ;
wire  nbb ;
wire  nbc ;
wire  nbd ;
wire  nca ;
wire  ncb ;
wire  ncc ;
wire  ncd ;
wire  nda ;
wire  ndb ;
wire  ndc ;
wire  ndd ;
wire  nea ;
wire  neb ;
wire  nec ;
wire  ned ;
wire  nfa ;
wire  nfb ;
wire  nfc ;
wire  nfd ;
wire  nga ;
wire  ngb ;
wire  ngc ;
wire  ngd ;
wire  nha ;
wire  nhb ;
wire  nhc ;
wire  nhd ;
wire  OAA ;
wire  OAB ;
wire  OAC ;
wire  OAD ;
wire  OAE ;
wire  OAF ;
wire  OAG ;
wire  OAH ;
wire  OBA ;
wire  OBB ;
wire  OBC ;
wire  OBD ;
wire  OBE ;
wire  OBF ;
wire  OBG ;
wire  OBH ;
wire  OCA ;
wire  OCB ;
wire  OCC ;
wire  OCD ;
wire  OCE ;
wire  OCF ;
wire  OCG ;
wire  OCH ;
wire  oda ;
wire  odb ;
wire  odc ;
wire  odd ;
wire  ode ;
wire  odf ;
wire  odg ;
wire  odh ;
wire  oea ;
wire  oeb ;
wire  oec ;
wire  oed ;
wire  oee ;
wire  oef ;
wire  oeg ;
wire  oeh ;
wire  ofa ;
wire  ofb ;
wire  ofc ;
wire  ofd ;
wire  ofe ;
wire  off ;
wire  ofg ;
wire  ofh ;
wire  oga ;
wire  ogb ;
wire  ogc ;
wire  ogd ;
wire  oge ;
wire  ogf ;
wire  ogg ;
wire  ogh ;
wire  oha ;
wire  ohb ;
wire  ohc ;
wire  ohd ;
wire  ohe ;
wire  ohf ;
wire  ohg ;
wire  ohh ;
wire  oia ;
wire  oib ;
wire  oic ;
wire  oid ;
wire  oie ;
wire  oif ;
wire  oig ;
wire  oih ;
wire  oja ;
wire  ojb ;
wire  ojc ;
wire  ojd ;
wire  oje ;
wire  ojf ;
wire  ojg ;
wire  ojh ;
wire  oka ;
wire  okb ;
wire  okc ;
wire  okd ;
wire  oke ;
wire  okf ;
wire  okg ;
wire  okh ;
wire  ola ;
wire  olb ;
wire  olc ;
wire  old ;
wire  ole ;
wire  olf ;
wire  olg ;
wire  olh ;
wire  oma ;
wire  omb ;
wire  omc ;
wire  omd ;
wire  ome ;
wire  omf ;
wire  omg ;
wire  omh ;
wire  ona ;
wire  onb ;
wire  onc ;
wire  ond ;
wire  one ;
wire  onf ;
wire  ong ;
wire  onh ;
wire  ooa ;
wire  oob ;
wire  ooc ;
wire  ood ;
wire  ooe ;
wire  oof ;
wire  oog ;
wire  ooh ;
wire  OQA ;
wire  oqb ;
wire  ora ;
wire  qaa ;
wire  qab ;
wire  qac ;
wire  qba ;
wire  QCA ;
wire  QCB ;
wire  QCC ;
wire  qda ;
wire  qdb ;
wire  qdc ;
wire  qea ;
wire  qeb ;
wire  qec ;

   wire RAA;
   wire RAB;
   wire RAC;
   wire RAD;
   wire RAE;
   wire RAF;
   wire RAG;
   wire RAH;
   wire RAI;
   wire RAJ;
   wire RAK;
   wire RAL;
   wire RAM;
   wire RAN;
   wire RAO;
   wire RAP;
   wire RBA;
   wire RBB;
   wire RBC;
   wire RBD;
   wire RBE;
   wire RBF;
   wire RBG;
   wire RBH;
   wire RBI;
   wire RBJ;
   wire RBK;
   wire RBL;
   wire RBM;
   wire RBN;
   wire RBO;
   wire RBP;

   wire RCA;
   wire RCB;
   wire RCC;
   wire RCD;
   wire RCE;
   wire RCF;
   wire RCG;
   wire RCH;
   wire RCI;
   wire RCJ;
   wire RCK;
   wire RCL;
   wire RCM;
   wire RCN;
   wire RCO;
   wire RCP;
   wire RDA;
   wire RDB;
   wire RDC;
   wire RDD;
   wire RDE;
   wire RDF;
   wire RDG;
   wire RDH;
   wire RDI;
   wire RDJ;
   wire RDK;
   wire RDL;
   wire RDM;
   wire RDN;
   wire RDO;
   wire RDP;

   wire REA;
   wire REB;
   wire REC;
   wire RED;
   wire REE;
   wire REFF;
   wire REG;
   wire REH;
   wire REI;
   wire REJ;
   wire REK;
   wire REL;
   wire REM;
   wire REN;
   wire REO;
   wire REP;
   wire RFA;
   wire RFB;
   wire RFC;
   wire RFD;
   wire RFE;
   wire RFF;
   wire RFG;
   wire RFH;
   wire RFI;
   wire RFJ;
   wire RFK;
   wire RFL;
   wire RFM;
   wire RFN;
   wire RFO;
   wire RFP;

   wire RGA;
   wire RGB;
   wire RGC;
   wire RGD;
   wire RGE;
   wire RGF;
   wire RGG;
   wire RGH;
   wire RGI;
   wire RGJ;
   wire RGK;
   wire RGL;
   wire RGM;
   wire RGN;
   wire RGO;
   wire RGP;
   wire RHA;
   wire RHB;
   wire RHC;
   wire RHD;
   wire RHE;
   wire RHF;
   wire RHG;
   wire RHH;
   wire RHI;
   wire RHJ;
   wire RHK;
   wire RHL;
   wire RHM;
   wire RHN;
   wire RHO;
   wire RHP;

   wire RIA;
   wire RIB;
   wire RIC;
   wire RID;
   wire RIE;
   wire RIF;
   wire RIG;
   wire RIH;
   wire RII;
   wire RIJ;
   wire RIK;
   wire RIL;
   wire RIM;
   wire RIN;
   wire RIO;
   wire RIP;
   wire RJA;
   wire RJB;
   wire RJC;
   wire RJD;
   wire RJE;
   wire RJF;
   wire RJG;
   wire RJH;
   wire RJI;
   wire RJJ;
   wire RJK;
   wire RJL;
   wire RJM;
   wire RJN;
   wire RJO;
   wire RJP;

   wire RKA;
   wire RKB;
   wire RKC;
   wire RKD;
   wire RKE;
   wire RKF;
   wire RKG;
   wire RKH;
   wire RKI;
   wire RKJ;
   wire RKK;
   wire RKL;
   wire RKM;
   wire RKN;
   wire RKO;
   wire RKP;
   wire RLA;
   wire RLB;
   wire RLC;
   wire RLD;
   wire RLE;
   wire RLF;
   wire RLG;
   wire RLH;
   wire RLI;
   wire RLJ;
   wire RLK;
   wire RLL;
   wire RLM;
   wire RLN;
   wire RLO;
   wire RLP;

   wire RMA;
   wire RMB;
   wire RMC;
   wire RMD;
   wire RME;
   wire RMF;
   wire RMG;
   wire RMH;
   wire RMI;
   wire RMJ;
   wire RMK;
   wire RML;
   wire RMM;
   wire RMN;
   wire RMO;
   wire RMP;
   wire RNA;
   wire RNB;
   wire RNC;
   wire RND;
   wire RNE;
   wire RNF;
   wire RNG;
   wire RNH;
   wire RNI;
   wire RNJ;
   wire RNK;
   wire RNL;
   wire RNM;
   wire RNN;
   wire RNO;
   wire RNP;

   wire ROA;
   wire ROB;
   wire ROC;
   wire ROD;
   wire ROE;
   wire ROF;
   wire ROG;
   wire ROH;
   wire ROI;
   wire ROJ;
   wire ROK;
   wire ROL;
   wire ROM;
   wire RON;
   wire ROO;
   wire ROP;
   wire RPA;
   wire RPB;
   wire RPC;
   wire RPD;
   wire RPE;
   wire RPF;
   wire RPG;
   wire RPH;
   wire RPI;
   wire RPJ;
   wire RPK;
   wire RPL;
   wire RPM;
   wire RPN;
   wire RPO;
   wire RPP;
   
wire  saa ;
wire  sab ;
wire  sac ;
wire  sad ;
wire  sae ;
wire  saf ;
wire  sag ;
wire  sah ;
wire  sba ;
wire  sbb ;
wire  sbc ;
wire  sbd ;
wire  sbe ;
wire  sbf ;
wire  sbg ;
wire  sbh ;
wire  sca ;
wire  scb ;
wire  scc ;
wire  scd ;
wire  sce ;
wire  scf ;
wire  scg ;
wire  sch ;
wire  sda ;
wire  sdb ;
wire  sdc ;
wire  sdd ;
wire  sde ;
wire  sdf ;
wire  sdg ;
wire  sdh ;
wire  sea ;
wire  seb ;
wire  sec ;
wire  sed ;
wire  see ;
wire  sef ;
wire  seg ;
wire  seh ;
wire  sfa ;
wire  sfb ;
wire  sfc ;
wire  sfd ;
wire  sfe ;
wire  sff ;
wire  sfg ;
wire  sfh ;
wire  sga ;
wire  sgb ;
wire  sgc ;
wire  sgd ;
wire  sge ;
wire  sgf ;
wire  sgg ;
wire  sgh ;
wire  sha ;
wire  shb ;
wire  shc ;
wire  shd ;
wire  she ;
wire  shf ;
wire  shg ;
wire  shh ;
wire  sja ;
wire  sjb ;
wire  sjc ;
wire  sjd ;
wire  sje ;
wire  sjf ;
wire  sjg ;
wire  sjh ;
wire  SKA ;
wire  SKB ;
wire  SKC ;
wire  SKD ;
wire  SKE ;
wire  SKF ;
wire  SKG ;
wire  SKH ;
wire  taa ;
wire  tab ;
wire  tac ;
wire  tad ;
wire  tba ;
wire  tbb ;
wire  tbc ;
wire  tbd ;
wire  tca ;
wire  tcb ;
wire  tcc ;
wire  tcd ;
wire  tda ;
wire  tdb ;
wire  tdc ;
wire  tdd ;
wire  tea ;
wire  teb ;
wire  tec ;
wire  ted ;
wire  tfa ;
wire  tfb ;
wire  tfc ;
wire  tfd ;
wire  tga ;
wire  tgb ;
wire  tgc ;
wire  tgd ;
wire  tha ;
wire  thb ;
wire  thc ;
wire  thd ;
wire  tib ;
wire  tic ;
wire  tid ;
wire  tie ;
wire  tif ;
wire  tig ;
wire  tjb ;
wire  tjc ;
wire  tjd ;
wire  tje ;
wire  tjf ;
wire  tjg ;
wire  tkb ;
wire  tkc ;
wire  tkd ;
wire  tke ;
wire  tkf ;
wire  tkg ;
wire  tsa ;
wire  tsb ;
wire  tsc ;
wire  tsd ;
wire  tse ;
wire  tsf ;
wire  tsg ;
wire  tsh ;
wire  uaa ;
wire  uab ;
wire  uac ;
wire  uad ;
wire  uae ;
wire  uaf ;
wire  uag ;
wire  uah ;
wire  uai ;
wire  uaj ;
wire  uak ;
wire  ual ;
wire  uam ;
wire  uan ;
wire  uao ;
wire  uap ;
wire  uaq ;
wire  uar ;
wire  uas ;
wire  uat ;
wire  uau ;
wire  uav ;
wire  uaw ;
wire  uax ;
wire  uba ;
wire  ubb ;
wire  ubc ;
wire  ubd ;
wire  ube ;
wire  ubf ;
wire  ubg ;
wire  ubh ;
wire  ubi ;
wire  ubj ;
wire  ubk ;
wire  ubl ;
wire  ubm ;
wire  ubn ;
wire  ubo ;
wire  ubp ;
wire  ubq ;
wire  ubr ;
wire  ubs ;
wire  ubt ;
wire  ubu ;
wire  ubv ;
wire  ubw ;
wire  ubx ;
wire  uca ;
wire  ucb ;
wire  ucc ;
wire  ucd ;
wire  uce ;
wire  ucf ;
wire  ucg ;
wire  uch ;
wire  uci ;
wire  ucj ;
wire  uck ;
wire  ucl ;
wire  ucm ;
wire  ucn ;
wire  uco ;
wire  ucp ;
wire  ucq ;
wire  ucr ;
wire  ucs ;
wire  uct ;
wire  ucu ;
wire  ucv ;
wire  ucw ;
wire  ucx ;
wire  uda ;
wire  udb ;
wire  udc ;
wire  udd ;
wire  ude ;
wire  udf ;
wire  udg ;
wire  udh ;
wire  udi ;
wire  udj ;
wire  udk ;
wire  udl ;
wire  udm ;
wire  udn ;
wire  udo ;
wire  udp ;
wire  udq ;
wire  udr ;
wire  uds ;
wire  udt ;
wire  udu ;
wire  udv ;
wire  udw ;
wire  udx ;
wire  uea ;
wire  ueb ;
wire  uec ;
wire  ued ;
wire  uee ;
wire  uef ;
wire  ueg ;
wire  ueh ;
wire  uei ;
wire  uej ;
wire  uek ;
wire  uel ;
wire  uem ;
wire  uen ;
wire  ueo ;
wire  uep ;
wire  ueq ;
wire  uer ;
wire  ues ;
wire  uet ;
wire  ueu ;
wire  uev ;
wire  uew ;
wire  uex ;
wire  ufa ;
wire  ufb ;
wire  ufc ;
wire  ufd ;
wire  ufe ;
wire  uff ;
wire  ufg ;
wire  ufh ;
wire  ufi ;
wire  ufj ;
wire  ufk ;
wire  ufl ;
wire  ufm ;
wire  ufn ;
wire  ufo ;
wire  ufp ;
wire  ufq ;
wire  ufr ;
wire  ufs ;
wire  uft ;
wire  ufu ;
wire  ufv ;
wire  ufw ;
wire  ufx ;
wire  uga ;
wire  ugb ;
wire  ugc ;
wire  ugd ;
wire  uge ;
wire  ugf ;
wire  ugg ;
wire  ugh ;
wire  ugi ;
wire  ugj ;
wire  ugk ;
wire  ugl ;
wire  ugm ;
wire  ugn ;
wire  ugo ;
wire  ugp ;
wire  ugq ;
wire  ugr ;
wire  ugs ;
wire  ugt ;
wire  ugu ;
wire  ugv ;
wire  ugw ;
wire  ugx ;
wire  uha ;
wire  uhb ;
wire  uhc ;
wire  uhd ;
wire  uhe ;
wire  uhf ;
wire  uhg ;
wire  uhh ;
wire  uhi ;
wire  uhj ;
wire  uhk ;
wire  uhl ;
wire  uhm ;
wire  uhn ;
wire  uho ;
wire  uhp ;
wire  uhq ;
wire  uhr ;
wire  uhs ;
wire  uht ;
wire  uhu ;
wire  uhv ;
wire  uhw ;
wire  uhx ;
wire  vaa ;
wire  vab ;
wire  vac ;
wire  vad ;
wire  vae ;
wire  vaf ;
wire  vag ;
wire  vah ;
wire  vai ;
wire  vaj ;
wire  vak ;
wire  val ;
wire  vam ;
wire  van ;
wire  vao ;
wire  vap ;
wire  vba ;
wire  vbb ;
wire  vbc ;
wire  vbd ;
wire  vbe ;
wire  vbf ;
wire  vbg ;
wire  vbh ;
wire  vbi ;
wire  vbj ;
wire  vbk ;
wire  vbl ;
wire  vbm ;
wire  vbn ;
wire  vbo ;
wire  vbp ;
wire  vca ;
wire  vcb ;
wire  vcc ;
wire  vcd ;
wire  vce ;
wire  vcf ;
wire  vcg ;
wire  vch ;
wire  vci ;
wire  vcj ;
wire  vck ;
wire  vcl ;
wire  vcm ;
wire  vcn ;
wire  vco ;
wire  vcp ;
wire  vda ;
wire  vdb ;
wire  vdc ;
wire  vdd ;
wire  vde ;
wire  vdf ;
wire  vdg ;
wire  vdh ;
wire  vdi ;
wire  vdj ;
wire  vdk ;
wire  vdl ;
wire  vdm ;
wire  vdn ;
wire  vdo ;
wire  vdp ;
wire  vea ;
wire  veb ;
wire  vec ;
wire  ved ;
wire  vee ;
wire  vef ;
wire  veg ;
wire  veh ;
wire  vei ;
wire  vej ;
wire  vek ;
wire  vel ;
wire  vem ;
wire  ven ;
wire  veo ;
wire  vep ;
wire  vfa ;
wire  vfb ;
wire  vfc ;
wire  vfd ;
wire  vfe ;
wire  vff ;
wire  vfg ;
wire  vfh ;
wire  vfi ;
wire  vfj ;
wire  vfk ;
wire  vfl ;
wire  vfm ;
wire  vfn ;
wire  vfo ;
wire  vfp ;
wire  vga ;
wire  vgb ;
wire  vgc ;
wire  vgd ;
wire  vge ;
wire  vgf ;
wire  vgg ;
wire  vgh ;
wire  vgi ;
wire  vgj ;
wire  vgk ;
wire  vgl ;
wire  vgm ;
wire  vgn ;
wire  vgo ;
wire  vgp ;
wire  vha ;
wire  vhb ;
wire  vhc ;
wire  vhd ;
wire  vhe ;
wire  vhf ;
wire  vhg ;
wire  vhh ;
wire  vhi ;
wire  vhj ;
wire  vhk ;
wire  vhl ;
wire  vhm ;
wire  vhn ;
wire  vho ;
wire  vhp ;
wire  waa ;
wire  wab ;
wire  wac ;
wire  wad ;
wire  wae ;
wire  waf ;
wire  wag ;
wire  wah ;
wire  wba ;
wire  wbb ;
wire  wbc ;
wire  wbd ;
wire  wbe ;
wire  wbf ;
wire  wbg ;
wire  wbh ;
wire  wca ;
wire  wcb ;
wire  wcc ;
wire  wcd ;
wire  wce ;
wire  wcf ;
wire  wcg ;
wire  wch ;
wire  wda ;
wire  wdb ;
wire  wdc ;
wire  wdd ;
wire  wde ;
wire  wdf ;
wire  wdg ;
wire  wdh ;
wire  wea ;
wire  web ;
wire  wec ;
wire  wed ;
wire  wee ;
wire  wef ;
wire  weg ;
wire  weh ;
wire  wfa ;
wire  wfb ;
wire  wfc ;
wire  wfd ;
wire  wfe ;
wire  wff ;
wire  wfg ;
wire  wfh ;
wire  wga ;
wire  wgb ;
wire  wgc ;
wire  wgd ;
wire  wge ;
wire  wgf ;
wire  wgg ;
wire  wgh ;
wire  wha ;
wire  whb ;
wire  whc ;
wire  whd ;
wire  whe ;
wire  whf ;
wire  whg ;
wire  whh ;
wire  ZZI ;
wire  ZZO ;
assign ZZI = 1'b1;
assign ZZO = 1'b0;
assign uaa = ~UAA;  //complement 
assign uab = ~UAB;  //complement 
assign uac = ~UAC;  //complement 
assign vaa = ~VAA;  //complement 
assign vai = ~VAI;  //complement 
assign hia = vaa & ~lib & ~lia & lic |  vba & ~lib & lia & lic |  vca & lib & ~lia & lic |  vda & lib & lia & lic; 
assign HIA = ~hia;  //complement 
assign hoa = vaa & ~lob & ~loa & loc |         vba & ~lob & loa & loc |  vca & lob & ~loa & loc |  vda & lob & loa & loc; 
assign HOA = ~hoa;  //complement 
assign uad = ~UAD;  //complement 
assign uae = ~UAE;  //complement 
assign uaf = ~UAF;  //complement 
assign vab = ~VAB;  //complement 
assign vaj = ~VAJ;  //complement 
assign hib = vab & ~lib & ~lia & lic |  vbb & ~lib & lia & lic |  vcb & lib & ~lia & lic |  vdb & lib & lia & lic; 
assign HIB = ~hib;  //complement 
assign hob = vab & ~lob & ~loa & loc |         vbb & ~lob & loa & loc |  vcb & lob & ~loa & loc |  vdb & lob & loa & loc; 
assign HOB = ~hob;  //complement 
assign uag = ~UAG;  //complement 
assign uah = ~UAH;  //complement 
assign uai = ~UAI;  //complement 
assign vac = ~VAC;  //complement 
assign vak = ~VAK;  //complement 
assign hic = vac & ~lib & ~lia & lic |  vbc & ~lib & lia & lic |  vcc & lib & ~lia & lic |  vdc & lib & lia & lic; 
assign HIC = ~hic;  //complement 
assign hoc = vac & ~lob & ~loa & loc |         vbc & ~lob & loa & loc |  vcc & lob & ~loa & loc |  vdc & lob & loa & loc; 
assign HOC = ~hoc;  //complement 
assign uaj = ~UAJ;  //complement 
assign uak = ~UAK;  //complement 
assign ual = ~UAL;  //complement 
assign vad = ~VAD;  //complement 
assign val = ~VAL;  //complement 
assign hid = vad & ~lib & ~lia & lic |  vbd & ~lib & lia & lic |  vcd & lib & ~lia & lic |  vdd & lib & lia & lic; 
assign HID = ~hid;  //complement 
assign hod = vad & ~lob & ~loa & loc |         vbd & ~lob & loa & loc |  vcd & lob & ~loa & loc |  vdd & lob & loa & loc; 
assign HOD = ~hod;  //complement 
assign uam = ~UAM;  //complement 
assign uan = ~UAN;  //complement 
assign uao = ~UAO;  //complement 
assign vae = ~VAE;  //complement 
assign vam = ~VAM;  //complement 
assign hie = vae & ~lib & ~lia & lic |  vbe & ~lib & lia & lic |  vce & lib & ~lia & lic |  vde & lib & lia & lic; 
assign HIE = ~hie;  //complement 
assign hoe = vae & ~lob & ~loa & loc |         vbe & ~lob & loa & loc |  vce & lob & ~loa & loc |  vde & lob & loa & loc; 
assign HOE = ~hoe;  //complement 
assign uap = ~UAP;  //complement 
assign uaq = ~UAQ;  //complement 
assign uar = ~UAR;  //complement 
assign vaf = ~VAF;  //complement 
assign van = ~VAN;  //complement 
assign hif = vaf & ~lib & ~lia & lic |  vbf & ~lib & lia & lic |  vcf & lib & ~lia & lic |  vdf & lib & lia & lic; 
assign HIF = ~hif;  //complement 
assign hof = vaf & ~lob & ~loa & loc |         vbf & ~lob & loa & loc |  vcf & lob & ~loa & loc |  vdf & lob & loa & loc; 
assign HOF = ~hof;  //complement 
assign uat = ~UAT;  //complement 
assign uau = ~UAU;  //complement 
assign uas = ~UAS;  //complement 
assign vag = ~VAG;  //complement 
assign vao = ~VAO;  //complement 
assign hig = vag & ~lib & ~lia & lic |  vbg & ~lib & lia & lic |  vcg & lib & ~lia & lic |  vdg & lib & lia & lic; 
assign HIG = ~hig;  //complement 
assign hog = vag & ~lob & ~loa & loc |         vbg & ~lob & loa & loc |  vcg & lob & ~loa & loc |  vdg & lob & loa & loc; 
assign HOG = ~hog;  //complement 
assign uav = ~UAV;  //complement 
assign uaw = ~UAW;  //complement 
assign uax = ~UAX;  //complement 
assign vah = ~VAH;  //complement 
assign vap = ~VAP;  //complement 
assign hih = vah & ~lib & ~lia & lic |  vbh & ~lib & lia & lic |  vch & lib & ~lia & lic |  vdh & lib & lia & lic; 
assign HIH = ~hih;  //complement 
assign hoh = vah & ~lob & ~loa & loc |         vbh & ~lob & loa & loc |  vch & lob & ~loa & loc |  vdh & lob & loa & loc; 
assign HOH = ~hoh;  //complement 
assign hii = vha & ~LIB & ~LIA & LIC |  vga & ~LIB & LIA & LIC |  vfa & LIB & ~LIA & LIC |  vea & LIB & LIA & LIC; 
assign HII = ~hii;  //complement 
assign hoi = vha & ~LOB & ~LOA & LOC |         vga & ~LOB & LOA & LOC |  vfa & LOB & ~LOA & LOC |  vea & LOB & LOA & LOC; 
assign HOI = ~hoi;  //complement 
assign HAA = ZZO & ~lab & ~laa & lac |  KAA & ~lab & laa & lac |  KBA & lab & ~laa & lac |  KCA & lab & laa & lac; 
assign haa = ~HAA;  //complement 
assign HBA = ZZO & ~lbb & ~lba & lbc |         KAA & ~lbb & lba & lbc |  KBA & lbb & ~lba & lbc |  KCA & lbb & lba & lbc; 
assign hba = ~HBA;  //complement 
assign waa = ~WAA;  //complement 
assign wab = ~WAB;  //complement 
assign hij = vhb & ~LIB & ~LIA & LIC |  vgb & ~LIB & LIA & LIC |  vfb & LIB & ~LIA & LIC |  veb & LIB & LIA & LIC; 
assign HIJ = ~hij;  //complement 
assign hoj = vhb & ~LOB & ~LOA & LOC |         vgb & ~LOB & LOA & LOC |  vfb & LOB & ~LOA & LOC |  veb & LOB & LOA & LOC; 
assign HOJ = ~hoj;  //complement 
assign HAB = ZZO & ~lab & ~laa & lac |  KAB & ~lab & laa & lac |  KBB & lab & ~laa & lac |  KCB & lab & laa & lac; 
assign hab = ~HAB;  //complement 
assign HBB = ZZO & ~lbb & ~lba & lbc |         KAB & ~lbb & lba & lbc |  KBB & lbb & ~lba & lbc |  KCB & lbb & lba & lbc; 
assign hbb = ~HBB;  //complement 
assign dam = ~DAM;  //complement 
assign dan = ~DAN;  //complement 
assign taa = ~TAA;  //complement 
assign tab = ~TAB;  //complement 
assign hik = vhc & ~LIB & ~LIA & LIC |  vgc & ~LIB & LIA & LIC |  vfc & LIB & ~LIA & LIC |  vec & LIB & LIA & LIC; 
assign HIK = ~hik;  //complement 
assign hok = vhc & ~LOB & ~LOA & LOC |         vgc & ~LOB & LOA & LOC |  vfc & LOB & ~LOA & LOC |  vec & LOB & LOA & LOC; 
assign HOK = ~hok;  //complement 
assign HAC = ZZO & ~lab & ~laa & lac |  KAC & ~lab & laa & lac |  KBC & lab & ~laa & lac |  KCC & lab & laa & lac; 
assign hac = ~HAC;  //complement 
assign HBC = ZZO & ~lbb & ~lba & lbc |         KAC & ~lbb & lba & lbc |  KBC & lbb & ~lba & lbc |  KCC & lbb & lba & lbc; 
assign hbc = ~HBC;  //complement 
assign KAA = ~kaa;  //complement 
assign KAB = ~kab;  //complement 
assign KAC = ~kac;  //complement 
assign KAD = ~kad;  //complement 
assign hil = vhd & ~LIB & ~LIA & LIC |  vgd & ~LIB & LIA & LIC |  vfd & LIB & ~LIA & LIC |  ved & LIB & LIA & LIC; 
assign HIL = ~hil;  //complement 
assign hol = vhd & ~LOB & ~LOA & LOC |         vgd & ~LOB & LOA & LOC |  vfd & LOB & ~LOA & LOC |  ved & LOB & LOA & LOC; 
assign HOL = ~hol;  //complement 
assign lia = ~LIA;  //complement 
assign lib = ~LIB;  //complement 
assign lic = ~LIC;  //complement 
assign HAD = ZZO & ~lab & ~laa & lac |  KAD & ~lab & laa & lac |  KBD & lab & ~laa & lac |  KCD & lab & laa & lac; 
assign had = ~HAD;  //complement 
assign HBD = ZZO & ~lbb & ~lba & lbc |         KAD & ~lbb & lba & lbc |  KBD & lbb & ~lba & lbc |  KCD & lbb & lba & lbc; 
assign hbd = ~HBD;  //complement 
assign wac = ~WAC;  //complement 
assign wad = ~WAD;  //complement 
assign hom = vhe & ~LOB & ~LOA & LOC |  vge & ~LOB & LOA & LOC |  vfe & LOB & ~LOA & LOC |  vee & LOB & LOA & LOC; 
assign HOM = ~hom;  //complement 
assign loa = ~LOA;  //complement 
assign lob = ~LOB;  //complement 
assign loc = ~LOC;  //complement 
assign HAE = ZZO & ~lab & ~laa & lac |  KAE & ~lab & laa & lac |  KBE & lab & ~laa & lac |  KCE & lab & laa & lac; 
assign hae = ~HAE;  //complement 
assign HBE = ZZO & ~lbb & ~lba & lbc |         KAE & ~lbb & lba & lbc |  KBE & lbb & ~lba & lbc |  KCE & lbb & lba & lbc; 
assign hbe = ~HBE;  //complement 
assign wae = ~WAE;  //complement 
assign waf = ~WAF;  //complement 
assign hin = vhf & ~LIB & ~LIA & LIC |  vgf & ~LIB & LIA & LIC |  vff & LIB & ~LIA & LIC |  vef & LIB & LIA & LIC; 
assign HIN = ~hin;  //complement 
assign hon = vhf & ~LOB & ~LOA & LOC |         vgf & ~LOB & LOA & LOC |  vff & LOB & ~LOA & LOC |  vef & LOB & LOA & LOC; 
assign HON = ~hon;  //complement 
assign HAF = ZZO & ~lab & ~laa & lac |  KAF & ~lab & laa & lac |  KBF & lab & ~laa & lac |  KCF & lab & laa & lac; 
assign haf = ~HAF;  //complement 
assign HBF = ZZO & ~lbb & ~lba & lbc |         KAF & ~lbb & lba & lbc |  KBF & lbb & ~lba & lbc |  KCF & lbb & lba & lbc; 
assign hbf = ~HBF;  //complement 
assign dao = ~DAO;  //complement 
assign dap = ~DAP;  //complement 
assign tac = ~TAC;  //complement 
assign tad = ~TAD;  //complement 
assign hio = vhg & ~LIB & ~LIA & LIC |  vgg & ~LIB & LIA & LIC |  vfg & LIB & ~LIA & LIC |  veg & LIB & LIA & LIC; 
assign HIO = ~hio;  //complement 
assign hoo = vhg & ~LOB & ~LOA & LOC |         vgg & ~LOB & LOA & LOC |  vfg & LOB & ~LOA & LOC |  veg & LOB & LOA & LOC; 
assign HOO = ~hoo;  //complement 
assign him = vhe & ~LIB & ~LIA & LIC |  vge & ~LIB & LIA & LIC |  vfe & LIB & ~LIA & LIC |  vee & LIB & LIA & LIC; 
assign HIM = ~him;  //complement 
assign HAG = ZZO & ~lab & ~laa & lac |  KAG & ~lab & laa & lac |  KBG & lab & ~laa & lac |  KCG & lab & laa & lac; 
assign hag = ~HAG;  //complement 
assign HBG = ZZO & ~lbb & ~lba & lbc |         KAG & ~lbb & lba & lbc |  KBG & lbb & ~lba & lbc |  KCG & lbb & lba & lbc; 
assign hbg = ~HBG;  //complement 
assign KAE = ~kae;  //complement 
assign KAF = ~kaf;  //complement 
assign KAG = ~kag;  //complement 
assign KAH = ~kah;  //complement 
assign hip = vhh & ~LIB & ~LIA & LIC |  vgh & ~LIB & LIA & LIC |  vfh & LIB & ~LIA & LIC |  veh & LIB & LIA & LIC; 
assign HIP = ~hip;  //complement 
assign hop = vhh & ~LOB & ~LOA & LOC |         vgh & ~LOB & LOA & LOC |  vfh & LOB & ~LOA & LOC |  veh & LOB & LOA & LOC; 
assign HOP = ~hop;  //complement 
assign HAH = ZZO & ~lab & ~laa & lac |  KAH & ~lab & laa & lac |  KBH & lab & ~laa & lac |  KCH & lab & laa & lac; 
assign hah = ~HAH;  //complement 
assign HBH = ZZO & ~lbb & ~lba & lbc |         KAH & ~lbb & lba & lbc |  KBH & lbb & ~lba & lbc |  KCH & lbb & lba & lbc; 
assign hbh = ~HBH;  //complement 
assign wag = ~WAG;  //complement 
assign wah = ~WAH;  //complement 
assign ofa = ~OFA;  //complement 
assign oea = ~OEA;  //complement 
assign DAI = ~dai;  //complement 
assign DAJ = ~daj;  //complement 
assign DAK = ~dak;  //complement 
assign DAL = ~dal;  //complement 
assign ofb = ~OFB;  //complement 
assign oeb = ~OEB;  //complement 
assign saa = ~SAA;  //complement 
assign sab = ~SAB;  //complement 
assign gaa = ~GAA;  //complement 
assign gai = ~GAI;  //complement 
assign ofc = ~OFC;  //complement 
assign oec = ~OEC;  //complement 
assign sba = ~SBA;  //complement 
assign sbb = ~SBB;  //complement 
assign MAA =  SJA & SKA & QDA  |  SJA & ska & QDB  |  sja & SKA & QDC  ; 
assign maa = ~MAA; //complement 
assign ofd = ~OFD;  //complement 
assign oed = ~OED;  //complement 
assign JAA =  SAA & NAA  |  SBA & NBA  |  SCA & NCA  |  SDA & NDA  ; 
assign jaa = ~JAA;  //complement 
assign JAI =  SAA & NAA  |  SBA & NBA  |  SCA & NCA  |  SDA & NDA  ; 
assign jai = ~JAI; //complement 
assign naa = ~NAA;  //complement 
assign nca = ~NCA;  //complement 
assign qda = ~QDA;  //complement 
assign sja = ~SJA;  //complement 
assign ofe = ~OFE;  //complement 
assign oee = ~OEE;  //complement 
assign JAB =  SAB & NAA  |  SBB & NBA  |  SCB & NCA  |  SDB & NDA  ; 
assign jab = ~JAB;  //complement 
assign JAJ =  SAB & NAA  |  SBB & NBA  |  SCB & NCA  |  SDB & NDA  ; 
assign jaj = ~JAJ; //complement 
assign dag = ~DAG;  //complement 
assign nba = ~NBA;  //complement 
assign nda = ~NDA;  //complement 
assign off = ~OFF;  //complement 
assign oef = ~OEF;  //complement 
assign sca = ~SCA;  //complement 
assign scb = ~SCB;  //complement 
assign OAA = ~oaa;  //complement 
assign OBA = ~oba;  //complement 
assign OCA = ~oca;  //complement 
assign SKA = ~ska;  //complement 
assign ofg = ~OFG;  //complement 
assign oeg = ~OEG;  //complement 
assign sda = ~SDA;  //complement 
assign sdb = ~SDB;  //complement 
assign gba = ~GBA;  //complement 
assign gbi = ~GBI;  //complement 
assign ofh = ~OFH;  //complement 
assign oeh = ~OEH;  //complement 
assign laa = ~LAA;  //complement 
assign lab = ~LAB;  //complement 
assign lac = ~LAC;  //complement 
assign dac = ~DAC;  //complement 
assign dad = ~DAD;  //complement 
assign dae = ~DAE;  //complement 
assign daf = ~DAF;  //complement 
assign uba = ~UBA;  //complement 
assign ubb = ~UBB;  //complement 
assign ubc = ~UBC;  //complement 
assign vba = ~VBA;  //complement 
assign vbi = ~VBI;  //complement 
assign hja = vaa & ~ljb & ~lja & ljc |  vba & ~ljb & lja & ljc |  vca & ljb & ~lja & ljc |  vda & ljb & lja & ljc; 
assign HJA = ~hja;  //complement 
assign hpa = vaa & ~lpb & ~lpa & lpc |         vba & ~lpb & lpa & lpc |  vca & lpb & ~lpa & lpc |  vda & lpb & lpa & lpc; 
assign HPA = ~hpa;  //complement 
assign ubd = ~UBD;  //complement 
assign ube = ~UBE;  //complement 
assign ubf = ~UBF;  //complement 
assign vbb = ~VBB;  //complement 
assign vbj = ~VBJ;  //complement 
assign hjb = vab & ~ljb & ~lja & ljc |  vbb & ~ljb & lja & ljc |  vcb & ljb & ~lja & ljc |  vdb & ljb & lja & ljc; 
assign HJB = ~hjb;  //complement 
assign hpb = vab & ~lpb & ~lpa & lpc |         vbb & ~lpb & lpa & lpc |  vcb & lpb & ~lpa & lpc |  vdb & lpb & lpa & lpc; 
assign HPB = ~hpb;  //complement 
assign ubg = ~UBG;  //complement 
assign ubh = ~UBH;  //complement 
assign ubi = ~UBI;  //complement 
assign vbc = ~VBC;  //complement 
assign vbk = ~VBK;  //complement 
assign hjc = vac & ~ljb & ~lja & ljc |  vbc & ~ljb & lja & ljc |  vcc & ljb & ~lja & ljc |  vdc & ljb & lja & ljc; 
assign HJC = ~hjc;  //complement 
assign hpc = vac & ~lpb & ~lpa & lpc |         vbc & ~lpb & lpa & lpc |  vcc & lpb & ~lpa & lpc |  vdc & lpb & lpa & lpc; 
assign HPC = ~hpc;  //complement 
assign ubj = ~UBJ;  //complement 
assign ubk = ~UBK;  //complement 
assign ubl = ~UBL;  //complement 
assign vbd = ~VBD;  //complement 
assign vbl = ~VBL;  //complement 
assign hpe = vae & ~lpb & ~lpa & lpc |  vbe & ~lpb & lpa & lpc |  vce & lpb & ~lpa & lpc |  vde & lpb & lpa & lpc; 
assign HPE = ~hpe;  //complement 
assign hqe = vae & ~lqb & ~lqa & lqc |         vbe & ~lqb & lqa & lqc |  vce & lqb & ~lqa & lqc |  vde & lqb & lqa & lqc; 
assign HQE = ~hqe;  //complement 
assign ubm = ~UBM;  //complement 
assign ubn = ~UBN;  //complement 
assign ubo = ~UBO;  //complement 
assign vbe = ~VBE;  //complement 
assign vbm = ~VBM;  //complement 
assign hpd = vad & ~lpb & ~lpa & lpc |  vbd & ~lpb & lpa & lpc |  vcd & lpb & ~lpa & lpc |  vdd & lpb & lpa & lpc; 
assign HPD = ~hpd;  //complement 
assign hjd = vad & ~ljb & ~lja & ljc |         vbd & ~ljb & lja & ljc |  vcd & ljb & ~lja & ljc |  vdd & ljb & lja & ljc; 
assign HJD = ~hjd;  //complement 
assign ubp = ~UBP;  //complement 
assign ubq = ~UBQ;  //complement 
assign ubr = ~UBR;  //complement 
assign vbn = ~VBN;  //complement 
assign vbf = ~VBF;  //complement 
assign hjf = vaf & ~ljb & ~lja & ljc |  vbf & ~ljb & lja & ljc |  vcf & ljb & ~lja & ljc |  vdf & ljb & lja & ljc; 
assign HJF = ~hjf;  //complement 
assign hpf = vaf & ~lpb & ~lpa & lpc |         vbf & ~lpb & lpa & lpc |  vcf & lpb & ~lpa & lpc |  vdf & lpb & lpa & lpc; 
assign HPF = ~hpf;  //complement 
assign ubs = ~UBS;  //complement 
assign ubt = ~UBT;  //complement 
assign ubu = ~UBU;  //complement 
assign vbg = ~VBG;  //complement 
assign vbo = ~VBO;  //complement 
assign hjg = vag & ~ljb & ~lja & ljc |  vbg & ~ljb & lja & ljc |  vcg & ljb & ~lja & ljc |  vdg & ljb & lja & ljc; 
assign HJG = ~hjg;  //complement 
assign hpg = vag & ~lpb & ~lpa & lpc |         vbg & ~lpb & lpa & lpc |  vcg & lpb & ~lpa & lpc |  vdg & lpb & lpa & lpc; 
assign HPG = ~hpg;  //complement 
assign ubv = ~UBV;  //complement 
assign ubw = ~UBW;  //complement 
assign ubx = ~UBX;  //complement 
assign vbh = ~VBH;  //complement 
assign vbp = ~VBP;  //complement 
assign hjh = vah & ~ljb & ~lja & ljc |  vbh & ~ljb & lja & ljc |  vch & ljb & ~lja & ljc |  vdh & ljb & lja & ljc; 
assign HJH = ~hjh;  //complement 
assign hph = vah & ~lpb & ~lpa & lpc |         vbh & ~lpb & lpa & lpc |  vch & lpb & ~lpa & lpc |  vdh & lpb & lpa & lpc; 
assign HPH = ~hph;  //complement 
assign hji = vha & ~LJB & ~LJA & LJC |  vga & ~LJB & LJA & LJC |  vfa & LJB & ~LJA & LJC |  vea & LJB & LJA & LJC; 
assign HJI = ~hji;  //complement 
assign hpi = vha & ~LPB & ~LPA & LPC |         vga & ~LPB & LPA & LPC |  vfa & LPB & ~LPA & LPC |  vea & LPB & LPA & LPC; 
assign HPI = ~hpi;  //complement 
assign HAI = ZZO & ~LAB & ~LAA & LAC |  KFA & ~LAB & LAA & LAC |  KEA & LAB & ~LAA & LAC |  KDA & LAB & LAA & LAC; 
assign hai = ~HAI;  //complement 
assign HBI = ZZO & ~LBB & ~LBA & LBC |         KFA & ~LBB & LBA & LBC |  KEA & LBB & ~LBA & LBC |  KDA & LBB & LBA & LBC; 
assign hbi = ~HBI;  //complement 
assign wba = ~WBA;  //complement 
assign wbb = ~WBB;  //complement 
assign hjj = vhb & ~LJB & ~LJA & LJC |  vgb & ~LJB & LJA & LJC |  vfb & LJB & ~LJA & LJC |  veb & LJB & LJA & LJC; 
assign HJJ = ~hjj;  //complement 
assign hpj = vhb & ~LPB & ~LPA & LPC |         vgb & ~LPB & LPA & LPC |  vfb & LPB & ~LPA & LPC |  veb & LPB & LPA & LPC; 
assign HPJ = ~hpj;  //complement 
assign HAJ = ZZO & ~LAB & ~LAA & LAC |  KFB & ~LAB & LAA & LAC |  KEB & LAB & ~LAA & LAC |  KDB & LAB & LAA & LAC; 
assign haj = ~HAJ;  //complement 
assign HBJ = ZZO & ~LBB & ~LBA & LBC |         KFB & ~LBB & LBA & LBC |  KEB & LBB & ~LBA & LBC |  KDB & LBB & LBA & LBC; 
assign hbj = ~HBJ;  //complement 
assign dbm = ~DBM;  //complement 
assign dbn = ~DBN;  //complement 
assign tba = ~TBA;  //complement 
assign tbb = ~TBB;  //complement 
assign hjk = vhc & ~LJB & ~LJA & LJC |  vgc & ~LJB & LJA & LJC |  vfc & LJB & ~LJA & LJC |  vec & LJB & LJA & LJC; 
assign HJK = ~hjk;  //complement 
assign hpk = vhc & ~LPB & ~LPA & LPC |         vgc & ~LPB & LPA & LPC |  vfc & LPB & ~LPA & LPC |  vec & LPB & LPA & LPC; 
assign HPK = ~hpk;  //complement 
assign HAK = ZZO & ~LAB & ~LAA & LAC |  KFC & ~LAB & LAA & LAC |  KEC & LAB & ~LAA & LAC |  KDC & LAB & LAA & LAC; 
assign hak = ~HAK;  //complement 
assign HBK = ZZO & ~LBB & ~LBA & LBC |         KFC & ~LBB & LBA & LBC |  KEC & LBB & ~LBA & LBC |  KDC & LBB & LBA & LBC; 
assign hbk = ~HBK;  //complement 
assign KBA = ~kba;  //complement 
assign KBB = ~kbb;  //complement 
assign KBC = ~kbc;  //complement 
assign KBD = ~kbd;  //complement 
assign lja = ~LJA;  //complement 
assign ljb = ~LJB;  //complement 
assign ljc = ~LJC;  //complement 
assign HAL = ZZO & ~LAB & ~LAA & LAC |  KFD & ~LAB & LAA & LAC |  KED & LAB & ~LAA & LAC |  KDD & LAB & LAA & LAC; 
assign hal = ~HAL;  //complement 
assign HBL = ZZO & ~LBB & ~LBA & LBC |         KFD & ~LBB & LBA & LBC |  KED & LBB & ~LBA & LBC |  KDD & LBB & LBA & LBC; 
assign hbl = ~HBL;  //complement 
assign wbc = ~WBC;  //complement 
assign wbd = ~WBD;  //complement 
assign hjm = vhe & ~LJB & ~LJA & LJC |  vge & ~LJB & LJA & LJC |  vfe & LJB & ~LJA & LJC |  vee & LJB & LJA & LJC; 
assign HJM = ~hjm;  //complement 
assign hpm = vhe & ~LPB & ~LPA & LPC |         vge & ~LPB & LPA & LPC |  vfe & LPB & ~LPA & LPC |  vee & LPB & LPA & LPC; 
assign HPM = ~hpm;  //complement 
assign lpa = ~LPA;  //complement 
assign lpb = ~LPB;  //complement 
assign lpc = ~LPC;  //complement 
assign HAM = ZZO & ~LAB & ~LAA & LAC |  KFE & ~LAB & LAA & LAC |  KEE & LAB & ~LAA & LAC |  KDE & LAB & LAA & LAC; 
assign ham = ~HAM;  //complement 
assign HBM = ZZO & ~LBB & ~LBA & LBC |         KFE & ~LBB & LBA & LBC |  KEE & LBB & ~LBA & LBC |  KDE & LBB & LBA & LBC; 
assign hbm = ~HBM;  //complement 
assign wbe = ~WBE;  //complement 
assign wbf = ~WBF;  //complement 
assign hjn = vhf & ~LJB & ~LJA & LJC |  vgf & ~LJB & LJA & LJC |  vff & LJB & ~LJA & LJC |  vef & LJB & LJA & LJC; 
assign HJN = ~hjn;  //complement 
assign hpn = vhf & ~LPB & ~LPA & LPC |         vgf & ~LPB & LPA & LPC |  vff & LPB & ~LPA & LPC |  vef & LPB & LPA & LPC; 
assign HPN = ~hpn;  //complement 
assign HAN = ZZO & ~LAB & ~LAA & LAC |  KFF & ~LAB & LAA & LAC |  KEF & LAB & ~LAA & LAC |  KDF & LAB & LAA & LAC; 
assign han = ~HAN;  //complement 
assign HBN = ZZO & ~LBB & ~LBA & LBC |         KFF & ~LBB & LBA & LBC |  KEF & LBB & ~LBA & LBC |  KDF & LBB & LBA & LBC; 
assign hbn = ~HBN;  //complement 
assign dbo = ~DBO;  //complement 
assign dbp = ~DBP;  //complement 
assign tbc = ~TBC;  //complement 
assign tbd = ~TBD;  //complement 
assign hjo = vhg & ~LJB & ~LJA & LJC |  vgg & ~LJB & LJA & LJC |  vfg & LJB & ~LJA & LJC |  veg & LJB & LJA & LJC; 
assign HJO = ~hjo;  //complement 
assign hpo = vhg & ~LPB & ~LPA & LPC |         vgg & ~LPB & LPA & LPC |  vfg & LPB & ~LPA & LPC |  veg & LPB & LPA & LPC; 
assign HPO = ~hpo;  //complement 
assign hpl = vhd & ~LPB & ~LPA & LPC |  vgd & ~LPB & LPA & LPC |  vfd & LPB & ~LPA & LPC |  ved & LPB & LPA & LPC; 
assign HPL = ~hpl;  //complement 
assign hql = vhd & ~LQB & ~LQA & LQC |         vgd & ~LQB & LQA & LQC |  vfd & LQB & ~LQA & LQC |  ved & LQB & LQA & LQC; 
assign HQL = ~hql;  //complement 
assign HAO = ZZO & ~LAB & ~LAA & LAC |  KFG & ~LAB & LAA & LAC |  KEG & LAB & ~LAA & LAC |  KDG & LAB & LAA & LAC; 
assign hao = ~HAO;  //complement 
assign HBO = ZZO & ~LBB & ~LBA & LBC |         KFG & ~LBB & LBA & LBC |  KEG & LBB & ~LBA & LBC |  KDG & LBB & LBA & LBC; 
assign hbo = ~HBO;  //complement 
assign KBE = ~kbe;  //complement 
assign KBF = ~kbf;  //complement 
assign KBG = ~kbg;  //complement 
assign KBH = ~kbh;  //complement 
assign hjp = vhh & ~LJB & ~LJA & LJC |  vgh & ~LJB & LJA & LJC |  vfh & LJB & ~LJA & LJC |  veh & LJB & LJA & LJC; 
assign HJP = ~hjp;  //complement 
assign hpp = vhh & ~LPB & ~LPA & LPC |         vgh & ~LPB & LPA & LPC |  vfh & LPB & ~LPA & LPC |  veh & LPB & LPA & LPC; 
assign HPP = ~hpp;  //complement 
assign HAP = ZZO & ~LAB & ~LAA & LAC |  KFH & ~LAB & LAA & LAC |  KEH & LAB & ~LAA & LAC |  KDH & LAB & LAA & LAC; 
assign hap = ~HAP;  //complement 
assign HBP = ZZO & ~LBB & ~LBA & LBC |         KFH & ~LBB & LBA & LBC |  KEH & LBB & ~LBA & LBC |  KDH & LBB & LBA & LBC; 
assign hbp = ~HBP;  //complement 
assign wbg = ~WBG;  //complement 
assign wbh = ~WBH;  //complement 
assign ona = ~ONA;  //complement 
assign ooa = ~OOA;  //complement 
assign DBI = ~dbi;  //complement 
assign DBJ = ~dbj;  //complement 
assign DBK = ~dbk;  //complement 
assign DBL = ~dbl;  //complement 
assign onb = ~ONB;  //complement 
assign oob = ~OOB;  //complement 
assign sea = ~SEA;  //complement 
assign seb = ~SEB;  //complement 
assign gab = ~GAB;  //complement 
assign gaj = ~GAJ;  //complement 
assign onc = ~ONC;  //complement 
assign ooc = ~OOC;  //complement 
assign sfa = ~SFA;  //complement 
assign sfb = ~SFB;  //complement 
assign MAB =  SJB & SKB & QDA  |  SJB & skb & QDB  |  sjb & SKB & QDC  ; 
assign mab = ~MAB; //complement 
assign ond = ~OND;  //complement 
assign ood = ~OOD;  //complement 
assign JBA =  SEA & NEA  |  SFA & NFA  |  SGA & NGA  |  SHA & NHA  ; 
assign jba = ~JBA;  //complement 
assign JBI =  SEA & NEA  |  SFA & NFA  |  SGA & NGA  |  SHA & NHA  ; 
assign jbi = ~JBI; //complement 
assign nea = ~NEA;  //complement 
assign nga = ~NGA;  //complement 
assign qdb = ~QDB;  //complement 
assign sjb = ~SJB;  //complement 
assign one = ~ONE;  //complement 
assign ooe = ~OOE;  //complement 
assign JBB =  SEB & NEA  |  SFB & NFA  |  SGB & NGA  |  SHB & NHA  ; 
assign jbb = ~JBB;  //complement 
assign JBJ =  SEB & NEA  |  SFB & NFA  |  SGB & NGA  |  SHB & NHA  ; 
assign jbj = ~JBJ; //complement 
assign dbg = ~DBG;  //complement 
assign nfa = ~NFA;  //complement 
assign nha = ~NHA;  //complement 
assign onf = ~ONF;  //complement 
assign oof = ~OOF;  //complement 
assign sga = ~SGA;  //complement 
assign sgb = ~SGB;  //complement 
assign OAB = ~oab;  //complement 
assign OBB = ~obb;  //complement 
assign OCB = ~ocb;  //complement 
assign SKB = ~skb;  //complement 
assign ong = ~ONG;  //complement 
assign oog = ~OOG;  //complement 
assign sha = ~SHA;  //complement 
assign shb = ~SHB;  //complement 
assign gbb = ~GBB;  //complement 
assign gbj = ~GBJ;  //complement 
assign onh = ~ONH;  //complement 
assign ooh = ~OOH;  //complement 
assign lba = ~LBA;  //complement 
assign lbb = ~LBB;  //complement 
assign lbc = ~LBC;  //complement 
assign dbc = ~DBC;  //complement 
assign dbd = ~DBD;  //complement 
assign dbe = ~DBE;  //complement 
assign dbf = ~DBF;  //complement 
assign uca = ~UCA;  //complement 
assign ucb = ~UCB;  //complement 
assign ucc = ~UCC;  //complement 
assign vca = ~VCA;  //complement 
assign vci = ~VCI;  //complement 
assign hka = vaa & ~lkb & ~lka & lkc |  vba & ~lkb & lka & lkc |  vca & lkb & ~lka & lkc |  vda & lkb & lka & lkc; 
assign HKA = ~hka;  //complement 
assign hqa = vaa & ~lqb & ~lqa & lqc |         vba & ~lqb & lqa & lqc |  vca & lqb & ~lqa & lqc |  vda & lqb & lqa & lqc; 
assign HQA = ~hqa;  //complement 
assign ucd = ~UCD;  //complement 
assign uce = ~UCE;  //complement 
assign ucf = ~UCF;  //complement 
assign vcb = ~VCB;  //complement 
assign vcj = ~VCJ;  //complement 
assign hkb = vab & ~lkb & ~lka & lkc |  vbb & ~lkb & lka & lkc |  vcb & lkb & ~lka & lkc |  vdb & lkb & lka & lkc; 
assign HKB = ~hkb;  //complement 
assign hqb = vab & ~lqb & ~lqa & lqc |         vbb & ~lqb & lqa & lqc |  vcb & lqb & ~lqa & lqc |  vdb & lqb & lqa & lqc; 
assign HQB = ~hqb;  //complement 
assign ucg = ~UCG;  //complement 
assign uci = ~UCI;  //complement 
assign uch = ~UCH;  //complement 
assign vcc = ~VCC;  //complement 
assign vck = ~VCK;  //complement 
assign hkc = vac & ~lkb & ~lka & lkc |  vbc & ~lkb & lka & lkc |  vcc & lkb & ~lka & lkc |  vdc & lkb & lka & lkc; 
assign HKC = ~hkc;  //complement 
assign hqc = vac & ~lqb & ~lqa & lqc |         vbc & ~lqb & lqa & lqc |  vcc & lqb & ~lqa & lqc |  vdc & lqb & lqa & lqc; 
assign HQC = ~hqc;  //complement 
assign ucj = ~UCJ;  //complement 
assign uck = ~UCK;  //complement 
assign ucl = ~UCL;  //complement 
assign vcd = ~VCD;  //complement 
assign vcl = ~VCL;  //complement 
assign hkd = vad & ~lkb & ~lka & lkc |  vbd & ~lkb & lka & lkc |  vcd & lkb & ~lka & lkc |  vdd & lkb & lka & lkc; 
assign HKD = ~hkd;  //complement 
assign hqd = vad & ~lqb & ~lqa & lqc |         vbd & ~lqb & lqa & lqc |  vcd & lqb & ~lqa & lqc |  vdd & lqb & lqa & lqc; 
assign HQD = ~hqd;  //complement 
assign ucm = ~UCM;  //complement 
assign ucn = ~UCN;  //complement 
assign uco = ~UCO;  //complement 
assign vce = ~VCE;  //complement 
assign vcm = ~VCM;  //complement 
assign hke = vae & ~lkb & ~lka & lkc |  vbe & ~lkb & lka & lkc |  vce & lkb & ~lka & lkc |  vde & lkb & lka & lkc; 
assign HKE = ~hke;  //complement 
assign ucp = ~UCP;  //complement 
assign ucq = ~UCQ;  //complement 
assign ucr = ~UCR;  //complement 
assign vcf = ~VCF;  //complement 
assign vcn = ~VCN;  //complement 
assign hkf = vaf & ~lkb & ~lka & lkc |  vbf & ~lkb & lka & lkc |  vcf & lkb & ~lka & lkc |  vdf & lkb & lka & lkc; 
assign HKF = ~hkf;  //complement 
assign hqf = vaf & ~lqb & ~lqa & lqc |         vbf & ~lqb & lqa & lqc |  vcf & lqb & ~lqa & lqc |  vdf & lqb & lqa & lqc; 
assign HQF = ~hqf;  //complement 
assign ucs = ~UCS;  //complement 
assign uct = ~UCT;  //complement 
assign ucu = ~UCU;  //complement 
assign vch = ~VCH;  //complement 
assign vcp = ~VCP;  //complement 
assign hkg = vag & ~lkb & ~lka & lkc |  vbg & ~lkb & lka & lkc |  vcg & lkb & ~lka & lkc |  vdg & lkb & lka & lkc; 
assign HKG = ~hkg;  //complement 
assign hqg = vag & ~lqb & ~lqa & lqc |         vbg & ~lqb & lqa & lqc |  vcg & lqb & ~lqa & lqc |  vdg & lqb & lqa & lqc; 
assign HQG = ~hqg;  //complement 
assign ucv = ~UCV;  //complement 
assign ucw = ~UCW;  //complement 
assign ucx = ~UCX;  //complement 
assign vcg = ~VCG;  //complement 
assign vco = ~VCO;  //complement 
assign hkh = vah & ~lkb & ~lka & lkc |  vbh & ~lkb & lka & lkc |  vch & lkb & ~lka & lkc |  vdh & lkb & lka & lkc; 
assign HKH = ~hkh;  //complement 
assign hqh = vah & ~lqb & ~lqa & lqc |         vbh & ~lqb & lqa & lqc |  vch & lqb & ~lqa & lqc |  vdh & lqb & lqa & lqc; 
assign HQH = ~hqh;  //complement 
assign hki = vha & ~LKB & ~LKA & LKC |  vga & ~LKB & LKA & LKC |  vfa & LKB & ~LKA & LKC |  vea & LKB & LKA & LKC; 
assign HKI = ~hki;  //complement 
assign hqi = vha & ~LQB & ~LQA & LQC |         vga & ~LQB & LQA & LQC |  vfa & LQB & ~LQA & LQC |  vea & LQB & LQA & LQC; 
assign HQI = ~hqi;  //complement 
assign dcm = ~DCM;  //complement 
assign dcn = ~DCN;  //complement 
assign tca = ~TCA;  //complement 
assign tcb = ~TCB;  //complement 
assign HCA = ZZO & ~lcb & ~lca & lcc |  KAA & ~lcb & lca & lcc |  KBA & lcb & ~lca & lcc |  KCA & lcb & lca & lcc; 
assign hca = ~HCA;  //complement 
assign HDA = ZZO & ~ldb & ~lda & ldc |         KAA & ~ldb & lda & ldc |  KBA & ldb & ~lda & ldc |  KCA & ldb & lda & ldc; 
assign hda = ~HDA;  //complement 
assign wca = ~WCA;  //complement 
assign wcb = ~WCB;  //complement 
assign hkj = vhb & ~LKB & ~LKA & LKC |  vgb & ~LKB & LKA & LKC |  vfb & LKB & ~LKA & LKC |  veb & LKB & LKA & LKC; 
assign HKJ = ~hkj;  //complement 
assign hqj = vhb & ~LQB & ~LQA & LQC |         vgb & ~LQB & LQA & LQC |  vfb & LQB & ~LQA & LQC |  veb & LQB & LQA & LQC; 
assign HQJ = ~hqj;  //complement 
assign HCB = ZZO & ~lcb & ~lca & lcc |  KAB & ~lcb & lca & lcc |  KBB & lcb & ~lca & lcc |  KCB & lcb & lca & lcc; 
assign hcb = ~HCB;  //complement 
assign HDB = ZZO & ~ldb & ~lda & ldc |         KAB & ~ldb & lda & ldc |  KBB & ldb & ~lda & ldc |  KCB & ldb & lda & ldc; 
assign hdb = ~HDB;  //complement 
assign HCF = ZZO & ~lcb & ~lca & lcc |  KAF & ~lcb & lca & lcc |  KBF & lcb & ~lca & lcc |  KCF & lcb & lca & lcc; 
assign hcf = ~HCF;  //complement 
assign HDF = ZZO & ~ldb & ~lda & ldc |         KAF & ~ldb & lda & ldc |  KBF & ldb & ~lda & ldc |  KCF & ldb & lda & ldc; 
assign hdf = ~HDF;  //complement 
assign hkk = vhc & ~LKB & ~LKA & LKC |  vgc & ~LKB & LKA & LKC |  vfc & LKB & ~LKA & LKC |  vec & LKB & LKA & LKC; 
assign HKK = ~hkk;  //complement 
assign hqk = vhc & ~LQB & ~LQA & LQC |         vgc & ~LQB & LQA & LQC |  vfc & LQB & ~LQA & LQC |  vec & LQB & LQA & LQC; 
assign HQK = ~hqk;  //complement 
assign HGM = ZZO & ~LGB & ~LGA & LGC |  KFE & ~LGB & LGA & LGC |  KEE & LGB & ~LGA & LGC |  KDE & LGB & LGA & LGC; 
assign hgm = ~HGM;  //complement 
assign HHM = ZZO & ~LHB & ~LHA & LHC |         KFE & ~LHB & LHA & LHC |  KEE & LHB & ~LHA & LHC |  KDE & LHB & LHA & LHC; 
assign hhm = ~HHM;  //complement 
assign HCC = ZZO & ~lcb & ~lca & lcc |  KAC & ~lcb & lca & lcc |  KBC & lcb & ~lca & lcc |  KCC & lcb & lca & lcc; 
assign hcc = ~HCC;  //complement 
assign HDC = ZZO & ~ldb & ~lda & ldc |         KAC & ~ldb & lda & ldc |  KBC & ldb & ~lda & ldc |  KCC & ldb & lda & ldc; 
assign hdc = ~HDC;  //complement 
assign KCA = ~kca;  //complement 
assign KCB = ~kcb;  //complement 
assign KCC = ~kcc;  //complement 
assign KCD = ~kcd;  //complement 
assign hnl = vhl & ~LNB & ~LNA & LNC |  vgl & ~LNB & LNA & LNC |  vfl & LNB & ~LNA & LNC |  vel & LNB & LNA & LNC; 
assign HNL = ~hnl;  //complement 
assign hml = vhl & ~LMB & ~LMA & LMC |         vgl & ~LMB & LMA & LMC |  vfl & LMB & ~LMA & LMC |  vel & LMB & LMA & LMC; 
assign HML = ~hml;  //complement 
assign lka = ~LKA;  //complement 
assign lkb = ~LKB;  //complement 
assign lkc = ~LKC;  //complement 
assign HCD = ZZO & ~lcb & ~lca & lcc |  KAD & ~lcb & lca & lcc |  KBD & lcb & ~lca & lcc |  KCD & lcb & lca & lcc; 
assign hcd = ~HCD;  //complement 
assign HDD = ZZO & ~ldb & ~lda & ldc |         KAD & ~ldb & lda & ldc |  KBD & ldb & ~lda & ldc |  KCD & ldb & lda & ldc; 
assign hdd = ~HDD;  //complement 
assign wcc = ~WCC;  //complement 
assign wcd = ~WCD;  //complement 
assign hkm = vhe & ~LKB & ~LKA & LKC |  vge & ~LKB & LKA & LKC |  vfe & LKB & ~LKA & LKC |  vee & LKB & LKA & LKC; 
assign HKM = ~hkm;  //complement 
assign hqm = vhe & ~LQB & ~LQA & LQC |         vge & ~LQB & LQA & LQC |  vfe & LQB & ~LQA & LQC |  vee & LQB & LQA & LQC; 
assign HQM = ~hqm;  //complement 
assign lqa = ~LQA;  //complement 
assign lqb = ~LQB;  //complement 
assign lqc = ~LQC;  //complement 
assign HCE = ZZO & ~lcb & ~lca & lcc |  KAE & ~lcb & lca & lcc |  KBE & lcb & ~lca & lcc |  KCE & lcb & lca & lcc; 
assign hce = ~HCE;  //complement 
assign HDE = ZZO & ~ldb & ~lda & ldc |         KAE & ~ldb & lda & ldc |  KBE & ldb & ~lda & ldc |  KCE & ldb & lda & ldc; 
assign hde = ~HDE;  //complement 
assign wce = ~WCE;  //complement 
assign wcf = ~WCF;  //complement 
assign hkn = vhf & ~LKB & ~LKA & LKC |  vgf & ~LKB & LKA & LKC |  vff & LKB & ~LKA & LKC |  vef & LKB & LKA & LKC; 
assign HKN = ~hkn;  //complement 
assign hqn = vhf & ~LQB & ~LQA & LQC |         vgf & ~LQB & LQA & LQC |  vff & LQB & ~LQA & LQC |  vef & LQB & LQA & LQC; 
assign HQN = ~hqn;  //complement 
assign hkl = vhd & ~LKB & ~LKA & LKC |  vgd & ~LKB & LKA & LKC |  vfd & LKB & ~LKA & LKC |  ved & LKB & LKA & LKC; 
assign HKL = ~hkl;  //complement 
assign hjl = vhd & ~LJB & ~LJA & LJC |         vgd & ~LJB & LJA & LJC |  vfd & LJB & ~LJA & LJC |  ved & LJB & LJA & LJC; 
assign HJL = ~hjl;  //complement 
assign dco = ~DCO;  //complement 
assign dcp = ~DCP;  //complement 
assign tcc = ~TCC;  //complement 
assign tcd = ~TCD;  //complement 
assign hko = vhg & ~LKB & ~LKA & LKC |  vgg & ~LKB & LKA & LKC |  vfg & LKB & ~LKA & LKC |  veg & LKB & LKA & LKC; 
assign HKO = ~hko;  //complement 
assign hqo = vhg & ~LQB & ~LQA & LQC |         vgg & ~LQB & LQA & LQC |  vfg & LQB & ~LQA & LQC |  veg & LQB & LQA & LQC; 
assign HQO = ~hqo;  //complement 
assign hje = vad & ~ljb & ~lja & ljc |  vbe & ~ljb & lja & ljc |  vce & ljb & ~lja & ljc |  vde & ljb & lja & ljc; 
assign HJE = ~hje;  //complement 
assign HCG = ZZO & ~lcb & ~lca & lcc |  KAG & ~lcb & lca & lcc |  KBG & lcb & ~lca & lcc |  KCG & lcb & lca & lcc; 
assign hcg = ~HCG;  //complement 
assign HDG = ZZO & ~ldb & ~lda & ldc |         KAG & ~ldb & lda & ldc |  KBG & ldb & ~lda & ldc |  KCG & ldb & lda & ldc; 
assign hdg = ~HDG;  //complement 
assign KCE = ~kce;  //complement 
assign KCF = ~kcf;  //complement 
assign KCG = ~kcg;  //complement 
assign KCH = ~kch;  //complement 
assign hkp = vhh & ~LKB & ~LKA & LKC |  vgh & ~LKB & LKA & LKC |  vfh & LKB & ~LKA & LKC |  veh & LKB & LKA & LKC; 
assign HKP = ~hkp;  //complement 
assign hqp = vhh & ~LQB & ~LQA & LQC |         vgh & ~LQB & LQA & LQC |  vfh & LQB & ~LQA & LQC |  veh & LQB & LQA & LQC; 
assign HQP = ~hqp;  //complement 
assign HCH = ZZO & ~lcb & ~lca & lcc |  KAH & ~lcb & lca & lcc |  KBH & lcb & ~lca & lcc |  KCH & lcb & lca & lcc; 
assign hch = ~HCH;  //complement 
assign HDH = ZZO & ~ldb & ~lda & ldc |         KAH & ~ldb & lda & ldc |  KBH & ldb & ~lda & ldc |  KCH & ldb & lda & ldc; 
assign hdh = ~HDH;  //complement 
assign wcg = ~WCG;  //complement 
assign wch = ~WCH;  //complement 
assign oda = ~ODA;  //complement 
assign oma = ~OMA;  //complement 
assign DCI = ~dci;  //complement 
assign DCJ = ~dcj;  //complement 
assign DCK = ~dck;  //complement 
assign DCL = ~dcl;  //complement 
assign odb = ~ODB;  //complement 
assign omb = ~OMB;  //complement 
assign sac = ~SAC;  //complement 
assign sad = ~SAD;  //complement 
assign gac = ~GAC;  //complement 
assign gak = ~GAK;  //complement 
assign odc = ~ODC;  //complement 
assign omc = ~OMC;  //complement 
assign sbc = ~SBC;  //complement 
assign sbd = ~SBD;  //complement 
assign MAC =  SJC & SKC & QDA  |  SJC & skc & QDB  |  sjc & SKC & QDC  ; 
assign mac = ~MAC; //complement 
assign odd = ~ODD;  //complement 
assign omd = ~OMD;  //complement 
assign JAC =  SAC & NAB  |  SBC & NBB  |  SCC & NCB  |  SDC & NDB  ; 
assign jac = ~JAC;  //complement 
assign JAK =  SAC & NAB  |  SBC & NBB  |  SCC & NCB  |  SDC & NDB  ; 
assign jak = ~JAK; //complement 
assign nab = ~NAB;  //complement 
assign ncb = ~NCB;  //complement 
assign qdc = ~QDC;  //complement 
assign sjc = ~SJC;  //complement 
assign ode = ~ODE;  //complement 
assign ome = ~OME;  //complement 
assign JAL =  SAD & NAB  |  SBD & NBB  |  SCD & NCB  |  SDD & NDB  ; 
assign jal = ~JAL;  //complement 
assign JAD =  SAD & NAB  |  SBD & NBB  |  SCD & NCB  |  SDD & NDB  ; 
assign jad = ~JAD; //complement 
assign dcg = ~DCG;  //complement 
assign nbb = ~NBB;  //complement 
assign ndb = ~NDB;  //complement 
assign odf = ~ODF;  //complement 
assign omf = ~OMF;  //complement 
assign scc = ~SCC;  //complement 
assign scd = ~SCD;  //complement 
assign OAC = ~oac;  //complement 
assign OBC = ~obc;  //complement 
assign OCC = ~occ;  //complement 
assign SKC = ~skc;  //complement 
assign odg = ~ODG;  //complement 
assign omg = ~OMG;  //complement 
assign sdc = ~SDC;  //complement 
assign sdd = ~SDD;  //complement 
assign gbc = ~GBC;  //complement 
assign gbk = ~GBK;  //complement 
assign odh = ~ODH;  //complement 
assign omh = ~OMH;  //complement 
assign lca = ~LCA;  //complement 
assign lcb = ~LCB;  //complement 
assign lcc = ~LCC;  //complement 
assign dcc = ~DCC;  //complement 
assign dcd = ~DCD;  //complement 
assign dce = ~DCE;  //complement 
assign dcf = ~DCF;  //complement 
assign uda = ~UDA;  //complement 
assign udb = ~UDB;  //complement 
assign udc = ~UDC;  //complement 
assign vda = ~VDA;  //complement 
assign vdi = ~VDI;  //complement 
assign udd = ~UDD;  //complement 
assign ude = ~UDE;  //complement 
assign udf = ~UDF;  //complement 
assign vdb = ~VDB;  //complement 
assign vdj = ~VDJ;  //complement 
assign udg = ~UDG;  //complement 
assign udh = ~UDH;  //complement 
assign udi = ~UDI;  //complement 
assign vdc = ~VDC;  //complement 
assign vdk = ~VDK;  //complement 
assign udj = ~UDJ;  //complement 
assign udk = ~UDK;  //complement 
assign udl = ~UDL;  //complement 
assign vdd = ~VDD;  //complement 
assign vdl = ~VDL;  //complement 
assign udm = ~UDM;  //complement 
assign udn = ~UDN;  //complement 
assign udo = ~UDO;  //complement 
assign vde = ~VDE;  //complement 
assign vdm = ~VDM;  //complement 
assign udp = ~UDP;  //complement 
assign udq = ~UDQ;  //complement 
assign udr = ~UDR;  //complement 
assign vdf = ~VDF;  //complement 
assign vdn = ~VDN;  //complement 
assign uds = ~UDS;  //complement 
assign udt = ~UDT;  //complement 
assign udu = ~UDU;  //complement 
assign vdg = ~VDG;  //complement 
assign vdo = ~VDO;  //complement 
assign udv = ~UDV;  //complement 
assign udw = ~UDW;  //complement 
assign udx = ~UDX;  //complement 
assign vdh = ~VDH;  //complement 
assign vdp = ~VDP;  //complement 
assign HCI = ZZO & ~LCB & ~LCA & LCC |  KFA & ~LCB & LCA & LCC |  KEA & LCB & ~LCA & LCC |  KDA & LCB & LCA & LCC; 
assign hci = ~HCI;  //complement 
assign HDI = ZZO & ~LDB & ~LDA & LDC |         KFA & ~LDB & LDA & LDC |  KEA & LDB & ~LDA & LDC |  KDA & LDB & LDA & LDC; 
assign hdi = ~HDI;  //complement 
assign wda = ~WDA;  //complement 
assign wdb = ~WDB;  //complement 
assign jea = kba; 
assign JEA = ~jea; //complement 
assign jeb = kbb; 
assign JEB = ~jeb;  //complement 
assign jec = kbc; 
assign JEC = ~jec;  //complement 
assign jed = kbd; 
assign JED = ~jed;  //complement 
assign HCJ = ZZO & ~LCB & ~LCA & LCC |  KFB & ~LCB & LCA & LCC |  KEB & LCB & ~LCA & LCC |  KDB & LCB & LCA & LCC; 
assign hcj = ~HCJ;  //complement 
assign HDJ = ZZO & ~LDB & ~LDA & LDC |         KFB & ~LDB & LDA & LDC |  KEB & LDB & ~LDA & LDC |  KDB & LDB & LDA & LDC; 
assign hdj = ~HDJ;  //complement 
assign ddm = ~DDM;  //complement 
assign tda = ~TDA;  //complement 
assign qea = ~QEA;  //complement 
assign HCK = ZZO & ~LCB & ~LCA & LCC |  KFC & ~LCB & LCA & LCC |  KEC & LCB & ~LCA & LCC |  KDC & LCB & LCA & LCC; 
assign hck = ~HCK;  //complement 
assign HDK = ZZO & ~LDB & ~LDA & LDC |         KFC & ~LDB & LDA & LDC |  KEC & LDB & ~LDA & LDC |  KDC & LDB & LDA & LDC; 
assign hdk = ~HDK;  //complement 
assign ddn = ~DDN;  //complement 
assign tdb = ~TDB;  //complement 
assign qeb = ~QEB;  //complement 
assign QCA = ~qca;  //complement 
assign QCB = ~qcb;  //complement 
assign HCL = ZZO & ~LCB & ~LCA & LCC |  KFD & ~LCB & LCA & LCC |  KED & LCB & ~LCA & LCC |  KDD & LCB & LCA & LCC; 
assign hcl = ~HCL;  //complement 
assign HDL = ZZO & ~LDB & ~LDA & LDC |         KFD & ~LDB & LDA & LDC |  KED & LDB & ~LDA & LDC |  KDD & LDB & LDA & LDC; 
assign hdl = ~HDL;  //complement 
assign wdc = ~WDC;  //complement 
assign wdd = ~WDD;  //complement 
assign qec = ~QEC;  //complement 
assign QCC = ~qcc;  //complement 
assign HCM = ZZO & ~LCB & ~LCA & LCC |  KFE & ~LCB & LCA & LCC |  KEE & LCB & ~LCA & LCC |  KDE & LCB & LCA & LCC; 
assign hcm = ~HCM;  //complement 
assign HDM = ZZO & ~LDB & ~LDA & LDC |         KFE & ~LDB & LDA & LDC |  KEE & LDB & ~LDA & LDC |  KDE & LDB & LDA & LDC; 
assign hdm = ~HDM;  //complement 
assign wde = ~WDE;  //complement 
assign wdf = ~WDF;  //complement 
assign HCN = ZZO & ~LCB & ~LCA & LCC |  KFF & ~LCB & LCA & LCC |  KEF & LCB & ~LCA & LCC |  KDF & LCB & LCA & LCC; 
assign hcn = ~HCN;  //complement 
assign HDN = ZZO & ~LDB & ~LDA & LDC |         KFF & ~LDB & LDA & LDC |  KEF & LDB & ~LDA & LDC |  KDF & LDB & LDA & LDC; 
assign hdn = ~HDN;  //complement 
assign ddo = ~DDO;  //complement 
assign tdc = ~TDC;  //complement 
assign ddp = ~DDP;  //complement 
assign jee = kbe; 
assign JEE = ~jee; //complement 
assign jef = kbf; 
assign JEF = ~jef;  //complement 
assign jeg = kbg; 
assign JEG = ~jeg;  //complement 
assign jeh = kbh; 
assign JEH = ~jeh;  //complement 
assign HCO = ZZO & ~LCB & ~LCA & LCC |  KFG & ~LCB & LCA & LCC |  KEG & LCB & ~LCA & LCC |  KDG & LCB & LCA & LCC; 
assign hco = ~HCO;  //complement 
assign HDO = ZZO & ~LDB & ~LDA & LDC |         KFG & ~LDB & LDA & LDC |  KEG & LDB & ~LDA & LDC |  KDG & LDB & LDA & LDC; 
assign hdo = ~HDO;  //complement 
assign tdd = ~TDD;  //complement 
assign HCP = ZZO & ~LCB & ~LCA & LCC |  KFH & ~LCB & LCA & LCC |  KEH & LCB & ~LCA & LCC |  KDH & LCB & LCA & LCC; 
assign hcp = ~HCP;  //complement 
assign HDP = ZZO & ~LDB & ~LDA & LDC |         KFH & ~LDB & LDA & LDC |  KEH & LDB & ~LDA & LDC |  KDH & LDB & LDA & LDC; 
assign hdp = ~HDP;  //complement 
assign wdg = ~WDG;  //complement 
assign wdh = ~WDH;  //complement 
assign tjb = ~TJB;  //complement 
assign tkb = ~TKB;  //complement 
assign ora = ~ORA;  //complement 
assign DDI = ~ddi;  //complement 
assign DDJ = ~ddj;  //complement 
assign DDK = ~ddk;  //complement 
assign DDL = ~ddl;  //complement 
assign tjc = ~TJC;  //complement 
assign tkc = ~TKC;  //complement 
assign CAE = ~cae;  //complement 
assign sec = ~SEC;  //complement 
assign sed = ~SED;  //complement 
assign gad = ~GAD;  //complement 
assign gal = ~GAL;  //complement 
assign tjd = ~TJD;  //complement 
assign tkd = ~TKD;  //complement 
assign CAF = ~caf;  //complement 
assign CAG = ~cag;  //complement 
assign sfc = ~SFC;  //complement 
assign sfd = ~SFD;  //complement 
assign MAD =  SJD & SKD & QDA  |  SJD & skd & QDB  |  sjd & SKD & QDC  ; 
assign mad = ~MAD; //complement 
assign CAH = ~cah;  //complement 
assign CAI = ~cai;  //complement 
assign JBC =  SEC & NEB  |  SFC & NFB  |  SGC & NGB  |  SHC & NHB  ; 
assign jbc = ~JBC;  //complement 
assign JBK =  SEC & NEB  |  SFC & NFB  |  SGC & NGB  |  SHC & NHB  ; 
assign jbk = ~JBK; //complement 
assign neb = ~NEB;  //complement 
assign ngb = ~NGB;  //complement 
assign sjd = ~SJD;  //complement 
assign tie = ~TIE;  //complement 
assign tif = ~TIF;  //complement 
assign tig = ~TIG;  //complement 
assign cad = ~CAD;  //complement 
assign CAJ = ~caj;  //complement 
assign JBD =  SED & NEB  |  SFD & NFB  |  SGD & NGB  |  SHD & NHB  ; 
assign jbd = ~JBD;  //complement 
assign JBL =  SED & NEB  |  SFD & NFB  |  SGD & NGB  |  SHD & NHB  ; 
assign jbl = ~JBL; //complement 
assign ddg = ~DDG;  //complement 
assign nfb = ~NFB;  //complement 
assign nhb = ~NHB;  //complement 
assign tje = ~TJE;  //complement 
assign tke = ~TKE;  //complement 
assign eaa =  ska & skb  ; 
assign EAA = ~eaa;  //complement 
assign eab =  skc & skd  ; 
assign EAB = ~eab;  //complement 
assign sgc = ~SGC;  //complement 
assign sgd = ~SGD;  //complement 
assign OAD = ~oad;  //complement 
assign OBD = ~obd;  //complement 
assign OCD = ~ocd;  //complement 
assign SKD = ~skd;  //complement 
assign tjf = ~TJF;  //complement 
assign tkf = ~TKF;  //complement 
assign OQA = ~oqa;  //complement 
assign shc = ~SHC;  //complement 
assign shd = ~SHD;  //complement 
assign gbd = ~GBD;  //complement 
assign gbl = ~GBL;  //complement 
assign tjg = ~TJG;  //complement 
assign tkg = ~TKG;  //complement 
assign lda = ~LDA;  //complement 
assign ldb = ~LDB;  //complement 
assign ldc = ~LDC;  //complement 
assign ddc = ~DDC;  //complement 
assign ddd = ~DDD;  //complement 
assign dde = ~DDE;  //complement 
assign ddf = ~DDF;  //complement 
assign uea = ~UEA;  //complement 
assign ueb = ~UEB;  //complement 
assign uec = ~UEC;  //complement 
assign vea = ~VEA;  //complement 
assign vei = ~VEI;  //complement 
assign ued = ~UED;  //complement 
assign uee = ~UEE;  //complement 
assign uef = ~UEF;  //complement 
assign hmj = vhj & ~LMB & ~LMA & LMC |  vgj & ~LMB & LMA & LMC |  vfj & LMB & ~LMA & LMC |  vej & LMB & LMA & LMC; 
assign HMJ = ~hmj;  //complement 
assign hnj = vhj & ~LNB & ~LNA & LNC |         vgj & ~LNB & LNA & LNC |  vfj & LNB & ~LNA & LNC |  vej & LNB & LNA & LNC; 
assign HNJ = ~hnj;  //complement 
assign veb = ~VEB;  //complement 
assign vej = ~VEJ;  //complement 
assign ueg = ~UEG;  //complement 
assign ueh = ~UEH;  //complement 
assign uei = ~UEI;  //complement 
assign hmk = vhk & ~LMB & ~LMA & LMC |  vgk & ~LMB & LMA & LMC |  vfk & LMB & ~LMA & LMC |  vek & LMB & LMA & LMC; 
assign HMK = ~hmk;  //complement 
assign hnk = vhk & ~LNB & ~LNA & LNC |         vgk & ~LNB & LNA & LNC |  vfk & LNB & ~LNA & LNC |  vek & LNB & LNA & LNC; 
assign HNK = ~hnk;  //complement 
assign vec = ~VEC;  //complement 
assign vek = ~VEK;  //complement 
assign veg = ~VEG;  //complement 
assign veo = ~VEO;  //complement 
assign uej = ~UEJ;  //complement 
assign uek = ~UEK;  //complement 
assign uel = ~UEL;  //complement 
assign ved = ~VED;  //complement 
assign vel = ~VEL;  //complement 
assign uem = ~UEM;  //complement 
assign uen = ~UEN;  //complement 
assign ueo = ~UEO;  //complement 
assign hmm = vhm & ~LMB & ~LMA & LMC |  vgm & ~LMB & LMA & LMC |  vfm & LMB & ~LMA & LMC |  vem & LMB & LMA & LMC; 
assign HMM = ~hmm;  //complement 
assign hnm = vhm & ~LNB & ~LNA & LNC |         vgm & ~LNB & LNA & LNC |  vfm & LNB & ~LNA & LNC |  vem & LNB & LNA & LNC; 
assign HNM = ~hnm;  //complement 
assign vee = ~VEE;  //complement 
assign vem = ~VEM;  //complement 
assign uep = ~UEP;  //complement 
assign ueq = ~UEQ;  //complement 
assign uer = ~UER;  //complement 
assign vef = ~VEF;  //complement 
assign ven = ~VEN;  //complement 
assign ueu = ~UEU;  //complement 
assign ues = ~UES;  //complement 
assign uet = ~UET;  //complement 
assign uev = ~UEV;  //complement 
assign uew = ~UEW;  //complement 
assign uex = ~UEX;  //complement 
assign veh = ~VEH;  //complement 
assign vep = ~VEP;  //complement 
assign HEA = ZZO & ~leb & ~lea & lec |  KAA & ~leb & lea & lec |  KBA & leb & ~lea & lec |  KCA & leb & lea & lec; 
assign hea = ~HEA;  //complement 
assign HFA = ZZO & ~lfb & ~lfa & lfc |         KAA & ~lfb & lfa & lfc |  KBA & lfb & ~lfa & lfc |  KCA & lfb & lfa & lfc; 
assign hfa = ~HFA;  //complement 
assign wea = ~WEA;  //complement 
assign web = ~WEB;  //complement 
assign HEB = ZZO & ~leb & ~lea & lec |  KAB & ~leb & lea & lec |  KBB & leb & ~lea & lec |  KCB & leb & lea & lec; 
assign heb = ~HEB;  //complement 
assign HFB = ZZO & ~lfb & ~lfa & lfc |         KAB & ~lfb & lfa & lfc |  KBB & lfb & ~lfa & lfc |  KCB & lfb & lfa & lfc; 
assign hfb = ~HFB;  //complement 
assign dem = ~DEM;  //complement 
assign tea = ~TEA;  //complement 
assign teb = ~TEB;  //complement 
assign HEC = ZZO & ~leb & ~lea & lec |  KAC & ~leb & lea & lec |  KBC & leb & ~lea & lec |  KCC & leb & lea & lec; 
assign hec = ~HEC;  //complement 
assign HFC = ZZO & ~lfb & ~lfa & lfc |         KAC & ~lfb & lfa & lfc |  KBC & lfb & ~lfa & lfc |  KCC & lfb & lfa & lfc; 
assign hfc = ~HFC;  //complement 
assign den = ~DEN;  //complement 
assign baj = ~BAJ;  //complement 
assign bak = ~BAK;  //complement 
assign bal = ~BAL;  //complement 
assign bba = ~BBA;  //complement 
assign bbb = ~BBB;  //complement 
assign bbc = ~BBC;  //complement 
assign HED = ZZO & ~leb & ~lea & lec |  KAD & ~leb & lea & lec |  KBD & leb & ~lea & lec |  KCD & leb & lea & lec; 
assign hed = ~HED;  //complement 
assign HFD = ZZO & ~lfb & ~lfa & lfc |         KAD & ~lfb & lfa & lfc |  KBD & lfb & ~lfa & lfc |  KCD & lfb & lfa & lfc; 
assign hfd = ~HFD;  //complement 
assign wec = ~WEC;  //complement 
assign wed = ~WED;  //complement 
assign bam = ~BAM;  //complement 
assign ban = ~BAN;  //complement 
assign bao = ~BAO;  //complement 
assign bap = ~BAP;  //complement 
assign FCH = ~aaf & ~aae & ~aad & QAA ; 
assign FCG = ~aaf & ~aae &  aad & QAA ; 
assign FCF = ~aaf &  aae & ~aad & QAA ; 
assign FCE = ~aaf &  aae &  aad & QAA ; 
assign FCD =  aaf & ~aae & ~aad & QAA ; 
assign FCC =  aaf & ~aae &  aad & QAA ; 
assign FCB =  aaf &  aae & ~aad & QAA ; 
assign FCA =  aaf &  aae &  aad & QAA ; 
assign FCI = ZZI ; 
assign HEE = ZZO & ~leb & ~lea & lec |  KAE & ~leb & lea & lec |  KBE & leb & ~lea & lec |  KCE & leb & lea & lec; 
assign hee = ~HEE;  //complement 
assign HFE = ZZO & ~lfb & ~lfa & lfc |         KAE & ~lfb & lfa & lfc |  KBE & lfb & ~lfa & lfc |  KCE & lfb & lfa & lfc; 
assign hfe = ~HFE;  //complement 
assign wee = ~WEE;  //complement 
assign wef = ~WEF;  //complement 
assign HEF = ZZO & ~leb & ~lea & lec |  KAF & ~leb & lea & lec |  KBF & leb & ~lea & lec |  KCF & leb & lea & lec; 
assign hef = ~HEF;  //complement 
assign HFF = ZZO & ~lfb & ~lfa & lfc |         KAF & ~lfb & lfa & lfc |  KBF & lfb & ~lfa & lfc |  KCF & lfb & lfa & lfc; 
assign hff = ~HFF;  //complement 
assign deo = ~DEO;  //complement 
assign tec = ~TEC;  //complement 
assign HEG = ZZO & ~leb & ~lea & lec |  KAG & ~leb & lea & lec |  KBG & leb & ~lea & lec |  KCG & leb & lea & lec; 
assign heg = ~HEG;  //complement 
assign HFG = ZZO & ~lfb & ~lfa & lfc |         KAG & ~lfb & lfa & lfc |  KBG & lfb & ~lfa & lfc |  KCG & lfb & lfa & lfc; 
assign hfg = ~HFG;  //complement 
assign dep = ~DEP;  //complement 
assign ted = ~TED;  //complement 
assign HEH = ZZO & ~leb & ~lea & lec |  KAH & ~leb & lea & lec |  KBH & leb & ~lea & lec |  KCH & leb & lea & lec; 
assign heh = ~HEH;  //complement 
assign HFH = ZZO & ~lfb & ~lfa & lfc |         KAH & ~lfb & lfa & lfc |  KBH & lfb & ~lfa & lfc |  KCH & lfb & lfa & lfc; 
assign hfh = ~HFH;  //complement 
assign weg = ~WEG;  //complement 
assign weh = ~WEH;  //complement 
assign tsa = ~TSA;  //complement 
assign tsb = ~TSB;  //complement 
assign tsc = ~TSC;  //complement 
assign tsd = ~TSD;  //complement 
assign DEI = ~dei;  //complement 
assign DEJ = ~dej;  //complement 
assign DEK = ~dek;  //complement 
assign DEL = ~del;  //complement 
assign tse = ~TSE;  //complement 
assign tsf = ~TSF;  //complement 
assign tsg = ~TSG;  //complement 
assign tsh = ~TSH;  //complement 
assign sae = ~SAE;  //complement 
assign saf = ~SAF;  //complement 
assign gae = ~GAE;  //complement 
assign gam = ~GAM;  //complement 
assign caa = ~CAA;  //complement 
assign cab = ~CAB;  //complement 
assign cac = ~CAC;  //complement 
assign FBA = ~CAC & ~CAB & ~CAA & CAD ; 
assign FBB = ~CAC & ~CAB &  CAA & CAD ; 
assign FBC = ~CAC &  CAB & ~CAA & CAD ; 
assign FBD = ~CAC &  CAB &  CAA & CAD ; 
assign FBE =  CAC & ~CAB & ~CAA & CAD ; 
assign FBF =  CAC & ~CAB &  CAA & CAD ; 
assign FBG =  CAC &  CAB & ~CAA & CAD ; 
assign FBH =  CAC &  CAB &  CAA & CAD ; 
assign FBI = ZZI ; 
assign sbe = ~SBE;  //complement 
assign sbf = ~SBF;  //complement 
assign MAE =  SJE & SKE & QDA  |  SJE & ske & QDB  |  sje & SKE & QDC  ; 
assign mae = ~MAE; //complement 
assign ABA = ~aba;  //complement 
assign ABB = ~abb;  //complement 
assign ABC = ~abc;  //complement 
assign FAA = ~AAC & ~AAB & ~AAA & ZZI ; 
assign FAB = ~AAC & ~AAB &  AAA & ZZI ; 
assign FAC = ~AAC &  AAB & ~AAA & ZZI ; 
assign FAD = ~AAC &  AAB &  AAA & ZZI ; 
assign FAE =  AAC & ~AAB & ~AAA & ZZI ; 
assign FAF =  AAC & ~AAB &  AAA & ZZI ; 
assign FAG =  AAC &  AAB & ~AAA & ZZI ; 
assign FAH =  AAC &  AAB &  AAA & ZZI ; 
assign FAI = ZZI ; 
assign JAE =  SAE & NAC  |  SBE & NBC  |  SCE & NCC  |  SDE & NDC  ; 
assign jae = ~JAE;  //complement 
assign JAM =  SAE & NAC  |  SBE & NBC  |  SCE & NCC  |  SDE & NDC  ; 
assign jam = ~JAM; //complement 
assign nac = ~NAC;  //complement 
assign ncc = ~NCC;  //complement 
assign sje = ~SJE;  //complement 
assign qaa = ~QAA;  //complement 
assign qab = ~QAB;  //complement 
assign qac = ~QAC;  //complement 
assign aaa = ~AAA;  //complement 
assign aab = ~AAB;  //complement 
assign aac = ~AAC;  //complement 
assign JAF =  SAF & NAC  |  SBF & NBC  |  SCF & NCC  |  SDF & NDC  ; 
assign jaf = ~JAF;  //complement 
assign JAN =  SAF & NAC  |  SBF & NBC  |  SCF & NCC  |  SDF & NDC  ; 
assign jan = ~JAN; //complement 
assign deg = ~DEG;  //complement 
assign nbc = ~NBC;  //complement 
assign ndc = ~NDC;  //complement 
assign oqb = ~OQB;  //complement 
assign qba = ~QBA;  //complement 
assign eac =  ske & skf  ; 
assign EAC = ~eac;  //complement 
assign ead =  skg & skh  ; 
assign EAD = ~ead;  //complement 
assign eae =  skh  ; 
assign EAE = ~eae;  //complement 
assign scf = ~SCF;  //complement 
assign sce = ~SCE;  //complement 
assign OAE = ~oae;  //complement 
assign OBE = ~obe;  //complement 
assign OCE = ~oce;  //complement 
assign SKE = ~ske;  //complement 
assign aad = ~AAD;  //complement 
assign aae = ~AAE;  //complement 
assign aaf = ~AAF;  //complement 
assign aag = ~AAG;  //complement 
assign FEA = ~AAF & ~AAE & ~AAD & QAB ; 
assign FEB = ~AAF & ~AAE &  AAD & QAB ; 
assign FEC = ~AAF &  AAE & ~AAD & QAB ; 
assign FED = ~AAF &  AAE &  AAD & QAB ; 
assign FEE =  AAF & ~AAE & ~AAD & QAB ; 
assign FEF =  AAF & ~AAE &  AAD & QAB ; 
assign FEG =  AAF &  AAE & ~AAD & QAB ; 
assign FEH =  AAF &  AAE &  AAD & QAB ; 
assign FEI = ZZI ; 
assign sde = ~SDE;  //complement 
assign sdf = ~SDF;  //complement 
assign gbe = ~GBE;  //complement 
assign gbm = ~GBM;  //complement 
assign bad = ~BAD;  //complement 
assign bae = ~BAE;  //complement 
assign baf = ~BAF;  //complement 
assign FDA = ~AAF & ~AAE & ~AAD & QBA ; 
assign FDB = ~AAF & ~AAE &  AAD & QBA ; 
assign FDC = ~AAF &  AAE & ~AAD & QBA ; 
assign FDD = ~AAF &  AAE &  AAD & QBA ; 
assign FDE =  AAF & ~AAE & ~AAD & QBA ; 
assign FDF =  AAF & ~AAE &  AAD & QBA ; 
assign FDG =  AAF &  AAE & ~AAD & QBA ; 
assign FDH =  AAF &  AAE &  AAD & QBA ; 
assign FDI = ZZI ;
assign fda = ~FDA;
assign fdb = ~FDB;
assign fdc = ~FDC;
assign fdd = ~FDD;
assign fde = ~FDE;
assign fdf = ~FDF;
assign fdg = ~FDG;
assign fdh = ~FDH;
   
assign lea = ~LEA;  //complement 
assign leb = ~LEB;  //complement 
assign lec = ~LEC;  //complement 
assign dec = ~DEC;  //complement 
assign ded = ~DED;  //complement 
assign dee = ~DEE;  //complement 
assign def = ~DEF;  //complement 
assign ufa = ~UFA;  //complement 
assign ufb = ~UFB;  //complement 
assign ufc = ~UFC;  //complement 
assign vfa = ~VFA;  //complement 
assign vfi = ~VFI;  //complement 
assign hla = vai & ~llb & ~lla & llc |  vbi & ~llb & lla & llc |  vci & llb & ~lla & llc |  vdi & llb & lla & llc; 
assign HLA = ~hla;  //complement 
assign hra = vai & ~lrb & ~lra & lrc |         vbi & ~lrb & lra & lrc |  vci & lrb & ~lra & lrc |  vdi & lrb & lra & lrc; 
assign HRA = ~hra;  //complement 
assign ufd = ~UFD;  //complement 
assign ufe = ~UFE;  //complement 
assign uff = ~UFF;  //complement 
assign vfb = ~VFB;  //complement 
assign vfj = ~VFJ;  //complement 
assign hlb = vaj & ~llb & ~lla & llc |  vbj & ~llb & lla & llc |  vcj & llb & ~lla & llc |  vdj & llb & lla & llc; 
assign HLB = ~hlb;  //complement 
assign hrb = vaj & ~lrb & ~lra & lrc |         vbj & ~lrb & lra & lrc |  vcj & lrb & ~lra & lrc |  vdj & lrb & lra & lrc; 
assign HRB = ~hrb;  //complement 
assign ufg = ~UFG;  //complement 
assign ufh = ~UFH;  //complement 
assign ufi = ~UFI;  //complement 
assign vfc = ~VFC;  //complement 
assign vfk = ~VFK;  //complement 
assign hlc = vak & ~llb & ~lla & llc |  vbk & ~llb & lla & llc |  vck & llb & ~lla & llc |  vdk & llb & lla & llc; 
assign HLC = ~hlc;  //complement 
assign hrc = vak & ~lrb & ~lra & lrc |         vbk & ~lrb & lra & lrc |  vck & lrb & ~lra & lrc |  vdk & lrb & lra & lrc; 
assign HRC = ~hrc;  //complement 
assign ufj = ~UFJ;  //complement 
assign ufk = ~UFK;  //complement 
assign ufl = ~UFL;  //complement 
assign vfd = ~VFD;  //complement 
assign vfl = ~VFL;  //complement 
assign hld = val & ~llb & ~lla & llc |  vbl & ~llb & lla & llc |  vcl & llb & ~lla & llc |  vdl & llb & lla & llc; 
assign HLD = ~hld;  //complement 
assign hrd = val & ~lrb & ~lra & lrc |         vbl & ~lrb & lra & lrc |  vcl & lrb & ~lra & lrc |  vdl & lrb & lra & lrc; 
assign HRD = ~hrd;  //complement 
assign ufm = ~UFM;  //complement 
assign ufn = ~UFN;  //complement 
assign ufo = ~UFO;  //complement 
assign vfe = ~VFE;  //complement 
assign vfm = ~VFM;  //complement 
assign hle = vam & ~llb & ~lla & llc |  vbm & ~llb & lla & llc |  vcm & llb & ~lla & llc |  vdm & llb & lla & llc; 
assign HLE = ~hle;  //complement 
assign hre = vam & ~lrb & ~lra & lrc |         vbm & ~lrb & lra & lrc |  vcm & lrb & ~lra & lrc |  vdm & lrb & lra & lrc; 
assign HRE = ~hre;  //complement 
assign ufp = ~UFP;  //complement 
assign ufq = ~UFQ;  //complement 
assign ufr = ~UFR;  //complement 
assign vff = ~VFF;  //complement 
assign vfn = ~VFN;  //complement 
assign hlf = van & ~llb & ~lla & llc |  vbn & ~llb & lla & llc |  vcn & llb & ~lla & llc |  vdn & llb & lla & llc; 
assign HLF = ~hlf;  //complement 
assign hrf = van & ~lrb & ~lra & lrc |         vbn & ~lrb & lra & lrc |  vcn & lrb & ~lra & lrc |  vdn & lrb & lra & lrc; 
assign HRF = ~hrf;  //complement 
assign uft = ~UFT;  //complement 
assign ufu = ~UFU;  //complement 
assign ufs = ~UFS;  //complement 
assign vfg = ~VFG;  //complement 
assign vfo = ~VFO;  //complement 
assign hlg = vao & ~llb & ~lla & llc |  vbo & ~llb & lla & llc |  vco & llb & ~lla & llc |  vdo & llb & lla & llc; 
assign HLG = ~hlg;  //complement 
assign hrg = vao & ~lrb & ~lra & lrc |         vbo & ~lrb & lra & lrc |  vco & lrb & ~lra & lrc |  vdo & lrb & lra & lrc; 
assign HRG = ~hrg;  //complement 
assign ufv = ~UFV;  //complement 
assign ufw = ~UFW;  //complement 
assign ufx = ~UFX;  //complement 
assign vfh = ~VFH;  //complement 
assign vfp = ~VFP;  //complement 
assign hlh = vap & ~llb & ~lla & llc |  vbp & ~llb & lla & llc |  vcp & llb & ~lla & llc |  vdp & llb & lla & llc; 
assign HLH = ~hlh;  //complement 
assign hrh = vap & ~lrb & ~lra & lrc |         vbp & ~lrb & lra & lrc |  vcp & lrb & ~lra & lrc |  vdp & lrb & lra & lrc; 
assign HRH = ~hrh;  //complement 
assign hli = vhi & ~LLB & ~LLA & LLC |  vgi & ~LLB & LLA & LLC |  vfi & LLB & ~LLA & LLC |  vei & LLB & LLA & LLC; 
assign HLI = ~hli;  //complement 
assign hri = vhi & ~LRB & ~LRA & LRC |         vgi & ~LRB & LRA & LRC |  vfi & LRB & ~LRA & LRC |  vei & LRB & LRA & LRC; 
assign HRI = ~hri;  //complement 
assign HEI = ZZO & ~LEB & ~LEA & LEC |  KFA & ~LEB & LEA & LEC |  KEA & LEB & ~LEA & LEC |  KDA & LEB & LEA & LEC; 
assign hei = ~HEI;  //complement 
assign HFI = ZZO & ~LFB & ~LFA & LFC |         KFA & ~LFB & LFA & LFC |  KEA & LFB & ~LFA & LFC |  KDA & LFB & LFA & LFC; 
assign hfi = ~HFI;  //complement 
assign wfa = ~WFA;  //complement 
assign wfb = ~WFB;  //complement 
assign hlj = vhj & ~LLB & ~LLA & LLC |  vgj & ~LLB & LLA & LLC |  vfj & LLB & ~LLA & LLC |  vej & LLB & LLA & LLC; 
assign HLJ = ~hlj;  //complement 
assign hrj = vhj & ~LRB & ~LRA & LRC |         vgj & ~LRB & LRA & LRC |  vfj & LRB & ~LRA & LRC |  vej & LRB & LRA & LRC; 
assign HRJ = ~hrj;  //complement 
assign HEJ = ZZO & ~LEB & ~LEA & LEC |  KFB & ~LEB & LEA & LEC |  KEB & LEB & ~LEA & LEC |  KDB & LEB & LEA & LEC; 
assign hej = ~HEJ;  //complement 
assign HFJ = ZZO & ~LFB & ~LFA & LFC |         KFB & ~LFB & LFA & LFC |  KEB & LFB & ~LFA & LFC |  KDB & LFB & LFA & LFC; 
assign hfj = ~HFJ;  //complement 
assign dfm = ~DFM;  //complement 
assign dfn = ~DFN;  //complement 
assign tfa = ~TFA;  //complement 
assign tfb = ~TFB;  //complement 
assign hlk = vhk & ~LLB & ~LLA & LLC |  vgk & ~LLB & LLA & LLC |  vfk & LLB & ~LLA & LLC |  vek & LLB & LLA & LLC; 
assign HLK = ~hlk;  //complement 
assign hrk = vhk & ~LRB & ~LRA & LRC |         vgk & ~LRB & LRA & LRC |  vfk & LRB & ~LRA & LRC |  vek & LRB & LRA & LRC; 
assign HRK = ~hrk;  //complement 
assign HEK = ZZO & ~LEB & ~LEA & LEC |  KFC & ~LEB & LEA & LEC |  KEC & LEB & ~LEA & LEC |  KDC & LEB & LEA & LEC; 
assign hek = ~HEK;  //complement 
assign HFK = ZZO & ~LFB & ~LFA & LFC |         KFC & ~LFB & LFA & LFC |  KEC & LFB & ~LFA & LFC |  KDC & LFB & LFA & LFC; 
assign hfk = ~HFK;  //complement 
assign KDA = ~kda;  //complement 
assign KDB = ~kdb;  //complement 
assign KDC = ~kdc;  //complement 
assign KDD = ~kdd;  //complement 
assign hll = vhl & ~LLB & ~LLA & LLC |  vgl & ~LLB & LLA & LLC |  vfl & LLB & ~LLA & LLC |  vel & LLB & LLA & LLC; 
assign HLL = ~hll;  //complement 
assign hrl = vhl & ~LRB & ~LRA & LRC |         vgl & ~LRB & LRA & LRC |  vfl & LRB & ~LRA & LRC |  vel & LRB & LRA & LRC; 
assign HRL = ~hrl;  //complement 
assign lla = ~LLA;  //complement 
assign llb = ~LLB;  //complement 
assign llc = ~LLC;  //complement 
assign HEL = ZZO & ~LEB & ~LEA & LEC |  KFD & ~LEB & LEA & LEC |  KED & LEB & ~LEA & LEC |  KDD & LEB & LEA & LEC; 
assign hel = ~HEL;  //complement 
assign HFL = ZZO & ~LFB & ~LFA & LFC |         KFD & ~LFB & LFA & LFC |  KED & LFB & ~LFA & LFC |  KDD & LFB & LFA & LFC; 
assign hfl = ~HFL;  //complement 
assign wfc = ~WFC;  //complement 
assign wfd = ~WFD;  //complement 
assign hlm = vhm & ~LLB & ~LLA & LLC |  vgm & ~LLB & LLA & LLC |  vfm & LLB & ~LLA & LLC |  vem & LLB & LLA & LLC; 
assign HLM = ~hlm;  //complement 
assign hrm = vhm & ~LRB & ~LRA & LRC |         vgm & ~LRB & LRA & LRC |  vfm & LRB & ~LRA & LRC |  vem & LRB & LRA & LRC; 
assign HRM = ~hrm;  //complement 
assign lra = ~LRA;  //complement 
assign lrb = ~LRB;  //complement 
assign lrc = ~LRC;  //complement 
assign HEM = ZZO & ~LEB & ~LEA & LEC |  KFE & ~LEB & LEA & LEC |  KEE & LEB & ~LEA & LEC |  KDE & LEB & LEA & LEC; 
assign hem = ~HEM;  //complement 
assign HFM = ZZO & ~LFB & ~LFA & LFC |         KFE & ~LFB & LFA & LFC |  KEE & LFB & ~LFA & LFC |  KDE & LFB & LFA & LFC; 
assign hfm = ~HFM;  //complement 
assign wfe = ~WFE;  //complement 
assign wff = ~WFF;  //complement 
assign hln = vhn & ~LLB & ~LLA & LLC |  vgn & ~LLB & LLA & LLC |  vfn & LLB & ~LLA & LLC |  ven & LLB & LLA & LLC; 
assign HLN = ~hln;  //complement 
assign hrn = vhn & ~LRB & ~LRA & LRC |         vgn & ~LRB & LRA & LRC |  vfn & LRB & ~LRA & LRC |  ven & LRB & LRA & LRC; 
assign HRN = ~hrn;  //complement 
assign HEN = ZZO & ~LEB & ~LEA & LEC |  KFF & ~LEB & LEA & LEC |  KEF & LEB & ~LEA & LEC |  KDF & LEB & LEA & LEC; 
assign hen = ~HEN;  //complement 
assign HFN = ZZO & ~LFB & ~LFA & LFC |         KFF & ~LFB & LFA & LFC |  KEF & LFB & ~LFA & LFC |  KDF & LFB & LFA & LFC; 
assign hfn = ~HFN;  //complement 
assign dfo = ~DFO;  //complement 
assign dfp = ~DFP;  //complement 
assign tfc = ~TFC;  //complement 
assign tfd = ~TFD;  //complement 
assign hlo = vho & ~LLB & ~LLA & LLC |  vgo & ~LLB & LLA & LLC |  vfo & LLB & ~LLA & LLC |  veo & LLB & LLA & LLC; 
assign HLO = ~hlo;  //complement 
assign hro = vho & ~LRB & ~LRA & LRC |         vgo & ~LRB & LRA & LRC |  vfo & LRB & ~LRA & LRC |  veo & LRB & LRA & LRC; 
assign HRO = ~hro;  //complement 
assign HEO = ZZO & ~LEB & ~LEA & LEC |  KFG & ~LEB & LEA & LEC |  KEG & LEB & ~LEA & LEC |  KDG & LEB & LEA & LEC; 
assign heo = ~HEO;  //complement 
assign HFO = ZZO & ~LFB & ~LFA & LFC |         KFG & ~LFB & LFA & LFC |  KEG & LFB & ~LFA & LFC |  KDG & LFB & LFA & LFC; 
assign hfo = ~HFO;  //complement 
assign KDE = ~kde;  //complement 
assign KDF = ~kdf;  //complement 
assign KDG = ~kdg;  //complement 
assign KDH = ~kdh;  //complement 
assign hlp = vhp & ~LLB & ~LLA & LLC |  vgp & ~LLB & LLA & LLC |  vfp & LLB & ~LLA & LLC |  vep & LLB & LLA & LLC; 
assign HLP = ~hlp;  //complement 
assign hrp = vhp & ~LRB & ~LRA & LRC |         vgp & ~LRB & LRA & LRC |  vfp & LRB & ~LRA & LRC |  vep & LRB & LRA & LRC; 
assign HRP = ~hrp;  //complement 
assign HEP = ZZO & ~LEB & ~LEA & LEC |  KFH & ~LEB & LEA & LEC |  KEH & LEB & ~LEA & LEC |  KDH & LEB & LEA & LEC; 
assign hep = ~HEP;  //complement 
assign HFP = ZZO & ~LFB & ~LFA & LFC |         KFH & ~LFB & LFA & LFC |  KEH & LFB & ~LFA & LFC |  KDH & LFB & LFA & LFC; 
assign hfp = ~HFP;  //complement 
assign wfg = ~WFG;  //complement 
assign wfh = ~WFH;  //complement 
assign oia = ~OIA;  //complement 
assign oja = ~OJA;  //complement 
assign DFI = ~dfi;  //complement 
assign DFJ = ~dfj;  //complement 
assign DFK = ~dfk;  //complement 
assign DFL = ~dfl;  //complement 
assign oib = ~OIB;  //complement 
assign ojb = ~OJB;  //complement 
assign see = ~SEE;  //complement 
assign sef = ~SEF;  //complement 
assign gaf = ~GAF;  //complement 
assign gan = ~GAN;  //complement 
assign oic = ~OIC;  //complement 
assign ojc = ~OJC;  //complement 
assign sfe = ~SFE;  //complement 
assign sff = ~SFF;  //complement 
assign MAF =  SJF & SKF & QDA  |  SJF & skf & QDB  |  sjf & SKF & QDC  ; 
assign maf = ~MAF; //complement 
assign oid = ~OID;  //complement 
assign ojd = ~OJD;  //complement 
assign JBE =  SEE & NEC  |  SFE & NFC  |  SGE & NGC  |  SHE & NHC  ; 
assign jbe = ~JBE;  //complement 
assign JBM =  SEE & NEC  |  SFE & NFC  |  SGE & NGC  |  SHE & NHC  ; 
assign jbm = ~JBM; //complement 
assign nec = ~NEC;  //complement 
assign ngc = ~NGC;  //complement 
assign sjf = ~SJF;  //complement 
assign oie = ~OIE;  //complement 
assign oje = ~OJE;  //complement 
assign JBF =  SEF & NEC  |  SFF & NFC  |  SGF & NGC  |  SHF & NHC  ; 
assign jbf = ~JBF;  //complement 
assign JBN =  SEF & NEC  |  SFF & NFC  |  SGF & NGC  |  SHF & NHC  ; 
assign jbn = ~JBN; //complement 
assign dfg = ~DFG;  //complement 
assign nfc = ~NFC;  //complement 
assign nhc = ~NHC;  //complement 
assign oif = ~OIF;  //complement 
assign ojf = ~OJF;  //complement 
assign sge = ~SGE;  //complement 
assign sgf = ~SGF;  //complement 
assign OAF = ~oaf;  //complement 
assign OBF = ~obf;  //complement 
assign OCF = ~ocf;  //complement 
assign SKF = ~skf;  //complement 
assign oig = ~OIG;  //complement 
assign ojg = ~OJG;  //complement 
assign she = ~SHE;  //complement 
assign shf = ~SHF;  //complement 
assign gbf = ~GBF;  //complement 
assign gbn = ~GBN;  //complement 
assign oih = ~OIH;  //complement 
assign ojh = ~OJH;  //complement 
assign lfa = ~LFA;  //complement 
assign lfb = ~LFB;  //complement 
assign lfc = ~LFC;  //complement 
assign dfc = ~DFC;  //complement 
assign dfd = ~DFD;  //complement 
assign dfe = ~DFE;  //complement 
assign dff = ~DFF;  //complement 
assign uga = ~UGA;  //complement 
assign ugb = ~UGB;  //complement 
assign ugc = ~UGC;  //complement 
assign vga = ~VGA;  //complement 
assign vgi = ~VGI;  //complement 
assign hsa = vai & ~lsb & ~lsa & lsc |  vbi & ~lsb & lsa & lsc |  vci & lsb & ~lsa & lsc |  vdi & lsb & lsa & lsc; 
assign HSA = ~hsa;  //complement 
assign ugd = ~UGD;  //complement 
assign uge = ~UGE;  //complement 
assign ugf = ~UGF;  //complement 
assign vgb = ~VGB;  //complement 
assign vgj = ~VGJ;  //complement 
assign ugg = ~UGG;  //complement 
assign ugh = ~UGH;  //complement 
assign ugi = ~UGI;  //complement 
assign vgg = ~VGG;  //complement 
assign vgo = ~VGO;  //complement 
assign vgc = ~VGC;  //complement 
assign vgk = ~VGK;  //complement 
assign hsc = vak & ~lsb & ~lsa & lsc |  vbk & ~lsb & lsa & lsc |  vck & lsb & ~lsa & lsc |  vdk & lsb & lsa & lsc; 
assign HSC = ~hsc;  //complement 
assign ugj = ~UGJ;  //complement 
assign ugk = ~UGK;  //complement 
assign ugl = ~UGL;  //complement 
assign vgd = ~VGD;  //complement 
assign vgl = ~VGL;  //complement 
assign hsd = val & ~lsb & ~lsa & lsc |  vbl & ~lsb & lsa & lsc |  vcl & lsb & ~lsa & lsc |  vdl & lsb & lsa & lsc; 
assign HSD = ~hsd;  //complement 
assign htd = val & ~ltb & ~lta & ltc |         vbl & ~ltb & lta & ltc |  vcl & ltb & ~lta & ltc |  vdl & ltb & lta & ltc; 
assign HTD = ~htd;  //complement 
assign ugm = ~UGM;  //complement 
assign ugn = ~UGN;  //complement 
assign ugo = ~UGO;  //complement 
assign vge = ~VGE;  //complement 
assign vgm = ~VGM;  //complement 
assign hte = vam & ~ltb & ~lta & ltc |  vbm & ~ltb & lta & ltc |  vcm & ltb & ~lta & ltc |  vdm & ltb & lta & ltc; 
assign HTE = ~hte;  //complement 
assign hse = vam & ~lsb & ~lsa & lsc |         vbm & ~lsb & lsa & lsc |  vcm & lsb & ~lsa & lsc |  vdm & lsb & lsa & lsc; 
assign HSE = ~hse;  //complement 
assign ugp = ~UGP;  //complement 
assign ugq = ~UGQ;  //complement 
assign ugr = ~UGR;  //complement 
assign vgf = ~VGF;  //complement 
assign vgn = ~VGN;  //complement 
assign hsf = van & ~lsb & ~lsa & lsc |  vbn & ~lsb & lsa & lsc |  vcn & lsb & ~lsa & lsc |  vdn & lsb & lsa & lsc; 
assign HSF = ~hsf;  //complement 
assign htf = van & ~ltb & ~lta & ltc |         vbn & ~ltb & lta & ltc |  vcn & ltb & ~lta & ltc |  vdn & ltb & lta & ltc; 
assign HTF = ~htf;  //complement 
assign ugs = ~UGS;  //complement 
assign ugt = ~UGT;  //complement 
assign ugu = ~UGU;  //complement 
assign hsb = vaj & ~lsb & ~lsa & lsc |  vbj & ~lsb & lsa & lsc |  vcj & lsb & ~lsa & lsc |  vdj & lsb & lsa & lsc; 
assign HSB = ~hsb;  //complement 
assign htb = vaj & ~ltb & ~lta & ltc |         vbj & ~ltb & lta & ltc |  vcj & ltb & ~lta & ltc |  vdj & ltb & lta & ltc; 
assign HTB = ~htb;  //complement 
assign ugv = ~UGV;  //complement 
assign ugw = ~UGW;  //complement 
assign ugx = ~UGX;  //complement 
assign vgh = ~VGH;  //complement 
assign vgp = ~VGP;  //complement 
assign hsh = vap & ~lsb & ~lsa & lsc |  vbp & ~lsb & lsa & lsc |  vcp & lsb & ~lsa & lsc |  vdp & lsb & lsa & lsc; 
assign HSH = ~hsh;  //complement 
assign hth = vap & ~ltb & ~lta & ltc |         vbp & ~ltb & lta & ltc |  vcp & ltb & ~lta & ltc |  vdp & ltb & lta & ltc; 
assign HTH = ~hth;  //complement 
assign hti = vhi & ~LTB & ~LTA & LTC |  vgi & ~LTB & LTA & LTC |  vfi & LTB & ~LTA & LTC |  vei & LTB & LTA & LTC; 
assign HTI = ~hti;  //complement 
assign hsi = vhi & ~LSB & ~LSA & LSC |         vgi & ~LSB & LSA & LSC |  vfi & LSB & ~LSA & LSC |  vei & LSB & LSA & LSC; 
assign HSI = ~hsi;  //complement 
assign HGA = ZZO & ~lgb & ~lga & lgc |  KAA & ~lgb & lga & lgc |  KBA & lgb & ~lga & lgc |  KCA & lgb & lga & lgc; 
assign hga = ~HGA;  //complement 
assign HHA = ZZO & ~lhb & ~lha & lhc |         KAA & ~lhb & lha & lhc |  KBA & lhb & ~lha & lhc |  KCA & lhb & lha & lhc; 
assign hha = ~HHA;  //complement 
assign wga = ~WGA;  //complement 
assign wgb = ~WGB;  //complement 
assign hsj = vhj & ~LSB & ~LSA & LSC |  vgj & ~LSB & LSA & LSC |  vfj & LSB & ~LSA & LSC |  vej & LSB & LSA & LSC; 
assign HSJ = ~hsj;  //complement 
assign HGB = ZZO & ~lgb & ~lga & lgc |  KAB & ~lgb & lga & lgc |  KBB & lgb & ~lga & lgc |  KCB & lgb & lga & lgc; 
assign hgb = ~HGB;  //complement 
assign HHB = ZZO & ~lhb & ~lha & lhc |         KAB & ~lhb & lha & lhc |  KBB & lhb & ~lha & lhc |  KCB & lhb & lha & lhc; 
assign hhb = ~HHB;  //complement 
assign dgm = ~DGM;  //complement 
assign dgn = ~DGN;  //complement 
assign tga = ~TGA;  //complement 
assign tgb = ~TGB;  //complement 
assign hsk = vhk & ~LSB & ~LSA & LSC |  vgk & ~LSB & LSA & LSC |  vfk & LSB & ~LSA & LSC |  vek & LSB & LSA & LSC; 
assign HSK = ~hsk;  //complement 
assign htk = vhk & ~LTB & ~LTA & LTC |         vgk & ~LTB & LTA & LTC |  vfk & LTB & ~LTA & LTC |  vek & LTB & LTA & LTC; 
assign HTK = ~htk;  //complement 
assign HGG = ZZO & ~lgb & ~lga & lgc |  KAG & ~lgb & lga & lgc |  KBG & lgb & ~lga & lgc |  KCG & lgb & lga & lgc; 
assign hgg = ~HGG;  //complement 
assign HHG = ZZO & ~lhb & ~lha & lhc |         KAG & ~lhb & lha & lhc |  KBG & lhb & ~lha & lhc |  KCG & lhb & lha & lhc; 
assign hhg = ~HHG;  //complement 
assign HGC = ZZO & ~lgb & ~lga & lgc |  KAC & ~lgb & lga & lgc |  KBC & lgb & ~lga & lgc |  KCC & lgb & lga & lgc; 
assign hgc = ~HGC;  //complement 
assign HHC = ZZO & ~lhb & ~lha & lhc |         KAC & ~lhb & lha & lhc |  KBC & lhb & ~lha & lhc |  KCC & lhb & lha & lhc; 
assign hhc = ~HHC;  //complement 
assign KEA = ~kea;  //complement 
assign KEB = ~keb;  //complement 
assign KEC = ~kec;  //complement 
assign KED = ~ked;  //complement 
assign hsl = vhl & ~LSB & ~LSA & LSC |  vgl & ~LSB & LSA & LSC |  vfl & LSB & ~LSA & LSC |  vel & LSB & LSA & LSC; 
assign HSL = ~hsl;  //complement 
assign lma = ~LMA;  //complement 
assign lmb = ~LMB;  //complement 
assign lmc = ~LMC;  //complement 
assign HGD = ZZO & ~lgb & ~lga & lgc |  KAD & ~lgb & lga & lgc |  KBD & lgb & ~lga & lgc |  KCD & lgb & lga & lgc; 
assign hgd = ~HGD;  //complement 
assign HHD = ZZO & ~lhb & ~lha & lhc |         KAD & ~lhb & lha & lhc |  KBD & lhb & ~lha & lhc |  KCD & lhb & lha & lhc; 
assign hhd = ~HHD;  //complement 
assign wgc = ~WGC;  //complement 
assign wgd = ~WGD;  //complement 
assign tib = ~TIB;  //complement 
assign tic = ~TIC;  //complement 
assign tid = ~TID;  //complement 
assign lsa = ~LSA;  //complement 
assign lsb = ~LSB;  //complement 
assign lsc = ~LSC;  //complement 
assign HGE = ZZO & ~lgb & ~lga & lgc |  KAE & ~lgb & lga & lgc |  KBE & lgb & ~lga & lgc |  KCE & lgb & lga & lgc; 
assign hge = ~HGE;  //complement 
assign HHE = ZZO & ~lhb & ~lha & lhc |         KAE & ~lhb & lha & lhc |  KBE & lhb & ~lha & lhc |  KCE & lhb & lha & lhc; 
assign hhe = ~HHE;  //complement 
assign wge = ~WGE;  //complement 
assign wgf = ~WGF;  //complement 
assign hsn = vhn & ~LSB & ~LSA & LSC |  vgn & ~LSB & LSA & LSC |  vfn & LSB & ~LSA & LSC |  ven & LSB & LSA & LSC; 
assign HSN = ~hsn;  //complement 
assign htn = vhn & ~LTB & ~LTA & LTC |         vgn & ~LTB & LTA & LTC |  vfn & LTB & ~LTA & LTC |  ven & LTB & LTA & LTC; 
assign HTN = ~htn;  //complement 
assign HGP = ZZO & ~LGB & ~LGA & LGC |  KFH & ~LGB & LGA & LGC |  KEH & LGB & ~LGA & LGC |  KDH & LGB & LGA & LGC; 
assign hgp = ~HGP;  //complement 
assign HHP = ZZO & ~LHB & ~LHA & LHC |         KFH & ~LHB & LHA & LHC |  KEH & LHB & ~LHA & LHC |  KDH & LHB & LHA & LHC; 
assign hhp = ~HHP;  //complement 
assign HGF = ZZO & ~lgb & ~lga & lgc |  KAF & ~lgb & lga & lgc |  KBF & lgb & ~lga & lgc |  KCF & lgb & lga & lgc; 
assign hgf = ~HGF;  //complement 
assign HHF = ZZO & ~lhb & ~lha & lhc |         KAF & ~lhb & lha & lhc |  KBF & lhb & ~lha & lhc |  KCF & lhb & lha & lhc; 
assign hhf = ~HHF;  //complement 
assign dgo = ~DGO;  //complement 
assign dgp = ~DGP;  //complement 
assign tgc = ~TGC;  //complement 
assign tgd = ~TGD;  //complement 
assign hso = vho & ~LSB & ~LSA & LSC |  vgo & ~LSB & LSA & LSC |  vfo & LSB & ~LSA & LSC |  veo & LSB & LSA & LSC; 
assign HSO = ~hso;  //complement 
assign KEE = ~kee;  //complement 
assign KEF = ~kef;  //complement 
assign KEG = ~keg;  //complement 
assign KEH = ~keh;  //complement 
assign hsp = vhp & ~LSB & ~LSA & LSC |  vgp & ~LSB & LSA & LSC |  vfp & LSB & ~LSA & LSC |  vep & LSB & LSA & LSC; 
assign HSP = ~hsp;  //complement 
assign htp = vhp & ~LTB & ~LTA & LTC |         vgp & ~LTB & LTA & LTC |  vfp & LTB & ~LTA & LTC |  vep & LTB & LTA & LTC; 
assign HTP = ~htp;  //complement 
assign HGH = ZZO & ~lgb & ~lga & lgc |  KAH & ~lgb & lga & lgc |  KBH & lgb & ~lga & lgc |  KCH & lgb & lga & lgc; 
assign hgh = ~HGH;  //complement 
assign HHH = ZZO & ~lhb & ~lha & lhc |         KAH & ~lhb & lha & lhc |  KBH & lhb & ~lha & lhc |  KCH & lhb & lha & lhc; 
assign hhh = ~HHH;  //complement 
assign wgg = ~WGG;  //complement 
assign wgh = ~WGH;  //complement 
assign oka = ~OKA;  //complement 
assign ola = ~OLA;  //complement 
assign DGI = ~dgi;  //complement 
assign DGJ = ~dgj;  //complement 
assign DGK = ~dgk;  //complement 
assign DGL = ~dgl;  //complement 
assign okb = ~OKB;  //complement 
assign olb = ~OLB;  //complement 
assign sag = ~SAG;  //complement 
assign sah = ~SAH;  //complement 
assign gag = ~GAG;  //complement 
assign gao = ~GAO;  //complement 
assign okc = ~OKC;  //complement 
assign olc = ~OLC;  //complement 
assign sbg = ~SBG;  //complement 
assign sbh = ~SBH;  //complement 
assign MAG =  SJG & SKG & QDA  |  SJG & skg & QDB  |  sjg & SKG & QDC  ; 
assign mag = ~MAG; //complement 
assign okd = ~OKD;  //complement 
assign old = ~OLD;  //complement 
assign JAG =  SAG & NAD  |  SBG & NBD  |  SCG & NCD  |  SDG & NDD  ; 
assign jag = ~JAG;  //complement 
assign JAO =  SAG & NAD  |  SBG & NBD  |  SCG & NCD  |  SDG & NDD  ; 
assign jao = ~JAO; //complement 
assign nad = ~NAD;  //complement 
assign ncd = ~NCD;  //complement 
assign sjg = ~SJG;  //complement 
assign oke = ~OKE;  //complement 
assign ole = ~OLE;  //complement 
assign JAH =  SAH & NAD  |  SBH & NBD  |  SCH & NCD  |  SDH & NDD  ; 
assign jah = ~JAH;  //complement 
assign JAP =  SAH & NAD  |  SBH & NBD  |  SCH & NCD  |  SDH & NDD  ; 
assign jap = ~JAP; //complement 
assign dgg = ~DGG;  //complement 
assign nbd = ~NBD;  //complement 
assign ndd = ~NDD;  //complement 
assign okf = ~OKF;  //complement 
assign olf = ~OLF;  //complement 
assign scg = ~SCG;  //complement 
assign sch = ~SCH;  //complement 
assign OAG = ~oag;  //complement 
assign OBG = ~obg;  //complement 
assign OCG = ~ocg;  //complement 
assign SKG = ~skg;  //complement 
assign okg = ~OKG;  //complement 
assign olg = ~OLG;  //complement 
assign sdg = ~SDG;  //complement 
assign sdh = ~SDH;  //complement 
assign gbg = ~GBG;  //complement 
assign gbo = ~GBO;  //complement 
assign okh = ~OKH;  //complement 
assign olh = ~OLH;  //complement 
assign lga = ~LGA;  //complement 
assign lgb = ~LGB;  //complement 
assign lgc = ~LGC;  //complement 
assign dgc = ~DGC;  //complement 
assign dgd = ~DGD;  //complement 
assign dge = ~DGE;  //complement 
assign dgf = ~DGF;  //complement 
assign uha = ~UHA;  //complement 
assign uhb = ~UHB;  //complement 
assign uhc = ~UHC;  //complement 
assign vha = ~VHA;  //complement 
assign vhi = ~VHI;  //complement 
assign hma = vai & ~lmb & ~lma & lmc |  vbi & ~lmb & lma & lmc |  vci & lmb & ~lma & lmc |  vdi & lmb & lma & lmc; 
assign HMA = ~hma;  //complement 
assign hna = vai & ~lnb & ~lna & lnc |         vbi & ~lnb & lna & lnc |  vci & lnb & ~lna & lnc |  vdi & lnb & lna & lnc; 
assign HNA = ~hna;  //complement 
assign uhd = ~UHD;  //complement 
assign uhe = ~UHE;  //complement 
assign uhf = ~UHF;  //complement 
assign vhb = ~VHB;  //complement 
assign vhj = ~VHJ;  //complement 
assign hmb = vaj & ~lmb & ~lma & lmc |  vbj & ~lmb & lma & lmc |  vcj & lmb & ~lma & lmc |  vdj & lmb & lma & lmc; 
assign HMB = ~hmb;  //complement 
assign hnb = vaj & ~lnb & ~lna & lnc |         vbj & ~lnb & lna & lnc |  vcj & lnb & ~lna & lnc |  vdj & lnb & lna & lnc; 
assign HNB = ~hnb;  //complement 
assign uhg = ~UHG;  //complement 
assign uhh = ~UHH;  //complement 
assign uhi = ~UHI;  //complement 
assign vhc = ~VHC;  //complement 
assign vhk = ~VHK;  //complement 
assign hmc = vak & ~lmb & ~lma & lmc |  vbk & ~lmb & lma & lmc |  vck & lmb & ~lma & lmc |  vdk & lmb & lma & lmc; 
assign HMC = ~hmc;  //complement 
assign hnc = vak & ~lnb & ~lna & lnc |         vbk & ~lnb & lna & lnc |  vck & lnb & ~lna & lnc |  vdk & lnb & lna & lnc; 
assign HNC = ~hnc;  //complement 
assign uhj = ~UHJ;  //complement 
assign uhk = ~UHK;  //complement 
assign uhl = ~UHL;  //complement 
assign vhd = ~VHD;  //complement 
assign vhl = ~VHL;  //complement 
assign hmd = val & ~lmb & ~lma & lmc |  vbl & ~lmb & lma & lmc |  vcl & lmb & ~lma & lmc |  vdl & lmb & lma & lmc; 
assign HMD = ~hmd;  //complement 
assign hnd = val & ~lnb & ~lna & lnc |         vbl & ~lnb & lna & lnc |  vcl & lnb & ~lna & lnc |  vdl & lnb & lna & lnc; 
assign HND = ~hnd;  //complement 
assign uhm = ~UHM;  //complement 
assign uhn = ~UHN;  //complement 
assign vhe = ~VHE;  //complement 
assign vhm = ~VHM;  //complement 
assign hme = vam & ~lmb & ~lma & lmc |  vbm & ~lmb & lma & lmc |  vcm & lmb & ~lma & lmc |  vdm & lmb & lma & lmc; 
assign HME = ~hme;  //complement 
assign hne = vam & ~lnb & ~lna & lnc |         vbm & ~lnb & lna & lnc |  vcm & lnb & ~lna & lnc |  vdm & lnb & lna & lnc; 
assign HNE = ~hne;  //complement 
assign uho = ~UHO;  //complement 
assign uhp = ~UHP;  //complement 
assign vhn = ~VHN;  //complement 
assign vhf = ~VHF;  //complement 
assign hmf = van & ~lmb & ~lma & lmc |  vbn & ~lmb & lma & lmc |  vcn & lmb & ~lma & lmc |  vdn & lmb & lma & lmc; 
assign HMF = ~hmf;  //complement 
assign hnf = van & ~lnb & ~lna & lnc |         vbn & ~lnb & lna & lnc |  vcn & lnb & ~lna & lnc |  vdn & lnb & lna & lnc; 
assign HNF = ~hnf;  //complement 
assign uhs = ~UHS;  //complement 
assign uht = ~UHT;  //complement 
assign uhu = ~UHU;  //complement 
assign vhg = ~VHG;  //complement 
assign vho = ~VHO;  //complement 
assign hmg = vao & ~lmb & ~lma & lmc |  vbo & ~lmb & lma & lmc |  vco & lmb & ~lma & lmc |  vdo & lmb & lma & lmc; 
assign HMG = ~hmg;  //complement 
assign hng = vao & ~lnb & ~lna & lnc |         vbo & ~lnb & lna & lnc |  vco & lnb & ~lna & lnc |  vdo & lnb & lna & lnc; 
assign HNG = ~hng;  //complement 
assign uhv = ~UHV;  //complement 
assign uhw = ~UHW;  //complement 
assign uhx = ~UHX;  //complement 
assign vhh = ~VHH;  //complement 
assign vhp = ~VHP;  //complement 
assign hmh = vap & ~lmb & ~lma & lmc |  vbp & ~lmb & lma & lmc |  vcp & lmb & ~lma & lmc |  vdp & lmb & lma & lmc; 
assign HMH = ~hmh;  //complement 
assign hnh = vap & ~lnb & ~lna & lnc |         vbp & ~lnb & lna & lnc |  vcp & lnb & ~lna & lnc |  vdp & lnb & lna & lnc; 
assign HNH = ~hnh;  //complement 
assign hmi = vhi & ~LMB & ~LMA & LMC |  vgi & ~LMB & LMA & LMC |  vfi & LMB & ~LMA & LMC |  vei & LMB & LMA & LMC; 
assign HMI = ~hmi;  //complement 
assign hni = vhi & ~LNB & ~LNA & LNC |         vgi & ~LNB & LNA & LNC |  vfi & LNB & ~LNA & LNC |  vei & LNB & LNA & LNC; 
assign HNI = ~hni;  //complement 
assign HGI = ZZO & ~LGB & ~LGA & LGC |  KFA & ~LGB & LGA & LGC |  KEA & LGB & ~LGA & LGC |  KDA & LGB & LGA & LGC; 
assign hgi = ~HGI;  //complement 
assign HHI = ZZO & ~LHB & ~LHA & LHC |         KFA & ~LHB & LHA & LHC |  KEA & LHB & ~LHA & LHC |  KDA & LHB & LHA & LHC; 
assign hhi = ~HHI;  //complement 
assign wha = ~WHA;  //complement 
assign whb = ~WHB;  //complement 
assign htj = vhj & ~LTB & ~LTA & LTC |  vgj & ~LTB & LTA & LTC |  vfj & LTB & ~LTA & LTC |  vej & LTB & LTA & LTC; 
assign HTJ = ~htj;  //complement 
assign HGN = ZZO & ~LGB & ~LGA & LGC |  KFF & ~LGB & LGA & LGC |  KEF & LGB & ~LGA & LGC |  KDF & LGB & LGA & LGC; 
assign hgn = ~HGN;  //complement 
assign HHN = ZZO & ~LHB & ~LHA & LHC |         KFF & ~LHB & LHA & LHC |  KEF & LHB & ~LHA & LHC |  KDF & LHB & LHA & LHC; 
assign hhn = ~HHN;  //complement 
assign HGJ = ZZO & ~LGB & ~LGA & LGC |  KFB & ~LGB & LGA & LGC |  KEB & LGB & ~LGA & LGC |  KDB & LGB & LGA & LGC; 
assign hgj = ~HGJ;  //complement 
assign HHJ = ZZO & ~LHB & ~LHA & LHC |         KFB & ~LHB & LHA & LHC |  KEB & LHB & ~LHA & LHC |  KDB & LHB & LHA & LHC; 
assign hhj = ~HHJ;  //complement 
assign dhm = ~DHM;  //complement 
assign dhn = ~DHN;  //complement 
assign tha = ~THA;  //complement 
assign thb = ~THB;  //complement 
assign htl = vhl & ~LTB & ~LTA & LTC |  vgl & ~LTB & LTA & LTC |  vfl & LTB & ~LTA & LTC |  vel & LTB & LTA & LTC; 
assign HTL = ~htl;  //complement 
assign hta = vai & ~ltb & ~lta & ltc |  vbi & ~ltb & lta & ltc |  vci & ltb & ~lta & ltc |  vdi & ltb & lta & ltc; 
assign HTA = ~hta;  //complement 
assign HGK = ZZO & ~LGB & ~LGA & LGC |  KFC & ~LGB & LGA & LGC |  KEC & LGB & ~LGA & LGC |  KDC & LGB & LGA & LGC; 
assign hgk = ~HGK;  //complement 
assign HHK = ZZO & ~LHB & ~LHA & LHC |         KFC & ~LHB & LHA & LHC |  KEC & LHB & ~LHA & LHC |  KDC & LHB & LHA & LHC; 
assign hhk = ~HHK;  //complement 
assign KFA = ~kfa;  //complement 
assign KFB = ~kfb;  //complement 
assign KFC = ~kfc;  //complement 
assign KFD = ~kfd;  //complement 
assign htg = vao & ~ltb & ~lta & ltc |  vbo & ~ltb & lta & ltc |  vco & ltb & ~lta & ltc |  vdo & ltb & lta & ltc; 
assign HTG = ~htg;  //complement 
assign hsg = vao & ~lsb & ~lsa & lsc |         vbo & ~lsb & lsa & lsc |  vco & lsb & ~lsa & lsc |  vdo & lsb & lsa & lsc; 
assign HSG = ~hsg;  //complement 
assign lna = ~LNA;  //complement 
assign lnb = ~LNB;  //complement 
assign lnc = ~LNC;  //complement 
assign HGL = ZZO & ~LGB & ~LGA & LGC |  KFD & ~LGB & LGA & LGC |  KED & LGB & ~LGA & LGC |  KDD & LGB & LGA & LGC; 
assign hgl = ~HGL;  //complement 
assign HHL = ZZO & ~LHB & ~LHA & LHC |         KFD & ~LHB & LHA & LHC |  KED & LHB & ~LHA & LHC |  KDD & LHB & LHA & LHC; 
assign hhl = ~HHL;  //complement 
assign whc = ~WHC;  //complement 
assign whd = ~WHD;  //complement 
assign KFE = ~kfe;  //complement 
assign KFF = ~kff;  //complement 
assign KFG = ~kfg;  //complement 
assign KFH = ~kfh;  //complement 
assign lta = ~LTA;  //complement 
assign ltb = ~LTB;  //complement 
assign ltc = ~LTC;  //complement 
assign whe = ~WHE;  //complement 
assign whf = ~WHF;  //complement 
assign hmn = vhn & ~LMB & ~LMA & LMC |  vgn & ~LMB & LMA & LMC |  vfn & LMB & ~LMA & LMC |  ven & LMB & LMA & LMC; 
assign HMN = ~hmn;  //complement 
assign hnn = vhn & ~LNB & ~LNA & LNC |         vgn & ~LNB & LNA & LNC |  vfn & LNB & ~LNA & LNC |  ven & LNB & LNA & LNC; 
assign HNN = ~hnn;  //complement 
assign htm = vhm & ~LTB & ~LTA & LTC |  vgm & ~LTB & LTA & LTC |  vfm & LTB & ~LTA & LTC |  vem & LTB & LTA & LTC; 
assign HTM = ~htm;  //complement 
assign hsm = vhm & ~LSB & ~LSA & LSC |         vgm & ~LSB & LSA & LSC |  vfm & LSB & ~LSA & LSC |  vem & LSB & LSA & LSC; 
assign HSM = ~hsm;  //complement 
assign dho = ~DHO;  //complement 
assign dhp = ~DHP;  //complement 
assign thd = ~THD;  //complement 
assign thc = ~THC;  //complement 
assign hmo = vho & ~LMB & ~LMA & LMC |  vgo & ~LMB & LMA & LMC |  vfo & LMB & ~LMA & LMC |  veo & LMB & LMA & LMC; 
assign HMO = ~hmo;  //complement 
assign hno = vho & ~LNB & ~LNA & LNC |         vgo & ~LNB & LNA & LNC |  vfo & LNB & ~LNA & LNC |  veo & LNB & LNA & LNC; 
assign HNO = ~hno;  //complement 
assign hto = vho & ~LTB & ~LTA & LTC |  vgo & ~LTB & LTA & LTC |  vfo & LTB & ~LTA & LTC |  veo & LTB & LTA & LTC; 
assign HTO = ~hto;  //complement 
assign uhq = ~UHQ;  //complement 
assign uhr = ~UHR;  //complement 
assign hmp = vhp & ~LMB & ~LMA & LMC |  vgp & ~LMB & LMA & LMC |  vfp & LMB & ~LMA & LMC |  vep & LMB & LMA & LMC; 
assign HMP = ~hmp;  //complement 
assign hnp = vhp & ~LNB & ~LNA & LNC |         vgp & ~LNB & LNA & LNC |  vfp & LNB & ~LNA & LNC |  vep & LNB & LNA & LNC; 
assign HNP = ~hnp;  //complement 
assign htc = vak & ~ltb & ~lta & ltc |  vbk & ~ltb & lta & ltc |  vck & ltb & ~lta & ltc |  vdk & ltb & lta & ltc; 
assign HTC = ~htc;  //complement 
assign HGO = ZZO & ~LGB & ~LGA & LGC |  KFG & ~LGB & LGA & LGC |  KEG & LGB & ~LGA & LGC |  KDG & LGB & LGA & LGC; 
assign hgo = ~HGO;  //complement 
assign HHO = ZZO & ~LHB & ~LHA & LHC |         KFG & ~LHB & LHA & LHC |  KEG & LHB & ~LHA & LHC |  KDG & LHB & LHA & LHC; 
assign hho = ~HHO;  //complement 
assign whg = ~WHG;  //complement 
assign whh = ~WHH;  //complement 
assign oga = ~OGA;  //complement 
assign oha = ~OHA;  //complement 
assign DHI = ~dhi;  //complement 
assign DHJ = ~dhj;  //complement 
assign DHK = ~dhk;  //complement 
assign DHL = ~dhl;  //complement 
assign ogb = ~OGB;  //complement 
assign ohb = ~OHB;  //complement 
assign seg = ~SEG;  //complement 
assign seh = ~SEH;  //complement 
assign gah = ~GAH;  //complement 
assign gap = ~GAP;  //complement 
assign ogc = ~OGC;  //complement 
assign ohc = ~OHC;  //complement 
assign sfg = ~SFG;  //complement 
assign sfh = ~SFH;  //complement 
assign MAH =  SJH & SKH & QDA  |  SJH & skh & QDB  |  sjh & SKH & QDC  ; 
assign mah = ~MAH; //complement 
assign ogd = ~OGD;  //complement 
assign ohd = ~OHD;  //complement 
assign JBG =  SEG & NED  |  SFG & NFD  |  SGG & NGD  |  SHG & NHD  ; 
assign jbg = ~JBG;  //complement 
assign JBO =  SEG & NED  |  SFG & NFD  |  SGG & NGD  |  SHG & NHD  ; 
assign jbo = ~JBO; //complement 
assign ned = ~NED;  //complement 
assign ngd = ~NGD;  //complement 
assign sjh = ~SJH;  //complement 
assign oge = ~OGE;  //complement 
assign ohe = ~OHE;  //complement 
assign JBH =  SEH & NED  |  SFH & NFD  |  SGH & NGD  |  SHH & NHD  ; 
assign jbh = ~JBH;  //complement 
assign JBP =  SEH & NED  |  SFH & NFD  |  SGH & NGD  |  SHH & NHD  ; 
assign jbp = ~JBP; //complement 
assign dhg = ~DHG;  //complement 
assign nfd = ~NFD;  //complement 
assign nhd = ~NHD;  //complement 
assign ogf = ~OGF;  //complement 
assign ohf = ~OHF;  //complement 
assign sgg = ~SGG;  //complement 
assign sgh = ~SGH;  //complement 
assign OAH = ~oah;  //complement 
assign OBH = ~obh;  //complement 
assign OCH = ~och;  //complement 
assign SKH = ~skh;  //complement 
assign ogg = ~OGG;  //complement 
assign ohg = ~OHG;  //complement 
assign shg = ~SHG;  //complement 
assign shh = ~SHH;  //complement 
assign gbh = ~GBH;  //complement 
assign gbp = ~GBP;  //complement 
assign ogh = ~OGH;  //complement 
assign ohh = ~OHH;  //complement 
assign lha = ~LHA;  //complement 
assign lhb = ~LHB;  //complement 
assign lhc = ~LHC;  //complement 
assign dhc = ~DHC;  //complement 
assign dhd = ~DHD;  //complement 
assign dhe = ~DHE;  //complement 
assign dhf = ~DHF;  //complement 
assign iaa = ~IAA; //complement 
assign iab = ~IAB; //complement 
assign iac = ~IAC; //complement 
assign iad = ~IAD; //complement 
assign iae = ~IAE; //complement 
assign iaf = ~IAF; //complement 
assign iag = ~IAG; //complement 
assign iah = ~IAH; //complement 
assign iba = ~IBA; //complement 
assign ibb = ~IBB; //complement 
assign ibc = ~IBC; //complement 
assign ibd = ~IBD; //complement 
assign ibe = ~IBE; //complement 
assign ibf = ~IBF; //complement 
assign ibg = ~IBG; //complement 
assign ibh = ~IBH; //complement 
assign ica = ~ICA; //complement 
assign icb = ~ICB; //complement 
assign icc = ~ICC; //complement 
assign icd = ~ICD; //complement 
assign ice = ~ICE; //complement 
assign icf = ~ICF; //complement 
assign icg = ~ICG; //complement 
assign ich = ~ICH; //complement 
assign ida = ~IDA; //complement 
assign idb = ~IDB; //complement 
assign idc = ~IDC; //complement 
assign idd = ~IDD; //complement 
assign ide = ~IDE; //complement 
assign idf = ~IDF; //complement 
assign idg = ~IDG; //complement 
assign idh = ~IDH; //complement 
assign iea = ~IEA; //complement 
assign ieb = ~IEB; //complement 
assign iec = ~IEC; //complement 
assign ied = ~IED; //complement 
assign iee = ~IEE; //complement 
assign ief = ~IEF; //complement 
assign ieg = ~IEG; //complement 
assign ieh = ~IEH; //complement 
assign ifa = ~IFA; //complement 
assign ifb = ~IFB; //complement 
assign ifc = ~IFC; //complement 
assign ifd = ~IFD; //complement 
assign ife = ~IFE; //complement 
assign ifff  = ~IFFF ; //complement 
assign ifg = ~IFG; //complement 
assign ifh = ~IFH; //complement 
assign iga = ~IGA; //complement 
assign igb = ~IGB; //complement 
assign igc = ~IGC; //complement 
assign igd = ~IGD; //complement 
assign ige = ~IGE; //complement 
assign igf = ~IGF; //complement 
assign igg = ~IGG; //complement 
assign igh = ~IGH; //complement 
assign iha = ~IHA; //complement 
assign ihb = ~IHB; //complement 
assign ihc = ~IHC; //complement 
assign ihd = ~IHD; //complement 
assign ihe = ~IHE; //complement 
assign ihf = ~IHF; //complement 
assign ihg = ~IHG; //complement 
assign ihh = ~IHH; //complement 
assign iia = ~IIA; //complement 
assign iib = ~IIB; //complement 
assign iic = ~IIC; //complement 
assign iid = ~IID; //complement 
assign iie = ~IIE; //complement 
assign iif = ~IIF; //complement 
assign iig = ~IIG; //complement 
assign iih = ~IIH; //complement 
assign ija = ~IJA; //complement 
assign ijb = ~IJB; //complement 
assign ijc = ~IJC; //complement 
assign ijd = ~IJD; //complement 
assign ije = ~IJE; //complement 
assign ijf = ~IJF; //complement 
assign ijg = ~IJG; //complement 
assign ijh = ~IJH; //complement 
assign ika = ~IKA; //complement 
assign ikb = ~IKB; //complement 
assign ikc = ~IKC; //complement 
assign ikd = ~IKD; //complement 
assign ike = ~IKE; //complement 
assign ikf = ~IKF; //complement 
assign ikg = ~IKG; //complement 
assign ikh = ~IKH; //complement 
assign ima = ~IMA; //complement 
assign imb = ~IMB; //complement 
assign imc = ~IMC; //complement 
assign imd = ~IMD; //complement 
assign ime = ~IME; //complement 
assign imf = ~IMF; //complement 
assign img = ~IMG; //complement 
assign imh = ~IMH; //complement 
assign ina = ~INA; //complement 
assign inb = ~INB; //complement 
assign inc = ~INC; //complement 
assign ind = ~IND; //complement 
assign ine = ~INE; //complement 
assign inf = ~INF; //complement 
assign ing = ~ING; //complement 
assign inh = ~INH; //complement 
assign ioa = ~IOA; //complement 
assign iob = ~IOB; //complement 
assign ioc = ~IOC; //complement 
assign iod = ~IOD; //complement 
assign ioe = ~IOE; //complement 
assign iof = ~IOF; //complement 
assign iog = ~IOG; //complement 
assign ioh = ~IOH; //complement 
assign ipa = ~IPA; //complement 
assign ipb = ~IPB; //complement 
assign ipc = ~IPC; //complement 
assign ipd = ~IPD; //complement 
assign ipe = ~IPE; //complement 
assign ipf = ~IPF; //complement 
assign ipg = ~IPG; //complement 
assign iph = ~IPH; //complement 
assign iqa = ~IQA; //complement 
assign iqb = ~IQB; //complement 
assign iqc = ~IQC; //complement 
assign iqd = ~IQD; //complement 
assign iqe = ~IQE; //complement 
assign iqf = ~IQF; //complement 
assign iqg = ~IQG; //complement 
assign iqh = ~IQH; //complement 
assign ira = ~IRA; //complement 
assign irb = ~IRB; //complement 
assign irc = ~IRC; //complement 
assign ird = ~IRD; //complement 
assign ire = ~IRE; //complement 
assign irf = ~IRF; //complement 
assign irg = ~IRG; //complement 
assign irh = ~IRH; //complement 
assign isa = ~ISA; //complement 
assign isb = ~ISB; //complement 
assign isc = ~ISC; //complement 
assign isd = ~ISD; //complement 
assign ise = ~ISE; //complement 
assign isf = ~ISF; //complement 
assign isg = ~ISG; //complement 
assign ita = ~ITA; //complement 
assign itb = ~ITB; //complement 
assign itc = ~ITC; //complement 
assign itd = ~ITD; //complement 
assign ite = ~ITE; //complement 
assign itf = ~ITF; //complement 
always@(posedge IZZ )
   begin 
 UAA <= DAG & DAI |  ZZO & dai ; 
 UAB <= UAA & DAI |  UAA & dai ; 
 UAC <= DAC & DAI |  UAC & dai ; 
 VAA <=  RAA & TAA  |  RAI & TAB  |  RIA & TAC  |  RII & TAD  ; 
 VAI <=  RAA & TAA  |  RAI & TAB  |  RIA & TAC  |  RII & TAD  ; 
 UAD <= DAD & DAI |  UAD & dai ; 
 UAE <= DAE & DAI |  UAE & dai ; 
 UAF <= DAF & DAI |  UAF & dai ; 
 VAB <=  RAB & TAA  |  RAJ & TAB  |  RIB & TAC  |  RIJ & TAD  ; 
 VAJ <=  RAB & TAA  |  RAJ & TAB  |  RIB & TAC  |  RIJ & TAD  ; 
 UAG <= DAG & DAJ |  ZZO & daj ; 
 UAH <= UAG & DAJ |  UAG & daj ; 
 UAI <= DAC & DAJ |  UAI & daj ; 
 VAC <=  RAC & TAA  |  RAK & TAB  |  RIC & TAC  |  RIK & TAD  ; 
 VAK <=  RAC & TAA  |  RAK & TAB  |  RIC & TAC  |  RIK & TAD  ; 
 UAJ <= DAD & DAJ |  UAJ & daj ; 
 UAK <= DAE & DAJ |  UAK & daj ; 
 UAL <= DAF & DAJ |  UAL & daj ; 
 VAD <=  RAD & TAA  |  RAL & TAB  |  RID & TAC  |  RIL & TAD  ; 
 VAL <=  RAD & TAA  |  RAL & TAB  |  RID & TAC  |  RIL & TAD  ; 
 UAM <= DAG & DAK |  ZZO & dak ; 
 UAN <= UAM & DAK |  UAM & dak ; 
 UAO <= DAC & DAK |  UAO & dak ; 
 VAE <=  RAE & TAA  |  RAM & TAB  |  RIE & TAC  |  RIM & TAD  ; 
 VAM <=  RAE & TAA  |  RAM & TAB  |  RIE & TAC  |  RIM & TAD  ; 
 UAP <= DAD & DAK |  UAP & dak ; 
 UAQ <= DAE & DAK |  UAQ & dak ; 
 UAR <= DAF & DAK |  UAR & dak ; 
 VAF <=  RAF & TAA  |  RAN & TAB  |  RIF & TAC  |  RIN & TAD  ; 
 VAN <=  RAF & TAA  |  RAN & TAB  |  RIF & TAC  |  RIN & TAD  ; 
 UAT <= UAS & DAL |  UAS & dal ; 
 UAU <= DAC & DAL |  UAU & dal ; 
 UAS <= DAG & DAL |  ZZO & dal ; 
 VAG <=  RAG & TAA  |  RAO & TAB  |  RIG & TAC  |  RIO & TAD  ; 
 VAO <=  RAG & TAA  |  RAO & TAB  |  RIG & TAC  |  RIO & TAD  ; 
 UAV <= DAD & DAL |  UAV & dal ; 
 UAW <= DAE & DAL |  UAW & dal ; 
 UAX <= DAF & DAL |  UAX & dal ; 
 VAH <=  RAH & TAA  |  RAP & TAB  |  RIH & TAC  |  RIP & TAD  ; 
 VAP <=  RAH & TAA  |  RAP & TAB  |  RIH & TAC  |  RIP & TAD  ; 
 WAA <=  HAA  |  HAI  ; 
 WAB <=  HAB  |  HAJ  ; 
 DAM <= dag & DAI ; 
 DAN <= dag & DAJ ; 
 TAA <= dag & DAM ; 
 TAB <= dag & DAN ; 
 kaa <= ika ; 
 kab <= ikb ; 
 kac <= ikc ; 
 kad <= ikd ; 
 LIA <= BBA & BAJ |  LIA & baj ; 
 LIB <= BBB & BAJ |  LIB & baj ; 
 LIC <= BBC & BAJ |  LIC & baj ; 
 WAC <=  HAC  |  HAK  ; 
 WAD <=  HAD  |  HAL  ; 
 LOA <= ABA & BAJ |  LOA & baj ; 
 LOB <= ABB & BAJ |  LOB & baj ; 
 LOC <= ABC & BAJ |  LOC & baj ; 
 WAE <=  HAE  |  HAM  ; 
 WAF <=  HAF  |  HAN  ; 
 DAO <= dag & DAK ; 
 DAP <= dag & DAL ; 
 TAC <= dag & DAO ; 
 TAD <= dag & DAP ; 
 kae <= ike ; 
 kaf <= ikf ; 
 kag <= ikg ; 
 kah <= ikh ; 
 WAG <=  HAG  |  HAO  ; 
 WAH <=  HAH  |  HAP  ; 
 OFA <=  HIA & HII  ; 
 OEA <=  HOA & HOI & tjb  |  JAA & TJB  |  JBA & TKB  ; 
 dai <=  iah  |  IAB  |  IAA  ; 
 daj <=  iah  |  IAB  |  iaa  ; 
 dak <=  iah  |  iab  |  IAA  ; 
 dal <=  iah  |  iab  |  iaa  ; 
 OFB <=  HIB & HIJ  ; 
 OEB <=  HOB & HOJ & tjb  |  JAB & TJB  |  JBB & TKB  ; 
 SAA <=  GAA & TSA  |  GBA & TSA  |  SAA & tsa  ; 
 SAB <=  GAB & TSA  |  GBB & TSA  |  SAB & tsa  ; 
 GAA <=  IRA & CAE  |  IPA & CAF  |  IQA & CAG  |  MAA  ; 
 GAI <=  IRA & CAE  |  IPA & CAF  |  IQA & CAG  |  MAA  ; 
 OFC <=  HIC & HIK  ; 
 OEC <=  HOC & HOK & tjb  |  JAC & TJB  |  JBC & TKB  ; 
 SBA <=  GAA & TSB  |  GBA & TSB  |  SBA & tsb  ; 
 SBB <=  GAB & TSB  |  GBB & TSB  |  SBB & tsb  ; 
 OFD <=  HID & HIL  ; 
 OED <=  HOD & HOL & tjb  |  JAD & TJB  |  JBD & TKB  ; 
 NAA <= FAA ; 
 NCA <= FAC ; 
 QDA <= QCA ; 
 SJA <= SKA ; 
 OFE <=  HIE & HIM  ; 
 OEE <=  HOE & HOM & tjb  |  JAE & TJB  |  JBE & TKB  ; 
 DAG <= IAG ; 
 NBA <= FAB ; 
 NDA <= FAD ; 
 OFF <=  HIF & HIN  ; 
 OEF <=  HOF & HON & tjb  |  JAF & TJB  |  JBF & TKB  ; 
 SCA <=  GAA & TSC  |  GBA & TSC  |  SCA & tsc  ; 
 SCB <=  GAB & TSC  |  GBB & TSC  |  SCB & tsc  ; 
 oaa <= jba & jaa ; 
 oba <= jba & jaa ; 
 oca <= jba & jaa ; 
 ska <= jba & jaa ; 
 OFG <=  HIG & HIO  ; 
 OEG <=  HOG & HOO & tjb  |  JAG & TJB  |  JBG & TKB  ; 
 SDA <=  GAA & TSD  |  GBA & TSD  |  SDA & tsd  ; 
 SDB <=  GAB & TSD  |  GBB & TSD  |  SDB & tsd  ; 
 GBA <=  INA & CAH  |  IOA & CAI  |  IMA & CAJ  |  IIA  |  IJA  ; 
 GBI <=  INA & CAH  |  IOA & CAI  |  IMA & CAJ  |  IIA  |  IJA  ; 
 OFH <=  HIH & HIP  ; 
 OEH <=  HOH & HOP & tjb  |  JAH & TJB  |  JBH & TKB  ; 
 LAA <= BAD & FDA |  LAA & fda ; 
 LAB <= BAE & FDA |  LAB & fda ; 
 LAC <= BAF & FDA |  LAC & fda ; 
 DAC <= IAC ; 
 DAD <= IAD ; 
 DAE <= IAE ; 
 DAF <= IAF ; 
 UBA <= DBG & DBI |  ZZO & dbi ; 
 UBB <= UBA & DBI |  UBA & dbi ; 
 UBC <= DBC & DBI |  UBC & dbi ; 
 VBA <=  RBA & TBA  |  RBI & TBB  |  RJA & TBC  |  RJI & TBD  ; 
 VBI <=  RBA & TBA  |  RBI & TBB  |  RJA & TBC  |  RJI & TBD  ; 
 UBD <= DBD & DBI |  UBD & dbi ; 
 UBE <= DBE & DBI |  UBE & dbi ; 
 UBF <= DBF & DBI |  UBF & dbi ; 
 VBB <=  RBB & TBA  |  RBJ & TBB  |  RJB & TBC  |  RJJ & TBD  ; 
 VBJ <=  RBB & TBA  |  RBJ & TBB  |  RJB & TBC  |  RJJ & TBD  ; 
 UBG <= DBG & DBJ |  ZZO & dbj ; 
 UBH <= UBG & DBJ |  UBG & dbj ; 
 UBI <= DBC & DBJ |  UBI & dbj ; 
 VBC <=  RBC & TBA  |  RBK & TBB  |  RJC & TBC  |  RJK & TBD  ; 
 VBK <=  RBC & TBA  |  RBK & TBB  |  RJC & TBC  |  RJK & TBD  ; 
 UBJ <= DBD & DBJ |  UBJ & dbj ; 
 UBK <= DBE & DBJ |  UBK & dbj ; 
 UBL <= DBF & DBJ |  UBL & dbj ; 
 VBD <=  RBD & TBA  |  RBL & TBB  |  RJD & TBC  |  RJL & TBD  ; 
 VBL <=  RBD & TBA  |  RBL & TBB  |  RJD & TBC  |  RJL & TBD  ; 
 UBM <= DBG & DBK |  ZZO & dbk ; 
 UBN <= UBM & DBK |  UBM & dbk ; 
 UBO <= DBC & DBK |  UBO & dbk ; 
 VBE <=  RBE & TBA  |  RBM & TBB  |  RJE & TBC  |  RJM & TBD  ; 
 VBM <=  RBE & TBA  |  RBM & TBB  |  RJE & TBC  |  RJM & TBD  ; 
 UBP <= DBD & DBK |  UBP & dbk ; 
 UBQ <= DBE & DBK |  UBQ & dbk ; 
 UBR <= DBF & DBK |  UBR & dbk ; 
 VBN <=  RBF & TBA  |  RBN & TBB  |  RJF & TBC  |  RJN & TBD  ; 
 VBF <=  RBF & TBA  |  RBN & TBB  |  RJF & TBC  |  RJN & TBD  ; 
 UBS <= DBG & DBL |  ZZO & dbl ; 
 UBT <= UBS & DBL |  UBS & dbl ; 
 UBU <= DBC & DBL |  UBU & dbl ; 
 VBG <=  RBG & TBA  |  RBO & TBB  |  RJG & TBC  |  RJO & TBD  ; 
 VBO <=  RBG & TBA  |  RBO & TBB  |  RJG & TBC  |  RJO & TBD  ; 
 UBV <= DBD & DBL |  UBV & dbl ; 
 UBW <= DBE & DBL |  UBW & dbl ; 
 UBX <= DBF & DBL |  UBX & dbl ; 
 VBH <=  RBH & TBA  |  RBP & TBB  |  RJH & TBC  |  RJP & TBD  ; 
 VBP <=  RBH & TBA  |  RBP & TBB  |  RJH & TBC  |  RJP & TBD  ; 
 WBA <=  HBA  |  HBI  ; 
 WBB <=  HBB  |  HBJ  ; 
 DBM <= dbg & DBI ; 
 DBN <= dbg & DBJ ; 
 TBA <= dbg & DBM ; 
 TBB <= dbg & DBN ; 
 kba <= ipa ; 
 kbb <= ipb ; 
 kbc <= ipc ; 
 kbd <= ipd ; 
 LJA <= BBA & BAL |  LJA & bal ; 
 LJB <= BBB & BAL |  LJB & bal ; 
 LJC <= BBC & BAL |  LJC & bal ; 
 WBC <=  HBC  |  HBK  ; 
 WBD <=  HBD  |  HBL  ; 
 LPA <= ABA & BAL |  LPA & bal ; 
 LPB <= ABB & BAL |  LPB & bal ; 
 LPC <= ABC & BAL |  LPC & bal ; 
 WBE <=  HBE  |  HBM  ; 
 WBF <=  HBF  |  HBN  ; 
 DBO <= dbg & DBK ; 
 DBP <= dbg & DBL ; 
 TBC <= dbg & DBO ; 
 TBD <= dbg & DBP ; 
 kbe <= ipe ; 
 kbf <= ipf ; 
 kbg <= ipg ; 
 kbh <= iph ; 
 WBG <=  HBG  |  HBO  ; 
 WBH <=  HBH  |  HBP  ; 
 ONA <=  HJA & HJI  ; 
 OOA <=  HPA & HPI & tjd  |  JAA & TJD  |  JBA & TKD  ; 
 dbi <=  ibh  |  IBB  |  IBA  ; 
 dbj <=  ibh  |  IBB  |  iba  ; 
 dbk <=  ibh  |  ibb  |  IBA  ; 
 dbl <=  ibh  |  ibb  |  iba  ; 
 ONB <=  HJB & HJJ  ; 
 OOB <=  HPB & HPJ & tjd  |  JAB & TJD  |  JBB & TKD  ; 
 SEA <=  GAI & TSE  |  GBI & TSE  |  SEA & tse  ; 
 SEB <=  GAJ & TSE  |  GBJ & TSE  |  SEB & tse  ; 
 GAB <=  IRB & CAE  |  IPB & CAF  |  IQB & CAG  |  MAB  ; 
 GAJ <=  IRB & CAE  |  IPB & CAF  |  IQB & CAG  |  MAB  ; 
 ONC <=  HJC & HJK  ; 
 OOC <=  HPC & HPK & tjd  |  JAC & TJD  |  JBC & TKD  ; 
 SFA <=  GAI & TSF  |  GBI & TSF  |  SFA & tsf  ; 
 SFB <=  GAJ & TSF  |  GBJ & TSF  |  SFB & tsf  ; 
 OND <=  HJD & HJL  ; 
 OOD <=  HPD & HPL & tjd  |  JAD & TJD  |  JBD & TKD  ; 
 NEA <= FAE ; 
 NGA <= FAG ; 
 QDB <= QCB ; 
 SJB <= SKB ; 
 ONE <=  HJE & HJM  ; 
 OOE <=  HPE & HPM & tjd  |  JAE & TJD  |  JBE & TKD  ; 
 DBG <= IBG ; 
 NFA <= FAF ; 
 NHA <= FAH ; 
 ONF <=  HJF & HJN  ; 
 OOF <=  HPF & HPN & tjd  |  JAF & TJD  |  JBF & TKD  ; 
 SGA <=  GAI & TSG  |  GBI & TSG  |  SGA & tsg  ; 
 SGB <=  GAJ & TSG  |  GBJ & TSG  |  SGB & tsg  ; 
 oab <= jbb & jab ; 
 obb <= jbb & jab ; 
 ocb <= jbb & jab ; 
 skb <= jbb & jab ; 
 ONG <=  HJG & HJO  ; 
 OOG <=  HPG & HPO & tjd  |  JAG & TJD  |  JBG & TKD  ; 
 SHA <=  GAI & TSH  |  GBI & TSH  |  SHA & tsg  ; 
 SHB <=  GAJ & TSH  |  GBJ & TSH  |  SHB & tsg  ; 
 GBB <=  INB & CAH  |  IOB & CAI  |  IMB & CAJ  |  IIB  |  IJB  ; 
 GBJ <=  INB & CAH  |  IOB & CAI  |  IMB & CAJ  |  IIB  |  IJB  ; 
 ONH <=  HJH & HJP  ; 
 OOH <=  HPH & HPP & tjd  |  JAH & TJD  |  JBH & TKD  ; 
 LBA <= BAD & FDB |  LBA & fdb ; 
 LBB <= BAE & FDB |  LBB & fdb ; 
 LBC <= BAF & FDB |  LBC & fdb ; 
 DBC <= IBC ; 
 DBD <= IBD ; 
 DBE <= IBE ; 
 DBF <= IBF ; 
 UCA <= DCG & DCI |  ZZO & dci ; 
 UCB <= UCA & DCI |  UCA & dci ; 
 UCC <= DCC & DCI |  UCC & dci ; 
 VCA <=  RCA & TCA  |  RCI & TCB  |  RKA & TCC  |  RKI & TCD  ; 
 VCI <=  RCA & TCA  |  RCI & TCB  |  RKA & TCC  |  RKI & TCD  ; 
 UCD <= DCD & DCI |  UCD & dci ; 
 UCE <= DCE & DCI |  UCE & dci ; 
 UCF <= DCF & DCI |  UCF & dci ; 
 VCB <=  RCB & TCA  |  RCJ & TCB  |  RKB & TCC  |  RKJ & TCD  ; 
 VCJ <=  RCB & TCA  |  RCJ & TCB  |  RKB & TCC  |  RKJ & TCD  ; 
 UCG <= DCG & DCJ |  ZZO & dcj ; 
 UCI <= DCC & DCJ |  UCI & dcj ; 
 UCH <= UCG & DCJ |  UCG & dcj ; 
 VCC <=  RCC & TCA  |  RCK & TCB  |  RKC & TCC  |  RKK & TCD  ; 
 VCK <=  RCC & TCA  |  RCK & TCB  |  RKC & TCC  |  RKK & TCD  ; 
 UCJ <= DCD & DCJ |  UCJ & dcj ; 
 UCK <= DCE & DCJ |  UCK & dcj ; 
 UCL <= DCF & DCJ |  UCL & dcj ; 
 VCD <=  RCD & TCA  |  RCL & TCB  |  RKD & TCC  |  RKL & TCD  ; 
 VCL <=  RCD & TCA  |  RCL & TCB  |  RKD & TCC  |  RKL & TCD  ; 
 UCM <= DCG & DCK |  ZZO & dck ; 
 UCN <= UCM & DCK |  UCM & dck ; 
 UCO <= DCC & DCK |  UCO & dck ; 
 VCE <=  RCE & TCA  |  RCM & TCB  |  RKE & TCC  |  RKM & TCD  ; 
 VCM <=  RCE & TCA  |  RCM & TCB  |  RKE & TCC  |  RKM & TCD  ; 
 UCP <= DCD & DCK |  UCP & dck ; 
 UCQ <= DCE & DCK |  UCQ & dck ; 
 UCR <= DCF & DCK |  UCR & dck ; 
 VCF <=  RCF & TCA  |  RCN & TCB  |  RKF & TCC  |  RKN & TCD  ; 
 VCN <=  RCF & TCA  |  RCN & TCB  |  RKF & TCC  |  RKN & TCD  ; 
 UCS <= DCG & DCL |  ZZO & dcl ; 
 UCT <= UCS & DCL |  UCS & dcl ; 
 UCU <= DCC & DCL |  UCU & dcl ; 
 VCH <=  RCH & TCA  |  RCP & TCB  |  RKH & TCC  |  RKP & TCD  ; 
 VCP <=  RCH & TCA  |  RCP & TCB  |  RKH & TCC  |  RKP & TCD  ; 
 UCV <= DCD & DCL |  UCV & dcl ; 
 UCW <= DCE & DCL |  UCW & dcl ; 
 UCX <= DCF & DCL |  UCX & dcl ; 
 VCG <=  RCG & TCA  |  RCO & TCB  |  RKG & TCC  |  RKO & TCD  ; 
 VCO <=  RCG & TCA  |  RCO & TCB  |  RKG & TCC  |  RKO & TCD  ; 
 DCM <= dcg & DCI ; 
 DCN <= dcg & DCJ ; 
 TCA <= dcg & DCM ; 
 TCB <= dcg & DCN ; 
 WCA <=  HCA  |  HCI  ; 
 WCB <=  HCB  |  HCJ  ; 
 kca <= iqa ; 
 kcb <= iqb ; 
 kcc <= iqc ; 
 kcd <= iqd ; 
 LKA <= BBA & BAJ |  LKA & baj ; 
 LKB <= BBB & BAJ |  LKB & baj ; 
 LKC <= BBC & BAJ |  LKC & baj ; 
 WCC <=  HCC  |  HCK  ; 
 WCD <=  HCD  |  HCL  ; 
 LQA <= ABA & BAK |  LQA & bak ; 
 LQB <= ABB & BAK |  LQB & bak ; 
 LQC <= ABC & BAK |  LQC & bak ; 
 WCE <=  HCE  |  HCM  ; 
 WCF <=  HCF  |  HCN  ; 
 DCO <= dcg & DCK ; 
 DCP <= dcg & DCL ; 
 TCC <= dcg & DCO ; 
 TCD <= dcg & DCP ; 
 kce <= iqe ; 
 kcf <= iqf ; 
 kcg <= iqg ; 
 kch <= iqh ; 
 WCG <=  HCG  |  HCO  ; 
 WCH <=  HCH  |  HCP  ; 
 ODA <=  HKA & HKI  ; 
 OMA <=  HQA & HQI & tjc  |  JAA & TJC  |  JBA & TKC  ; 
 dci <=  ich  |  ICB  |  ICA  ; 
 dcj <=  ich  |  ICB  |  ica  ; 
 dck <=  ich  |  icb  |  ICA  ; 
 dcl <=  ich  |  icb  |  ica  ; 
 ODB <=  HKB & HKJ  ; 
 OMB <=  HQB & HQJ & tjc  |  JAB & TJC  |  JBB & TKC  ; 
 SAC <=  GAC & TSA  |  GBC & TSA  |  SAC & tsa  ; 
 SAD <=  GAD & TSA  |  GBD & TSA  |  SAD & tsa  ; 
 GAC <=  IRC & CAE  |  IPC & CAF  |  IQC & CAG  |  MAC  ; 
 GAK <=  IRC & CAE  |  IPC & CAF  |  IQC & CAG  |  MAC  ; 
 ODC <=  HKC & HKK  ; 
 OMC <=  HQC & HQK & tjc  |  JAC & TJC  |  JBC & TKC  ; 
 SBC <=  GAC & TSB  |  GBC & TSB  |  SBC & tsb  ; 
 SBD <=  GAD & TSB  |  GBD & TSB  |  SBD & tsb  ; 
 ODD <=  HKD & HKL  ; 
 OMD <=  HQD & HQL & tjc  |  JAD & TJC  |  JBD & TKC  ; 
 NAB <= FAA ; 
 NCB <= FAC ; 
 QDC <= QCC ; 
 SJC <= SKC ; 
 ODE <=  HKE & HKM  ; 
 OME <=  HQE & HQM & tjc  |  JAE & TJC  |  JBE & TKC  ; 
 DCG <= ICG ; 
 NBB <= FAB ; 
 NDB <= FAD ; 
 ODF <=  HKF & HKN  ; 
 OMF <=  HQF & HQN & tjc  |  JAF & TJC  |  JBF & TKC  ; 
 SCC <=  GAC & TSC  |  GBC & TSC  |  SCC & tsc  ; 
 SCD <=  GAD & TSC  |  GBD & TSC  |  SCD & tsc  ; 
 oac <= jbc & jac ; 
 obc <= jbc & jac ; 
 occ <= jbc & jac ; 
 skc <= jbc & jac ; 
 ODG <=  HKG & HKO  ; 
 OMG <=  HQG & HQO & tjc  |  JAG & TJC  |  JBG & TKC  ; 
 SDC <=  GAC & TSD  |  GBC & TSD  |  SDC & tsd  ; 
 SDD <=  GAD & TSD  |  GBD & TSD  |  SDD & tsd  ; 
 GBC <=  INC & CAH  |  IOC & CAI  |  IMC & CAJ  |  IIC  |  IJC  ; 
 GBK <=  INC & CAH  |  IOC & CAI  |  IMC & CAJ  |  IIC  |  IJC  ; 
 ODH <=  HKH & HKP  ; 
 OMH <=  HQH & HQP & tjc  |  JAH & TJC  |  JBH & TKC  ; 
 LCA <= BAD & FDC |  LCA & fdc ; 
 LCB <= BAE & FDC |  LCB & fdc ; 
 LCC <= BAF & FDC |  LCC & fdc ; 
 DCC <= ICC ; 
 DCD <= ICD ; 
 DCE <= ICE ; 
 DCF <= ICF ; 
 UDA <= DDG & DDI |  ZZO & ddi ; 
 UDB <= UDA & DDI |  UDA & ddi ; 
 UDC <= DDC & DDI |  UDC & ddi ; 
 VDA <=  RDA & TDA  |  RDI & TDB  |  RLA & TDC  |  RLI & TDD  ; 
 VDI <=  RDA & TDA  |  RDI & TDB  |  RLA & TDC  |  RLI & TDD  ; 
 UDD <= DDD & DDI |  UDD & ddi ; 
 UDE <= DDE & DDI |  UDE & ddi ; 
 UDF <= DDF & DDI |  UDF & ddi ; 
 VDB <=  RDB & TDA  |  RDJ & TDB  |  RLB & TDC  |  RLJ & TDD  ; 
 VDJ <=  RDB & TDA  |  RDJ & TDB  |  RLB & TDC  |  RLJ & TDD  ; 
 UDG <= DDG & DDJ |  ZZO & ddj ; 
 UDH <= UDG & DDJ |  UDG & ddj ; 
 UDI <= DDC & DDJ |  UDI & ddj ; 
 VDC <=  RDC & TDA  |  RDK & TDB  |  RLC & TDC  |  RLK & TDD  ; 
 VDK <=  RDC & TDA  |  RDK & TDB  |  RLC & TDC  |  RLK & TDD  ; 
 UDJ <= DDD & DDJ |  UDJ & ddj ; 
 UDK <= DDE & DDJ |  UDK & ddj ; 
 UDL <= DDF & DDJ |  UDL & ddj ; 
 VDD <=  RDD & TDA  |  RDL & TDB  |  RLD & TDC  |  RLL & TDD  ; 
 VDL <=  RDD & TDA  |  RDL & TDB  |  RLD & TDC  |  RLL & TDD  ; 
 UDM <= DDG & DDK |  ZZO & ddk ; 
 UDN <= UDM & DDK |  UDM & ddk ; 
 UDO <= DDC & DDK |  UDO & ddk ; 
 VDE <=  RDE & TDA  |  RDM & TDB  |  RLE & TDC  |  RLM & TDD  ; 
 VDM <=  RDE & TDA  |  RDM & TDB  |  RLE & TDC  |  RLM & TDD  ; 
 UDP <= DDD & DDK |  UDP & ddk ; 
 UDQ <= DDE & DDK |  UDQ & ddk ; 
 UDR <= DDF & DDK |  UDR & ddk ; 
 VDF <=  RDF & TDA  |  RDN & TDB  |  RLF & TDC  |  RLN & TDD  ; 
 VDN <=  RDF & TDA  |  RDN & TDB  |  RLF & TDC  |  RLN & TDD  ; 
 UDS <= DDG & DDL |  ZZO & ddl ; 
 UDT <= UDS & DDL |  UDS & ddl ; 
 UDU <= DDC & DDL |  UDU & ddl ; 
 VDG <=  RDG & TDA  |  RDO & TDB  |  RLG & TDC  |  RLO & TDD  ; 
 VDO <=  RDG & TDA  |  RDO & TDB  |  RLG & TDC  |  RLO & TDD  ; 
 UDV <= DDD & DDL |  UDV & ddl ; 
 UDW <= DDE & DDL |  UDW & ddl ; 
 UDX <= DDF & DDL |  UDX & ddl ; 
 VDH <=  RDH & TDA  |  RDP & TDB  |  RLH & TDC  |  RLP & TDD  ; 
 VDP <=  RDH & TDA  |  RDP & TDB  |  RLH & TDC  |  RLP & TDD  ; 
 WDA <=  HDA  |  HDI  ; 
 WDB <=  HDB  |  HDJ  ; 
 DDM <= ddg & DDI ; 
 TDA <= ddg & DDM ; 
 QEA <=  JEA & jeb & jec  |  jea & JEB & jec  |  jea & jeb & JEC  |  JEA & JEB & JEC  ;
 DDN <= ddg & DDJ ; 
 TDB <= ddg & DDN ; 
 QEB <=  JED & jee & jef  |  jed & JEE & jef  |  jed & jee & JEF  |  JED & JEE & JEF  ;
 qca <=  aad  |  bap  ; 
 qcb <=  aae  |  bap  ; 
 WDC <=  HDC  |  HDK  ; 
 WDD <=  HDD  |  HDL  ; 
 QEC <=  JEG & jeh  |  jeg & JEH  ; 
 qcc <=  aaf  |  bap  ; 
 WDE <=  HDE  |  HDM  ; 
 WDF <=  HDF  |  HDN  ; 
 DDO <= ddg & DDK ; 
 TDC <= ddg & DDO ; 
 DDP <= ddg & DDL ; 
 TDD <= ddg & DDP ; 
 WDG <=  HDG  |  HDO  ; 
 WDH <=  HDH  |  HDP  ; 
 TJB <=  FEB  |  TIB  ; 
 TKB <=  FEB  |  TIB  ; 
 ORA <=  QEA & qeb & qec  |  qea & QEB & qec  |  qea & qeb & QEC  |  QEA & QEB & QEC  ;
 ddi <=  idh  |  IDB  |  IDA  ; 
 ddj <=  idh  |  IDB  |  ida  ; 
 ddk <=  idh  |  idb  |  IDA  ; 
 ddl <=  idh  |  idb  |  ida  ; 
 TJC <=  FEC  |  TIC  ; 
 TKC <=  FEC  |  TIC  ; 
 cae <=  ITF  |  ITE  |  itd  ; 
 SEC <=  GAK & TSE  |  GBK & TSE  |  SEC & tse  ; 
 SED <=  GAL & TSE  |  GBL & TSE  |  SED & tse  ; 
 GAD <=  IRD & CAE  |  IPD & CAF  |  IQD & CAG  |  MAD  ; 
 GAL <=  IRD & CAE  |  IPD & CAF  |  IQD & CAG  |  MAD  ; 
 TJD <=  FED  |  TID  ; 
 TKD <=  FED  |  TID  ; 
 caf <=  ITF  |  ite  |  ITD  ; 
 cag <=  ITF  |  ite  |  itd  ; 
 SFC <=  GAK & TSF  |  GBK & TSF  |  SFC & tsf  ; 
 SFD <=  GAL & TSF  |  GBL & TSF  |  SFD & tsf  ; 
 cah <=  itf  |  ITE  |  ITD  ; 
 cai <=  itf  |  ITE  |  itd  ; 
 NEB <= FAE ; 
 NGB <= FAG ; 
 SJD <= SKD ; 
 TIE <= FEE ; 
 TIF <= FEF ; 
 TIG <= FEG ; 
 CAD <=  ITF  |  ITE  |  ITD  ; 
 caj <=  itf  |  ite  |  ITD  ; 
 DDG <= IDG ; 
 NFB <= FAF ; 
 NHB <= FAH ; 
 TJE <=  FEE  |  TIE  ; 
 TKE <=  FEE  |  TIE  ; 
 SGC <=  GAK & TSG  |  GBK & TSG  |  SGC & tsg  ; 
 SGD <=  GAL & TSG  |  GBL & TSG  |  SGD & tsg  ; 
 oad <= jbd & jad ; 
 obd <= jbd & jad ; 
 ocd <= jbd & jad ; 
 skd <= jbd & jad ; 
 TJF <=  FEF  |  TIF  ; 
 TKF <=  FEF  |  TIF  ; 
 oqa <=  EAA  |  EAB  |  EAC  |  EAD  ; 
 SHC <=  GAK & TSH  |  GBK & TSH  |  SHC & tsg  ; 
 SHD <=  GAL & TSH  |  GBL & TSH  |  SHD & tsg  ; 
 GBD <=  IND & CAH  |  IOD & CAI  |  IMD & CAJ  |  IID  |  IJD  ; 
 GBL <=  IND & CAH  |  IOD & CAI  |  IMD & CAJ  |  IID  |  IJD  ; 
 TJG <=  FEG  |  TIG  ; 
 TKG <=  FEG  |  TIG  ; 
 LDA <= BAD & FDD |  LDA & fdd ; 
 LDB <= BAE & FDD |  LDB & fdd ; 
 LDC <= BAF & FDD |  LDC & fdd ; 
 DDC <= IDC ; 
 DDD <= IDD ; 
 DDE <= IDE ; 
 DDF <= IDF ; 
 UEA <= DEG & DEI |  ZZO & dei ; 
 UEB <= UEA & DEI |  UEA & dei ; 
 UEC <= DEC & DEI |  UEC & dei ; 
 VEA <=  REA & TEA  |  REI & TEB  |  RMA & TEC  |  RMI & TED  ; 
 VEI <=  REA & TEA  |  REI & TEB  |  RMA & TEC  |  RMI & TED  ; 
 UED <= DED & DEI |  UED & dei ; 
 UEE <= DEE & DEI |  UEE & dei ; 
 UEF <= DEF & DEI |  UEF & dei ; 
 VEB <=  REB & TEA  |  REJ & TEB  |  RMB & TEC  |  RMJ & TED  ; 
 VEJ <=  REB & TEA  |  REJ & TEB  |  RMB & TEC  |  RMJ & TED  ; 
 UEG <= DEG & DEJ |  ZZO & dej ; 
 UEH <= UEG & DEJ |  UEG & dej ; 
 UEI <= DEC & DEJ |  UEI & dej ; 
 VEC <=  REC & TEA  |  REK & TEB  |  RMC & TEC  |  RMK & TED  ; 
 VEK <=  REC & TEA  |  REK & TEB  |  RMC & TEC  |  RMK & TED  ; 
 VEG <=  REG & TEA  |  REO & TEB  |  RMG & TEC  |  RMO & TED  ; 
 VEO <=  REG & TEA  |  REO & TEB  |  RMG & TEC  |  RMO & TED  ; 
 UEJ <= DED & DEJ |  UEJ & dej ; 
 UEK <= DEE & DEJ |  UEK & dej ; 
 UEL <= DEF & DEJ |  UEL & dej ; 
 VED <=  RED & TEA  |  REL & TEB  |  RMD & TEC  |  RML & TED  ; 
 VEL <=  RED & TEA  |  REL & TEB  |  RMD & TEC  |  RML & TED  ; 
 UEM <= DEG & DEK |  ZZO & dek ; 
 UEN <= UEM & DEK |  UEM & dek ; 
 UEO <= DEC & DEK |  UEO & dek ; 
 VEE <=  REE & TEA  |  REM & TEB  |  RME & TEC  |  RMM & TED  ; 
 VEM <=  REE & TEA  |  REM & TEB  |  RME & TEC  |  RMM & TED  ; 
 UEP <= DED & DEK |  UEP & dek ; 
 UEQ <= DEE & DEK |  UEQ & dek ; 
 UER <= DEF & DEK |  UER & dek ; 
 VEF <=  REFF  & TEA  |  REN & TEB  |  RMF & TEC  |  RMN & TED  ; 
 VEN <=  REFF  & TEA  |  REN & TEB  |  RMF & TEC  |  RMN & TED  ; 
 UEU <= DEC & DEL |  UEU & del ; 
 UES <= DEG & DEL |  ZZO & del ; 
 UET <= UES & DEL |  UES & del ; 
 UEV <= DED & DEL |  UEV & del ; 
 UEW <= DEE & DEL |  UEW & del ; 
 UEX <= DEF & DEL |  UEX & del ; 
 VEH <=  REH & TEA  |  REP & TEB  |  RMH & TEC  |  RMP & TED  ; 
 VEP <=  REH & TEA  |  REP & TEB  |  RMH & TEC  |  RMP & TED  ; 
 WEA <=  HEA  |  HEI  ; 
 WEB <=  HEB  |  HEJ  ; 
 DEM <= deg & DEI ; 
 TEA <= deg & DEM ; 
 TEB <= deg & DEN ; 
 DEN <= deg & DEJ ; 
 BAJ <= FCB ; 
 BAK <= FCC ; 
 BAL <= FCD ; 
 BBA <= ABA ; 
 BBB <= ABB ; 
 BBC <= ABC ; 
 WEC <=  HEC  |  HEK  ; 
 WED <=  HED  |  HEL  ; 
 BAM <= FCE ; 
 BAN <= FCF ; 
 BAO <= FCG ; 
 BAP <= FCH ; 
 WEE <=  HEE  |  HEM  ; 
 WEF <=  HEF  |  HEN  ; 
 DEO <= deg & DEK ; 
 TEC <= deg & DEO ; 
 DEP <= deg & DEL ; 
 TED <= deg & DEP ; 
 WEG <=  HEG  |  HEO  ; 
 WEH <=  HEH  |  HEP  ; 
 TSA <= FBA ; 
 TSB <= FBB ; 
 TSC <= FBC ; 
 TSD <= FBD ; 
 dei <=  ieh  |  IEB  |  IEA  ; 
 dej <=  ieh  |  IEB  |  iea  ; 
 dek <=  ieh  |  ieb  |  IEA  ; 
 del <=  ieh  |  ieb  |  iea  ; 
 TSE <= FBE ; 
 TSF <= FBF ; 
 TSG <= FBG ; 
 TSH <= FBH ; 
 SAE <=  GAE & TSA  |  GBE & TSA  |  SAE & tsa  ; 
 SAF <=  GAF & TSA  |  GBF & TSA  |  SAF & tsa  ; 
 GAE <=  IRE & CAE  |  IPE & CAF  |  IQE & CAG  |  MAE  ; 
 GAM <=  IRE & CAE  |  IPE & CAF  |  IQE & CAG  |  MAE  ; 
 CAA <= ITA ; 
 CAB <= ITB ; 
 CAC <= ITC ; 
 SBE <=  GAE & TSB  |  GBE & TSB  |  SBE & tsb  ; 
 SBF <=  GAF & TSB  |  GBF & TSB  |  SBF & tsb  ; 
 aba <= isa ; 
 abb <= isb ; 
 abc <= isc ; 
 NAC <= FAA ; 
 NCC <= FAC ; 
 SJE <= SKE ; 
 QAA <=  ISF & qaa  |  ISE & qaa  |  ISD & qaa  ; 
 QAB <=  ISF & qaa  |  ISE & qaa  |  ISD & qaa  ; 
 QAC <=  ISF & qaa  |  ISE & qaa  |  ISD & qaa  ; 
 AAA <= ISA ; 
 AAB <= ISB ; 
 AAC <= ISC ; 
 DEG <= IEG ; 
 NBC <= FAB ; 
 NDC <= FAD ; 
 OQB <= EAE ; 
 QBA <=  QAC & AAG  ; 
 SCF <=  GAF & TSC  |  GBF & TSC  |  SCF & tsc  ; 
 SCE <=  GAE & TSC  |  GBE & TSC  |  SCE & tsc  ; 
 oae <= jbe & jae ; 
 obe <= jbe & jae ; 
 oce <= jbe & jae ; 
 ske <= jbe & jae ; 
 AAD <= ISD ; 
 AAE <= ISE ; 
 AAF <= ISF ; 
 AAG <= ISG ; 
 SDE <=  GAE & TSD  |  GBE & TSD  |  SDE & tsd  ; 
 SDF <=  GAF & TSD  |  GBF & TSD  |  SDF & tsd  ; 
 GBE <=  INE & CAH  |  IOE & CAI  |  IME & CAJ  |  IIE  |  IJE  ; 
 GBM <=  INE & CAH  |  IOE & CAI  |  IME & CAJ  |  IIE  |  IJE  ; 
 BAD <= AAD ; 
 BAE <= AAE ; 
 BAF <= AAF ; 
 LEA <= BAD & FDE |  LEA & fde ; 
 LEB <= BAE & FDE |  LEB & fde ; 
 LEC <= BAF & FDE |  LEC & fde ; 
 DEC <= IEC ; 
 DED <= IED ; 
 DEE <= IEE ; 
 DEF <= IEF ; 
 UFA <= DFG & DFI |  ZZO & dfi ; 
 UFB <= UFA & DFI |  UFA & dfi ; 
 UFC <= DFC & DFI |  UFC & dfi ; 
 VFA <=  RFA & TFA  |  RFI & TFB  |  RNA & TFC  |  RNI & TFD  ; 
 VFI <=  RFA & TFA  |  RFI & TFB  |  RNA & TFC  |  RNI & TFD  ; 
 UFD <= DFD & DFI |  UFD & dfi ; 
 UFE <= DFE & DFI |  UFE & dfi ; 
 UFF <= DFF & DFI |  UFF & dfi ; 
 VFB <=  RFB & TFA  |  RFJ & TFB  |  RNB & TFC  |  RNJ & TFD  ; 
 VFJ <=  RFB & TFA  |  RFJ & TFB  |  RNB & TFC  |  RNJ & TFD  ; 
 UFG <= DFG & DFJ |  ZZO & dfj ; 
 UFH <= UFG & DFJ |  UFG & dfj ; 
 UFI <= DFC & DFJ |  UFI & dfj ; 
 VFC <=  RFC & TFA  |  RFK & TFB  |  RNC & TFC  |  RNK & TFD  ; 
 VFK <=  RFC & TFA  |  RFK & TFB  |  RNC & TFC  |  RNK & TFD  ; 
 UFJ <= DFD & DFJ |  UFJ & dfj ; 
 UFK <= DFE & DFJ |  UFK & dfj ; 
 UFL <= DFF & DFJ |  UFL & dfj ; 
 VFD <=  RFD & TFA  |  RFL & TFB  |  RND & TFC  |  RNL & TFD  ; 
 VFL <=  RFD & TFA  |  RFL & TFB  |  RND & TFC  |  RNL & TFD  ; 
 UFM <= DFG & DFK |  ZZO & dfk ; 
 UFN <= UFM & DFK |  UFM & dfk ; 
 UFO <= DFC & DFK |  UFO & dfk ; 
 VFE <=  RFE & TFA  |  RFM & TFB  |  RNE & TFC  |  RNM & TFD  ; 
 VFM <=  RFE & TFA  |  RFM & TFB  |  RNE & TFC  |  RNM & TFD  ; 
 UFP <= DFD & DFK |  UFP & dfk ; 
 UFQ <= DFE & DFK |  UFQ & dfk ; 
 UFR <= DFF & DFK |  UFR & dfk ; 
 VFF <=  RFF & TFA  |  RFN & TFB  |  RNF & TFC  |  RNN & TFD  ; 
 VFN <=  RFF & TFA  |  RFN & TFB  |  RNF & TFC  |  RNN & TFD  ; 
 UFT <= UFS & DFL |  UFS & dfl ; 
 UFU <= DFC & DFL |  UFU & dfl ; 
 UFS <= DFG & DFL |  ZZO & dfl ; 
 VFG <=  RFG & TFA  |  RFO & TFB  |  RNG & TFC  |  RNO & TFD  ; 
 VFO <=  RFG & TFA  |  RFO & TFB  |  RNG & TFC  |  RNO & TFD  ; 
 UFV <= DFD & DFL |  UFV & dfl ; 
 UFW <= DFE & DFL |  UFW & dfl ; 
 UFX <= DFF & DFL |  UFX & dfl ; 
 VFH <=  RFH & TFA  |  RFP & TFB  |  RNH & TFC  |  RNP & TFD  ; 
 VFP <=  RFH & TFA  |  RFP & TFB  |  RNH & TFC  |  RNP & TFD  ; 
 WFA <=  HFA  |  HFI  ; 
 WFB <=  HFB  |  HFJ  ; 
 DFM <= dfg & DFI ; 
 DFN <= dfg & DFJ ; 
 TFA <= dfg & DFM ; 
 TFB <= dfg & DFN ; 
 kda <= ina ; 
 kdb <= inb ; 
 kdc <= inc ; 
 kdd <= ind ; 
 LLA <= BBA & BAM |  LLA & bam ; 
 LLB <= BBB & BAM |  LLB & bam ; 
 LLC <= BBC & BAM |  LLC & bam ; 
 WFC <=  HFC  |  HFK  ; 
 WFD <=  HFD  |  HFL  ; 
 LRA <= ABA & BAM |  LRA & bam ; 
 LRB <= ABB & BAM |  LRB & bam ; 
 LRC <= ABC & BAM |  LRC & bam ; 
 WFE <=  HFE  |  HFM  ; 
 WFF <=  HFF  |  HFN  ; 
 DFO <= dfg & DFK ; 
 DFP <= dfg & DFL ; 
 TFC <= dfg & DFO ; 
 TFD <= dfg & DFP ; 
 kde <= ine ; 
 kdf <= inf ; 
 kdg <= ing ; 
 kdh <= inh ; 
 WFG <=  HFG  |  HFO  ; 
 WFH <=  HFH  |  HFP  ; 
 OIA <=  HLA & HLI  ; 
 OJA <=  HRA & HRI & tje  |  JAI & TJE  |  JBI & TKE  ; 
 dfi <=  ifh  |  IFB  |  IFA  ; 
 dfj <=  ifh  |  IFB  |  ifa  ; 
 dfk <=  ifh  |  ifb  |  IFA  ; 
 dfl <=  ifh  |  ifb  |  ifa  ; 
 OIB <=  HLB & HLJ  ; 
 OJB <=  HRB & HRJ & tje  |  JAJ & TJE  |  JBJ & TKE  ; 
 SEE <=  GAM & TSE  |  GBM & TSE  |  SEE & tse  ; 
 SEF <=  GAN & TSE  |  GBN & TSE  |  SEF & tse  ; 
 GAF <=  IRF & CAE  |  IPF & CAF  |  IQF & CAG  |  MAF  ; 
 GAN <=  IRF & CAE  |  IPF & CAF  |  IQF & CAG  |  MAF  ; 
 OIC <=  HLC & HLK  ; 
 OJC <=  HRC & HRK & tje  |  JAK & TJE  |  JBK & TKE  ; 
 SFE <=  GAM & TSF  |  GBM & TSF  |  SFE & tsf  ; 
 SFF <=  GAN & TSF  |  GBN & TSF  |  SFF & tsf  ; 
 OID <=  HLD & HLL  ; 
 OJD <=  HRD & HRL & tje  |  JAL & TJE  |  JBL & TKE  ; 
 NEC <= FAE ; 
 NGC <= FAG ; 
 SJF <= SKF ; 
 OIE <=  HLE & HLM  ; 
 OJE <=  HRE & HRM & tje  |  JAM & TJE  |  JBM & TKE  ; 
 DFG <= IFG ; 
 NFC <= FAF ; 
 NHC <= FAH ; 
 OIF <=  HLF & HLN  ; 
 OJF <=  HRF & HRN & tje  |  JAN & TJE  |  JBN & TKE  ; 
 SGE <=  GAM & TSG  |  GBM & TSG  |  SGE & tsg  ; 
 SGF <=  GAN & TSG  |  GBN & TSG  |  SGF & tsg  ; 
 oaf <= jbf & jaf ; 
 obf <= jbf & jaf ; 
 ocf <= jbf & jaf ; 
 skf <= jbf & jaf ; 
 OIG <=  HLG & HLO  ; 
 OJG <=  HRG & HRO & tje  |  JAO & TJE  |  JBO & TKE  ; 
 SHE <=  GAM & TSH  |  GBM & TSH  |  SHE & tsg  ; 
 SHF <=  GAN & TSH  |  GBN & TSH  |  SHF & tsg  ; 
 GBF <=  INF & CAH  |  IOF & CAI  |  IMF & CAJ  |  IIF  |  IJF  ; 
 GBN <=  INF & CAH  |  IOF & CAI  |  IMF & CAJ  |  IIF  |  IJF  ; 
 OIH <=  HLH & HLP  ; 
 OJH <=  HRH & HRP & tje  |  JAP & TJE  |  JBP & TKE  ; 
 LFA <= BAD & FDF |  LFA & fdf ; 
 LFB <= BAE & FDF |  LFB & fdf ; 
 LFC <= BAF & FDF |  LFC & fdf ; 
 DFC <= IFC ; 
 DFD <= IFD ; 
 DFE <= IFE ; 
 DFF <= IFFF  ; 
 UGA <= DGG & DGI |  ZZO & dgi ; 
 UGB <= UGA & DGI |  UGA & dgi ; 
 UGC <= DGC & DGI |  UGC & dgi ; 
 VGA <=  RGA & TGA  |  RGI & TGB  |  ROA & TGC  |  ROI & TGD  ; 
 VGI <=  RGA & TGA  |  RGI & TGB  |  ROA & TGC  |  ROI & TGD  ; 
 UGD <= DGD & DGI |  UGD & dgi ; 
 UGE <= DGE & DGI |  UGE & dgi ; 
 UGF <= DGF & DGI |  UGF & dgi ; 
 VGB <=  RGB & TGA  |  RGJ & TGB  |  ROB & TGC  |  ROJ & TGD  ; 
 VGJ <=  RGB & TGA  |  RGJ & TGB  |  ROB & TGC  |  ROJ & TGD  ; 
 UGG <= DGG & DGJ |  ZZO & dgj ; 
 UGH <= UGG & DGJ |  UGG & dgj ; 
 UGI <= DGC & DGJ |  UGI & dgj ; 
 VGG <=  RGG & TGA  |  RGO & TGB  |  ROG & TGC  |  ROO & TGD  ; 
 VGO <=  RGG & TGA  |  RGO & TGB  |  ROG & TGC  |  ROO & TGD  ; 
 VGC <=  RGC & TGA  |  RGK & TGB  |  ROC & TGC  |  ROK & TGD  ; 
 VGK <=  RGC & TGA  |  RGK & TGB  |  ROC & TGC  |  ROK & TGD  ; 
 UGJ <= DGD & DGJ |  UGJ & dgj ; 
 UGK <= DGE & DGJ |  UGK & dgj ; 
 UGL <= DGF & DGJ |  UGL & dgj ; 
 VGD <=  RGD & TGA  |  RGL & TGB  |  ROD & TGC  |  ROL & TGD  ; 
 VGL <=  RGD & TGA  |  RGL & TGB  |  ROD & TGC  |  ROL & TGD  ; 
 UGM <= DGG & DGK |  ZZO & dgk ; 
 UGN <= UGM & DGK |  UGM & dgk ; 
 UGO <= DGC & DGK |  UGO & dgk ; 
 VGE <=  RGE & TGA  |  RGM & TGB  |  ROE & TGC  |  ROM & TGD  ; 
 VGM <=  RGE & TGA  |  RGM & TGB  |  ROE & TGC  |  ROM & TGD  ; 
 UGP <= DGD & DGK |  UGP & dgk ; 
 UGQ <= DGE & DGK |  UGQ & dgk ; 
 UGR <= DGF & DGK |  UGR & dgk ; 
 VGF <=  RGF & TGA  |  RGN & TGB  |  ROF & TGC  |  RON & TGD  ; 
 VGN <=  RGF & TGA  |  RGN & TGB  |  ROF & TGC  |  RON & TGD  ; 
 UGS <= DGG & DGL |  ZZO & dgl ; 
 UGT <= UGS & DGL |  UGS & dgl ; 
 UGU <= DGC & DGL |  UGU & dgl ; 
 UGV <= DGD & DGL |  UGV & dgl ; 
 UGW <= DGE & DGL |  UGW & dgl ; 
 UGX <= DGF & DGL |  UGX & dgl ; 
 VGH <=  RGH & TGA  |  RGP & TGB  |  ROH & TGC  |  ROP & TGD  ; 
 VGP <=  RGH & TGA  |  RGP & TGB  |  ROH & TGC  |  ROP & TGD  ; 
 WGA <=  HGA  |  HGI  ; 
 WGB <=  HGB  |  HGJ  ; 
 DGM <= dgg & DGI ; 
 DGN <= dgg & DGJ ; 
 TGA <= dgg & DGM ; 
 TGB <= dgg & DGN ; 
 kea <= ioa ; 
 keb <= iob ; 
 kec <= ioc ; 
 ked <= iod ; 
 LMA <= BBA & BAN |  LMA & ban ; 
 LMB <= BBB & BAN |  LMB & ban ; 
 LMC <= BBC & BAN |  LMC & ban ; 
 WGC <=  HGC  |  HGK  ; 
 WGD <=  HGD  |  HGL  ; 
 TIB <= FEB ; 
 TIC <= FEC ; 
 TID <= FED ; 
 LSA <= ABA & BAN |  LSA & ban ; 
 LSB <= ABB & BAN |  LSB & ban ; 
 LSC <= ABC & BAN |  LSC & ban ; 
 WGE <=  HGE  |  HGM  ; 
 WGF <=  HGF  |  HGN  ; 
 DGO <= dgg & DGK ; 
 DGP <= dgg & DGL ; 
 TGC <= dgg & DGO ; 
 TGD <= dgg & DGP ; 
 kee <= ioe ; 
 kef <= iof ; 
 keg <= iog ; 
 keh <= ioh ; 
 WGG <=  HGG  |  HGO  ; 
 WGH <=  HGH  |  HGP  ; 
 OKA <=  HMA & HMI  ; 
 OLA <=  HSA & HSI & tjf  |  JAI & TJF  |  JBI & TKF  ; 
 dgi <=  igh  |  IGB  |  IGA  ; 
 dgj <=  igh  |  IGB  |  iga  ; 
 dgk <=  igh  |  igb  |  IGA  ; 
 dgl <=  igh  |  igb  |  iga  ; 
 OKB <=  HMB & HMJ  ; 
 OLB <=  HSB & HSJ & tjf  |  JAJ & TJF  |  JBJ & TKF  ; 
 SAG <=  GAG & TSA  |  GBG & TSA  |  SAG & tsa  ; 
 SAH <=  GAH & TSA  |  GBH & TSA  |  SAH & tsa  ; 
 GAG <=  IRG & CAE  |  IPG & CAF  |  IQG & CAG  |  MAG  ; 
 GAO <=  IRG & CAE  |  IPG & CAF  |  IQG & CAG  |  MAG  ; 
 OKC <=  HMC & HMK  ; 
 OLC <=  HSC & HSK & tjf  |  JAK & TJF  |  JBK & TKF  ; 
 SBG <=  GAG & TSB  |  GBG & TSB  |  SBG & tsb  ; 
 SBH <=  GAH & TSB  |  GBH & TSB  |  SBH & tsb  ; 
 OKD <=  HMD & HML  ; 
 OLD <=  HSD & HSL & tjf  |  JAL & TJF  |  JBL & TKF  ; 
 NAD <= FAA ; 
 NCD <= FAC ; 
 SJG <= SKG ; 
 OKE <=  HME & HMM  ; 
 OLE <=  HSE & HSM & tjf  |  JAM & TJF  |  JBM & TKF  ; 
 DGG <= IGG ; 
 NBD <= FAB ; 
 NDD <= FAD ; 
 OKF <=  HMF & HMM  ; 
 OLF <=  HSF & HSN & tjf  |  JAN & TJF  |  JBN & TKF  ; 
 SCG <=  GAG & TSC  |  GBG & TSC  |  SCG & tsc  ; 
 SCH <=  GAH & TSC  |  GBH & TSC  |  SCH & tsc  ; 
 oag <= jbg & jag ; 
 obg <= jbg & jag ; 
 ocg <= jbg & jag ; 
 skg <= jbg & jag ; 
 OKG <=  HMG & HMO  ; 
 OLG <=  HSG & HSO & tjf  |  JAO & TJF  |  JBO & TKF  ; 
 SDG <=  GAG & TSD  |  GBG & TSD  |  SDG & tsd  ; 
 SDH <=  GAH & TSD  |  GBH & TSD  |  SDH & tsd  ; 
 GBG <=  ING & CAH  |  IOG & CAI  |  IMG & CAJ  |  IIG  |  IJG  ; 
 GBO <=  ING & CAH  |  IOG & CAI  |  IMG & CAJ  |  IIG  |  IJG  ; 
 OKH <=  HMH & HMP  ; 
 OLH <=  HSH & HSP & tjf  |  JAP & TJF  |  JBP & TKF  ; 
 LGA <= BAD & FDG |  LGA & fdg ; 
 LGB <= BAE & FDG |  LGB & fdg ; 
 LGC <= BAF & FDG |  LGC & fdg ; 
 DGC <= IGC ; 
 DGD <= IGD ; 
 DGE <= IGE ; 
 DGF <= IGF ; 
 UHA <= DHG & DHI |  ZZO & dhi ; 
 UHB <= UHA & DHI |  UHA & dhi ; 
 UHC <= DHC & DHI |  UHC & dhi ; 
 VHA <=  RHA & THA  |  RHI & THB  |  RPA & THC  |  RPI & THD  ; 
 VHI <=  RHA & THA  |  RHI & THB  |  RPA & THC  |  RPI & THD  ; 
 UHD <= DHD & DHI |  UHD & dhi ; 
 UHE <= DHE & DHI |  UHE & dhi ; 
 UHF <= DHF & DHI |  UHF & dhi ; 
 VHB <=  RHB & THA  |  RHJ & THB  |  RPB & THC  |  RPJ & THD  ; 
 VHJ <=  RHB & THA  |  RHJ & THB  |  RPB & THC  |  RPJ & THD  ; 
 UHG <= DHG & DHJ |  ZZO & dhj ; 
 UHH <= UHG & DHJ |  UHG & dhj ; 
 UHI <= DHC & DHJ |  UHI & dhj ; 
 VHC <=  RHC & THA  |  RHK & THB  |  RPC & THC  |  RPK & THD  ; 
 VHK <=  RHC & THA  |  RHK & THB  |  RPC & THC  |  RPK & THD  ; 
 UHJ <= DHD & DHJ |  UHJ & dhj ; 
 UHK <= DHE & DHJ |  UHK & dhj ; 
 UHL <= DHF & DHJ |  UHL & dhj ; 
 VHD <=  RHD & THA  |  RHL & THB  |  RPD & THC  |  RPL & THD  ; 
 VHL <=  RHD & THA  |  RHL & THB  |  RPD & THC  |  RPL & THD  ; 
 UHM <= DHG & DHK |  ZZO & dhk ; 
 UHN <= UHM & DHK |  UHM & dhk ; 
 VHE <=  RHE & THA  |  RHM & THB  |  RPE & THC  |  RPM & THD  ; 
 VHM <=  RHE & THA  |  RHM & THB  |  RPE & THC  |  RPM & THD  ; 
 UHO <= DHC & DHK |  UHO & dhk ; 
 UHP <= DHD & DHK |  UHP & dhk ; 
 VHN <=  RHF & THA  |  RHN & THB  |  RPF & THC  |  RPN & THD  ; 
 VHF <=  RHF & THA  |  RHN & THB  |  RPF & THC  |  RPN & THD  ; 
 UHS <= DHG & DHL |  ZZO & dhl ; 
 UHT <= UHS & DHL |  UHS & dhl ; 
 UHU <= DHC & DHL |  UHU & dhl ; 
 VHG <=  RHG & THA  |  RHO & THB  |  RPG & THC  |  RPO & THD  ; 
 VHO <=  RHG & THA  |  RHO & THB  |  RPG & THC  |  RPO & THD  ; 
 UHV <= DHD & DHL |  UHV & dhl ; 
 UHW <= DHE & DHL |  UHW & dhl ; 
 UHX <= DHF & DHL |  UHX & dhl ; 
 VHH <=  RHH & THA  |  RHP & THB  |  RPH & THC  |  RPP & THD  ; 
 VHP <=  RHH & THA  |  RHP & THB  |  RPH & THC  |  RPP & THD  ; 
 WHA <=  HHA  |  HHI  ; 
 WHB <=  HHB  |  HHJ  ; 
 DHM <= dhg & DHI ; 
 DHN <= dhg & DHJ ; 
 THA <= dhg & DHM ; 
 THB <= dhg & DHN ; 
 kfa <= ima ; 
 kfb <= imb ; 
 kfc <= imc ; 
 kfd <= imd ; 
 LNA <= BBA & BAO |  LNA & bao ; 
 LNB <= BBB & BAO |  LNB & bao ; 
 LNC <= BBC & BAO |  LNC & bao ; 
 WHC <=  HHC  |  HHK  ; 
 WHD <=  HHD  |  HHL  ; 
 kfe <= ime ; 
 kff <= imf ; 
 kfg <= img ; 
 kfh <= imh ; 
 LTA <= ABA & BAO |  LTA & bao ; 
 LTB <= ABB & BAO |  LTB & bao ; 
 LTC <= ABC & BAO |  LTC & bao ; 
 WHE <=  HHE  |  HHM  ; 
 WHF <=  HHF  |  HHN  ; 
 DHO <= dhg & DHK ; 
 DHP <= dhg & DHL ; 
 THD <= dhg & DHP ; 
 THC <= dhg & DHO ; 
 UHQ <= DHE & DHK |  UHQ & dhk ; 
 UHR <= DHF & DHK |  UHR & dhk ; 
 WHG <=  HHG  |  HHO  ; 
 WHH <=  HHH  |  HHP  ; 
 OGA <=  HNA & HNI  ; 
 OHA <=  HTA & HTI & tjg  |  JAI & TJG  |  JBI & TKG  ; 
 dhi <=  ihh  |  IHB  |  IHA  ; 
 dhj <=  ihh  |  IHB  |  iha  ; 
 dhk <=  ihh  |  ihb  |  IHA  ; 
 dhl <=  ihh  |  ihb  |  iha  ; 
 OGB <=  HNB & HNJ  ; 
 OHB <=  HTB & HTJ & tjg  |  JAJ & TJG  |  JBJ & TKG  ; 
 SEG <=  GAO & TSE  |  GBO & TSE  |  SEG & tse  ; 
 SEH <=  GAP & TSE  |  GBP & TSE  |  SEH & tse  ; 
 GAH <=  IRH & CAE  |  IPH & CAF  |  IQH & CAG  |  MAH  ; 
 GAP <=  IRH & CAE  |  IPH & CAF  |  IQH & CAG  |  MAH  ; 
 OGC <=  HNC & HNK  ; 
 OHC <=  HTC & HTK & tjg  |  JAK & TJG  |  JBK & TKG  ; 
 SFG <=  GAO & TSF  |  GBO & TSF  |  SFG & tsf  ; 
 SFH <=  GAP & TSF  |  GBP & TSF  |  SFH & tsf  ; 
 OGD <=  HND & HNL  ; 
 OHD <=  HTD & HTL & tjg  |  JAL & TJG  |  JBL & TKG  ; 
 NED <= FAE ; 
 NGD <= FAG ; 
 SJH <= SKH ; 
 OGE <=  HNE & HNM  ; 
 OHE <=  HTE & HTM & tjg  |  JAM & TJG  |  JBM & TKG  ; 
 DHG <= IHG ; 
 NFD <= FAF ; 
 NHD <= FAH ; 
 OGF <=  HNF & HNN  ; 
 OHF <=  HTF & HTN & tjg  |  JAN & TJG  |  JBN & TKG  ; 
 SGG <=  GAO & TSG  |  GBO & TSG  |  SGG & tsg  ; 
 SGH <=  GAP & TSG  |  GBP & TSG  |  SGH & tsg  ; 
 oah <= jbh & jah ; 
 obh <= jbh & jah ; 
 och <= jbh & jah ; 
 skh <= jbh & jah ; 
 OGG <=  HNG & HNO  ; 
 OHG <=  HTG & HTO & tjg  |  JAO & TJG  |  JBO & TKG  ; 
 SHG <=  GAO & TSH  |  GBO & TSH  |  SHG & tsg  ; 
 SHH <=  GAP & TSH  |  GBP & TSH  |  SHH & tsg  ; 
 GBH <=  INH & CAH  |  IOH & CAI  |  IMH & CAJ  |  IIH  |  IJH  ; 
 GBP <=  INH & CAH  |  IOH & CAI  |  IMH & CAJ  |  IIH  |  IJH  ; 
 OGH <=  HNH & HNP  ; 
 OHH <=  HTH & HTP & tjg  |  JAP & TJG  |  JBP & TKG  ; 
 LHA <= BAD & FDH |  LHA & fdh ; 
 LHB <= BAE & FDH |  LHB & fdh ; 
 LHC <= BAF & FDH |  LHC & fdh ; 
 DHC <= IHC ; 
 DHD <= IHD ; 
 DHE <= IHE ; 
 DHF <= IHF ; 
end 
ram_16x4 rinst_0( RAA,RAB,RAC,RAD, WAA,WAB,WAC,WAD, UAC,UAD,UAE,UAF, ZZI, UAB, IZZ); 
ram_16x4 rinst_1( RAE,RAF,RAG,RAH, WAE,WAF,WAG,WAH, UAC,UAD,UAE,UAF, ZZI, UAB, IZZ); 
ram_16x4 rinst_2( RAI,RAJ,RAK,RAL, WAA,WAB,WAC,WAD, UAI,UAJ,UAK,UAL, ZZI, UAH, IZZ); 
ram_16x4 rinst_3( RAM,RAN,RAO,RAP, WAE,WAF,WAG,WAH, UAI,UAJ,UAK,UAL, ZZI, UAH, IZZ); 
ram_16x4 rinst_4( RIA,RIB,RIC,RID, WAA,WAB,WAC,WAD, UAO,UAP,UAQ,UAR, ZZI, UAN, IZZ); 
ram_16x4 rinst_5( RIE,RIF,RIG,RIH, WAE,WAF,WAG,WAH, UAO,UAP,UAQ,UAR, ZZI, UAN, IZZ); 
ram_16x4 rinst_6( RII,RIJ,RIK,RIL, WAA,WAB,WAC,WAD, UAU,UAV,UAW,UAX, ZZI, UAT, IZZ); 
ram_16x4 rinst_7( RIM,RIN,RIO,RIP, WAE,WAF,WAG,WAH, UAU,UAV,UAW,UAX, ZZI, UAT, IZZ); 
ram_16x4 rinst_8( RBA,RBB,RBC,RBD, WBA,WBB,WBC,WBD, UBC,UBD,UBE,UBF, ZZI, UBB, IZZ); 
ram_16x4 rinst_9( RBE,RBF,RBG,RBH, WBE,WBF,WBG,WBH, UBC,UBD,UBE,UBF, ZZI, UBB, IZZ); 
ram_16x4 rinst_10( RBI,RBJ,RBK,RBL, WBA,WBB,WBC,WBD, UBI,UBJ,UBK,UBL, ZZI, UBH, IZZ); 
ram_16x4 rinst_11( RBM,RBN,RBO,RBP, WBE,WBF,WBG,WBH, UBI,UBJ,UBK,UBL, ZZI, UBH, IZZ); 
ram_16x4 rinst_12( RJA,RJB,RJC,RJD, WBA,WBB,WBC,WBD, UBO,UBP,UBQ,UBR, ZZI, UBN, IZZ); 
ram_16x4 rinst_13( RJE,RJF,RJG,RJH, WBE,WBF,WBG,WBH, UBO,UBP,UBQ,UBR, ZZI, UBN, IZZ); 
ram_16x4 rinst_14( RJI,RJJ,RJK,RJL, WBA,WBB,WBC,WBD, UBU,UBV,UBW,UBX, ZZI, UBT, IZZ); 
ram_16x4 rinst_15( RJM,RJN,RJO,RJP, WBE,WBF,WBG,WBH, UBU,UBV,UBW,UBX, ZZI, UBT, IZZ); 
ram_16x4 rinst_16( RCA,RCB,RCC,RCD, WCA,WCB,WCC,WCD, UCC,UCD,UCE,UCF, ZZI, UCB, IZZ); 
ram_16x4 rinst_17( RCE,RCF,RCG,RCH, WCE,WCF,WCG,WCH, UCC,UCD,UCE,UCF, ZZI, UCB, IZZ); 
ram_16x4 rinst_18( RCI,RCJ,RCK,RCL, WCA,WCB,WCC,WCD, UCI,UCJ,UCK,UCL, ZZI, UCH, IZZ); 
ram_16x4 rinst_19( RCM,RCN,RCO,RCP, WCE,WCF,WCG,WCH, UCI,UCJ,UCK,UCL, ZZI, UCH, IZZ); 
ram_16x4 rinst_20( RKA,RKB,RKC,RKD, WCA,WCB,WCC,WCD, UCO,UCP,UCQ,UCR, ZZI, UCN, IZZ); 
ram_16x4 rinst_21( RKE,RKF,RKG,RKH, WCE,WCF,WCG,WCH, UCO,UCP,UCQ,UCR, ZZI, UCN, IZZ); 
ram_16x4 rinst_22( RKI,RKJ,RKK,RKL, WCA,WCB,WCC,WCD, UCU,UCV,UCW,UCX, ZZI, UCT, IZZ); 
ram_16x4 rinst_23( RKM,RKN,RKO,RKP, WCE,WCF,WCG,WGH, UCU,UCV,UCW,UCX, ZZI, UCT, IZZ); 
ram_16x4 rinst_24( RDA,RDB,RDC,RDD, WDA,WDB,WDC,WDD, UDC,UDD,UDE,UDF, ZZI, UDB, IZZ); 
ram_16x4 rinst_25( RDE,RDF,RDG,RDH, WDE,WDF,WDG,WDH, UDC,UDD,UDE,UDF, ZZI, UDB, IZZ); 
ram_16x4 rinst_26( RDI,RDJ,RDK,RDL, WDA,WDB,WDC,WDD, UDI,UDJ,UDK,UDL, ZZI, UDH, IZZ); 
ram_16x4 rinst_27( RDM,RDN,RDO,RDP, WDE,WDF,WDG,WDH, UDI,UDJ,UDK,UDL, ZZI, UDH, IZZ); 
ram_16x4 rinst_28( RLA,RLB,RLC,RLD, WDA,WDB,WDC,WDD, UDO,UDP,UDQ,UDR, ZZI, UDN, IZZ); 
ram_16x4 rinst_29( RLE,RLF,RLG,RLH, WDE,WDF,WDG,WDH, UDO,UDP,UDQ,UDR, ZZI, UDN, IZZ); 
ram_16x4 rinst_30( RLI,RLJ,RLK,RLL, WDA,WDB,WDC,WDD, UDU,UDV,UDW,UDX, ZZI, UDT, IZZ); 
ram_16x4 rinst_31( RLM,RLN,RLO,RLP, WDE,WDF,WDG,WDH, UDU,UDV,UDW,UDX, ZZI, UDT, IZZ); 
ram_16x4 rinst_32( REA,REB,REC,RED, WEA,WEB,WEC,WED, UEC,UED,UEE,UEF, ZZI, UEB, IZZ); 
ram_16x4 rinst_33( REE,REFF ,REG,REH, WEE,WEF,WEG,WEH, UEC,UED,UEE,UEF, ZZI, UEB, IZZ); 
ram_16x4 rinst_34( REI,REJ,REK,REL, WEA,WEB,WEC,WED, UEI,UEJ,UEK,UEL, ZZI, UEH, IZZ); 
ram_16x4 rinst_35( REM,REN,REO,REP, WEE,WEF,WEG,WEH, UEI,UEJ,UEK,UEL, ZZI, UEH, IZZ); 
ram_16x4 rinst_36( RMA,RMB,RMC,RMD, WEA,WEB,WEC,WED, UEO,UEP,UEQ,UER, ZZI, UEN, IZZ); 
ram_16x4 rinst_37( RME,RMF,RMG,RMH, WEE,WEF,WEG,WEH, UEO,UEP,UEQ,UER, ZZI, UEN, IZZ); 
ram_16x4 rinst_38( RMI,RMJ,RMK,RML, WEA,WEB,WEC,WED, UEU,UEV,UEW,UEX, ZZI, UET, IZZ); 
ram_16x4 rinst_39( RMM,RMN,RMO,RMP, WEE,WEF,WEG,WEH, UEU,UEV,UEW,UEX, ZZI, UET, IZZ); 
ram_16x4 rinst_40( RFA,RFB,RFC,RFD, WFA,WFB,WFC,WFD, UFC,UFD,UFE,UFF, ZZI, UFB, IZZ); 
ram_16x4 rinst_41( RFE,RFF,RFG,RFH, WFE,WFF,WFG,WFH, UFC,UFD,UFE,UFF, ZZI, UFB, IZZ); 
ram_16x4 rinst_42( RFI,RFJ,RFK,RFL, WFA,WFB,WFC,WFD, UFI,UFJ,UFK,UFL, ZZI, UFH, IZZ); 
ram_16x4 rinst_43( RFM,RFN,RFO,RFP, WFE,WFF,WFG,WFH, UFI,UFJ,UFK,UFL, ZZI, UFH, IZZ); 
ram_16x4 rinst_44( RNA,RNB,RNC,RND, WFA,WFB,WFC,WFD, UFO,UFP,UFQ,UFR, ZZI, UFN, IZZ); 
ram_16x4 rinst_45( RNE,RNF,RNG,RNH, WFE,WFF,WFG,WFH, UFO,UFP,UFQ,UFR, ZZI, UFN, IZZ); 
ram_16x4 rinst_46( RNI,RNJ,RNK,RNL, WFA,WFB,WFC,WFD, UFU,UFV,UFW,UFX, ZZI, UFT, IZZ); 
ram_16x4 rinst_47( RNM,RNN,RNO,RNP, WFE,WFF,WFG,WFH, UFU,UFV,UFW,UFX, ZZI, UFT, IZZ); 
ram_16x4 rinst_48( RGA,RGB,RGC,RGD, WGA,WGB,WGC,WGD, UGC,UGD,UGE,UGF, ZZI, UGB, IZZ); 
ram_16x4 rinst_49( RGE,RGF,RGG,RGH, WGE,WGF,WGG,WGH, UGC,UGD,UGE,UGF, ZZI, UGB, IZZ); 
ram_16x4 rinst_50( RGM,RGN,RGO,RGP, WGE,WGF,WGG,WGH, UGI,UGJ,UGK,UGL, ZZI, UGH, IZZ); 
ram_16x4 rinst_51( ROA,ROB,ROC,ROD, WGA,WGB,WGC,WGD, UGO,UGP,UGQ,UGR, ZZI, UGN, IZZ); 
ram_16x4 rinst_52( ROE,ROF,ROG,ROH, WGE,WGF,WGG,WGH, UGO,UGP,UGQ,UGR, ZZI, UGN, IZZ); 
ram_16x4 rinst_53( ROI,ROJ,ROK,ROL, WGA,WGB,WGC,WGD, UGU,UGV,UGW,UGX, ZZI, UGT, IZZ); 
ram_16x4 rinst_54( RGI,RGJ,RGK,RGL, WGA,WGB,WGC,WGD, UGI,UGJ,UGK,UGL, ZZI, UGH, IZZ); 
ram_16x4 rinst_55( ROM,RON,ROO,ROP, WGE,WGF,WGG,WGH, UGU,UGV,UGW,UGX, ZZI, UGT, IZZ); 
ram_16x4 rinst_56( RHA,RHB,RHC,RHD, WHA,WHB,WHC,WHD, UHC,UHD,UHE,UHF, ZZI, UHB, IZZ); 
ram_16x4 rinst_57( RHE,RHF,RHG,RHH, WHE,WHF,WHG,WHH, UHC,UHD,UHE,UHF, ZZI, UHB, IZZ); 
ram_16x4 rinst_58( RHI,RHJ,RHK,RHL, WHA,WHB,WHC,WHD, UHI,UHJ,UHK,UHL, ZZI, UHH, IZZ); 
ram_16x4 rinst_59( RHM,RHN,RHO,RHP, WHE,WHF,WHG,WHH, UHI,UHJ,UHK,UHL, ZZI, UHH, IZZ); 
ram_16x4 rinst_60( RPA,RPB,RPC,RPD, WHA,WHB,WHC,WHD, UHO,UHP,UHQ,UHR, ZZI, UHN, IZZ); 
ram_16x4 rinst_61( RPE,RPF,RPG,RPH, WHE,WHF,WHG,WHH, UHO,UHP,UHQ,UHR, ZZI, UHN, IZZ); 
ram_16x4 rinst_62( RPI,RPJ,RPK,RPL, WHA,WHB,WHC,WHD, UHU,UHV,UHW,UHX, ZZI, UHT, IZZ); 
ram_16x4 rinst_63( RPM,RPN,RPO,RPP, WHE,WHF,WHG,WHH, UHU,UHV,UHH,UHX, ZZI, UHT, IZZ); 
endmodule;
