module as( IZZ,
 IAA, 
 IAB, 
 IAC, 
 IAD, 
 IAE, 
 IAF, 
 IAG, 
 IAH, 
 ICA, 
 ICB, 
 ICC, 
 ICD, 
 ICE, 
 ICF, 
 ICG, 
 ICH, 
 IEA, 
 IEB, 
 IEC, 
 IED, 
 IEE, 
 IEF, 
 IEG, 
 IEH, 
 IGA, 
 IGB, 
 IGC, 
 IGD, 
 IGE, 
 IGF, 
 IGG, 
 IGH, 
 IIA, 
 IJA, 
 IKA, 
 ILA, 
 IPA, 
 IQA, 
 IQB, 
 IQC, 
 IRA, 
 IRB, 
 IRC, 
 ISA, 
 ISB, 
 ISC, 
 ITA, 
 ITB, 
 ITC, 
 IUA, 
 IUB, 
 IUC, 
 IVA, 
 IVB, 
 IVC, 
 IWA, 
 IWB, 
 IWC, 
 IXA, 
 IXB, 
 IXC, 
 IYA,  
 OAA, 
 OAB, 
 OAC, 
 OAD, 
 OAE, 
 OAF, 
 OAG, 
 OAH, 
 OBA, 
 OBB, 
 OBC, 
 OBD, 
 OBE, 
 OBF, 
 OBG, 
 OBH, 
 OCA, 
 OCB, 
 OCC, 
 OCD, 
 OCE, 
 OCF, 
 OCG, 
 OCH, 
 ODA, 
 ODB, 
 ODC, 
 ODD, 
 ODE, 
 ODF, 
 ODG, 
 ODH, 
 OKA, 
 OKB, 
 OKC, 
OKD ); 
    
 input IZZ; 
 input IAA; 
 input IAB; 
 input IAC; 
 input IAD; 
 input IAE; 
 input IAF; 
 input IAG; 
 input IAH; 
 input ICA; 
 input ICB; 
 input ICC; 
 input ICD; 
 input ICE; 
 input ICF; 
 input ICG; 
 input ICH; 
 input IEA; 
 input IEB; 
 input IEC; 
 input IED; 
 input IEE; 
 input IEF; 
 input IEG; 
 input IEH; 
 input IGA; 
 input IGB; 
 input IGC; 
 input IGD; 
 input IGE; 
 input IGF; 
 input IGG; 
 input IGH; 
 input IIA; 
 input IJA; 
 input IKA; 
 input ILA; 
 input IPA; 
 input IQA; 
 input IQB; 
 input IQC; 
 input IRA; 
 input IRB; 
 input IRC; 
 input ISA; 
 input ISB; 
 input ISC; 
 input ITA; 
 input ITB; 
 input ITC; 
 input IUA; 
 input IUB; 
 input IUC; 
 input IVA; 
 input IVB; 
 input IVC; 
 input IWA; 
 input IWB; 
 input IWC; 
 input IXA; 
 input IXB; 
 input IXC; 
 input IYA;  
 output OAA; 
 output OAB; 
 output OAC; 
 output OAD; 
 output OAE; 
 output OAF; 
 output OAG; 
 output OAH; 
 output OBA; 
 output OBB; 
 output OBC; 
 output OBD; 
 output OBE; 
 output OBF; 
 output OBG; 
 output OBH; 
 output OCA; 
 output OCB; 
 output OCC; 
 output OCD; 
 output OCE; 
 output OCF; 
 output OCG; 
 output OCH; 
 output ODA; 
 output ODB; 
 output ODC; 
 output ODD; 
 output ODE; 
 output ODF; 
 output ODG; 
 output ODH; 
 output OKA; 
 output OKB; 
 output OKC; 
 output OKD; 
  
  
reg  AAA ;
reg  AAB ;
reg  AAC ;
reg  AAD ;
reg  AAE ;
reg  AAF ;
reg  AAG ;
reg  AAH ;
reg  AAI ;
reg  AAJ ;
reg  AAK ;
reg  AAL ;
reg  AAM ;
reg  AAN ;
reg  AAO ;
reg  AAP ;
reg  ABA ;
reg  ABB ;
reg  ABC ;
reg  ABD ;
reg  ABE ;
reg  ABF ;
reg  ABG ;
reg  ABH ;
reg  ABI ;
reg  ABJ ;
reg  ABK ;
reg  ABL ;
reg  ABM ;
reg  ABN ;
reg  ABO ;
reg  ABP ;
reg  ACA ;
reg  ACB ;
reg  ACC ;
reg  ACD ;
reg  ACE ;
reg  ACF ;
reg  ACG ;
reg  ACH ;
reg  ACI ;
reg  ACJ ;
reg  ACK ;
reg  ACL ;
reg  ACM ;
reg  ACN ;
reg  ACO ;
reg  ACP ;
reg  ADA ;
reg  ADB ;
reg  ADC ;
reg  ADD ;
reg  ADE ;
reg  ADF ;
reg  ADG ;
reg  ADH ;
reg  ADI ;
reg  ADJ ;
reg  ADK ;
reg  ADL ;
reg  ADM ;
reg  ADN ;
reg  ADO ;
reg  ADP ;
reg  AEA ;
reg  AEB ;
reg  AEC ;
reg  AED ;
reg  AEE ;
reg  AEF ;
reg  AEG ;
reg  AEH ;
reg  AEI ;
reg  AEJ ;
reg  AEK ;
reg  AEL ;
reg  AEM ;
reg  AEN ;
reg  AEO ;
reg  AEP ;
reg  AFA ;
reg  AFB ;
reg  AFC ;
reg  AFD ;
reg  AFE ;
reg  AFF ;
reg  AFG ;
reg  AFH ;
reg  AFI ;
reg  AFJ ;
reg  AFK ;
reg  AFL ;
reg  AFM ;
reg  AFN ;
reg  AFO ;
reg  AFP ;
reg  AGA ;
reg  AGB ;
reg  AGC ;
reg  AGD ;
reg  AGE ;
reg  AGF ;
reg  AGG ;
reg  AGH ;
reg  AGI ;
reg  AGJ ;
reg  AGK ;
reg  AGL ;
reg  AGM ;
reg  AGN ;
reg  AGO ;
reg  AGP ;
reg  AHA ;
reg  AHB ;
reg  AHC ;
reg  AHD ;
reg  AHE ;
reg  AHF ;
reg  AHG ;
reg  AHH ;
reg  AHI ;
reg  AHJ ;
reg  AHK ;
reg  AHL ;
reg  AHM ;
reg  AHN ;
reg  AHO ;
reg  AHP ;
reg  AIA ;
reg  AIB ;
reg  AIC ;
reg  AID ;
reg  AIE ;
reg  AIF ;
reg  AIG ;
reg  AIH ;
reg  AII ;
reg  AIJ ;
reg  AIK ;
reg  AIL ;
reg  AIM ;
reg  AIN ;
reg  AIO ;
reg  AIP ;
reg  AJA ;
reg  AJB ;
reg  AJC ;
reg  AJD ;
reg  AJE ;
reg  AJF ;
reg  AJG ;
reg  AJH ;
reg  AJI ;
reg  AJJ ;
reg  AJK ;
reg  AJL ;
reg  AJM ;
reg  AJN ;
reg  AJO ;
reg  AJP ;
reg  AKA ;
reg  AKB ;
reg  AKC ;
reg  AKD ;
reg  AKE ;
reg  AKF ;
reg  AKG ;
reg  AKH ;
reg  AKI ;
reg  AKJ ;
reg  AKK ;
reg  AKL ;
reg  AKM ;
reg  AKN ;
reg  AKO ;
reg  AKP ;
reg  ALA ;
reg  ALB ;
reg  ALC ;
reg  ALD ;
reg  ALE ;
reg  ALF ;
reg  ALG ;
reg  ALH ;
reg  ALI ;
reg  ALJ ;
reg  ALK ;
reg  ALL ;
reg  ALM ;
reg  ALN ;
reg  ALO ;
reg  ALP ;
reg  AMA ;
reg  AMB ;
reg  AMC ;
reg  AMD ;
reg  AME ;
reg  AMF ;
reg  AMG ;
reg  AMH ;
reg  AMI ;
reg  AMJ ;
reg  AMK ;
reg  AML ;
reg  AMM ;
reg  AMN ;
reg  AMO ;
reg  AMP ;
reg  ANA ;
reg  ANB ;
reg  ANC ;
reg  ANDD ;
reg  ANE ;
reg  ANF ;
reg  ANG ;
reg  ANH ;
reg  ANI ;
reg  ANJ ;
reg  ANK ;
reg  ANL ;
reg  ANM ;
reg  ANN ;
reg  ANO ;
reg  ANP ;
reg  AOA ;
reg  AOB ;
reg  AOC ;
reg  AOD ;
reg  AOE ;
reg  AOF ;
reg  AOG ;
reg  AOH ;
reg  AOI ;
reg  AOJ ;
reg  AOK ;
reg  AOL ;
reg  AOM ;
reg  AON ;
reg  AOO ;
reg  AOP ;
reg  APA ;
reg  APB ;
reg  APC ;
reg  APD ;
reg  APE ;
reg  APF ;
reg  APG ;
reg  APH ;
reg  API ;
reg  APJ ;
reg  APK ;
reg  APL ;
reg  APM ;
reg  APN ;
reg  APO ;
reg  APP ;
reg  CAA ;
reg  CAB ;
reg  CAC ;
reg  CAD ;
reg  CBA ;
reg  CBB ;
reg  CBC ;
reg  CBD ;
reg  CCA ;
reg  CCB ;
reg  CCC ;
reg  CCD ;
reg  CDA ;
reg  CDB ;
reg  CDC ;
reg  CDD ;
reg  CDE ;
reg  CEA ;
reg  CEB ;
reg  CEC ;
reg  CED ;
reg  CFA ;
reg  CFB ;
reg  CFC ;
reg  CFD ;
reg  CGA ;
reg  CGB ;
reg  CGC ;
reg  CGD ;
reg  CHA ;
reg  CHB ;
reg  CHC ;
reg  CHD ;
reg  EAA ;
reg  EAB ;
reg  EAC ;
reg  EAD ;
reg  EAE ;
reg  EAF ;
reg  EAG ;
reg  EAH ;
reg  EBA ;
reg  EBB ;
reg  EBC ;
reg  EBD ;
reg  EBE ;
reg  EBF ;
reg  EBG ;
reg  EBH ;
reg  ECA ;
reg  ECB ;
reg  ECC ;
reg  ECD ;
reg  ECE ;
reg  ECF ;
reg  ECG ;
reg  ECH ;
reg  EDA ;
reg  EDB ;
reg  EDC ;
reg  EDD ;
reg  EDE ;
reg  EDF ;
reg  EDG ;
reg  EDH ;
reg  EEA ;
reg  EEB ;
reg  EEC ;
reg  EED ;
reg  EEE ;
reg  EEF ;
reg  EEG ;
reg  EEH ;
reg  EFA ;
reg  EFB ;
reg  EFC ;
reg  EFD ;
reg  EFE ;
reg  EFF ;
reg  EFG ;
reg  EFH ;
reg  EGA ;
reg  EGB ;
reg  EGC ;
reg  EGD ;
reg  EGE ;
reg  EGF ;
reg  EGG ;
reg  EGH ;
reg  EHA ;
reg  EHB ;
reg  EHC ;
reg  EHD ;
reg  EHE ;
reg  EHF ;
reg  EHG ;
reg  EHH ;
reg  eia ;
reg  eib ;
reg  eic ;
reg  eid ;
reg  eie ;
reg  eif ;
reg  eig ;
reg  eih ;
reg  eja ;
reg  ejb ;
reg  ejc ;
reg  ejd ;
reg  eje ;
reg  ejf ;
reg  ejg ;
reg  ejh ;
reg  eka ;
reg  ekb ;
reg  ekc ;
reg  ekd ;
reg  eke ;
reg  ekf ;
reg  ekg ;
reg  ekh ;
reg  ela ;
reg  elb ;
reg  elc ;
reg  eld ;
reg  ele ;
reg  elf ;
reg  elg ;
reg  elh ;
reg  ema ;
reg  emb ;
reg  emc ;
reg  emd ;
reg  eme ;
reg  emf ;
reg  emg ;
reg  emh ;
reg  ena ;
reg  enb ;
reg  enc ;
reg  endd ;
reg  ene ;
reg  enf ;
reg  eng ;
reg  enh ;
reg  eoa ;
reg  eob ;
reg  eoc ;
reg  eod ;
reg  eoe ;
reg  eof ;
reg  eog ;
reg  eoh ;
reg  epa ;
reg  epb ;
reg  epc ;
reg  epd ;
reg  epe ;
reg  epf ;
reg  epg ;
reg  eph ;
reg  KAA ;
reg  KAB ;
reg  KAC ;
reg  KAD ;
reg  KBA ;
reg  KBB ;
reg  KBC ;
reg  KBD ;
reg  KBE ;
reg  KBF ;
reg  KBG ;
reg  KBH ;
reg  KCA ;
reg  KCB ;
reg  KCC ;
reg  KCD ;
reg  KCE ;
reg  KCF ;
reg  KCG ;
reg  KCH ;
reg  KDA ;
reg  KDB ;
reg  KDC ;
reg  KDD ;
reg  KDE ;
reg  KDF ;
reg  KDG ;
reg  KDH ;
reg  KEA ;
reg  KEB ;
reg  KEC ;
reg  KED ;
reg  KEE ;
reg  KEF ;
reg  KEG ;
reg  KEH ;
reg  KFA ;
reg  KFB ;
reg  KFC ;
reg  KFD ;
reg  KFE ;
reg  KFF ;
reg  KFG ;
reg  KFH ;
reg  KGA ;
reg  KGB ;
reg  KGC ;
reg  KGD ;
reg  KGE ;
reg  KGF ;
reg  KGG ;
reg  KGH ;
reg  KHA ;
reg  KHB ;
reg  KHC ;
reg  KHD ;
reg  KHE ;
reg  KHF ;
reg  KHG ;
reg  KHH ;
reg  maa ;
reg  mab ;
reg  mac ;
reg  mae ;
reg  maf ;
reg  mag ;
reg  NAA ;
reg  NAB ;
reg  NAC ;
reg  NAD ;
reg  NAE ;
reg  NAF ;
reg  NAG ;
reg  NAH ;
reg  NAI ;
reg  NAJ ;
reg  NAK ;
reg  NAL ;
reg  NAM ;
reg  NAN ;
reg  NAO ;
reg  NAP ;
reg  NBA ;
reg  NBB ;
reg  NBC ;
reg  NBD ;
reg  NBE ;
reg  NBF ;
reg  NBG ;
reg  NBH ;
reg  NBI ;
reg  NBJ ;
reg  NBK ;
reg  NBL ;
reg  NBM ;
reg  NBN ;
reg  NBO ;
reg  NBP ;
reg  nca ;
reg  ncb ;
reg  ncc ;
reg  ncd ;
reg  nce ;
reg  ncf ;
reg  ncg ;
reg  nch ;
reg  nci ;
reg  ncj ;
reg  nck ;
reg  ncl ;
reg  ncm ;
reg  ncn ;
reg  nco ;
reg  ncp ;
reg  nda ;
reg  ndb ;
reg  ndc ;
reg  ndd ;
reg  nde ;
reg  ndf ;
reg  ndg ;
reg  ndh ;
reg  nea ;
reg  neb ;
reg  nec ;
reg  ned ;
reg  nee ;
reg  nef ;
reg  neg ;
reg  neh ;
reg  nei ;
reg  nej ;
reg  nek ;
reg  nel ;
reg  nem ;
reg  nen ;
reg  neo ;
reg  nep ;
reg  nfa ;
reg  nfb ;
reg  nfc ;
reg  nfd ;
reg  nfe ;
reg  nff ;
reg  nfg ;
reg  nfh ;
reg  NGA ;
reg  NGB ;
reg  NGC ;
reg  NGD ;
reg  NGE ;
reg  NGF ;
reg  NGG ;
reg  NGH ;
reg  nha ;
reg  nhb ;
reg  nhc ;
reg  nhd ;
reg  nhe ;
reg  nhf ;
reg  nhg ;
reg  nhh ;
reg  OAA ;
reg  OAB ;
reg  OAC ;
reg  OAD ;
reg  OAE ;
reg  OAF ;
reg  OAG ;
reg  OAH ;
reg  OBA ;
reg  OBB ;
reg  OBC ;
reg  OBD ;
reg  OBE ;
reg  OBF ;
reg  OBG ;
reg  OBH ;
reg  OCA ;
reg  OCB ;
reg  OCC ;
reg  OCD ;
reg  OCE ;
reg  OCF ;
reg  OCG ;
reg  OCH ;
reg  ODA ;
reg  ODB ;
reg  ODC ;
reg  ODD ;
reg  ODE ;
reg  ODF ;
reg  ODG ;
reg  ODH ;
reg  OKA ;
reg  OKB ;
reg  OKC ;
reg  OKD ;
reg  QAF ;
reg  QCA ;
reg  QCC ;
reg  QCD ;
reg  QCE ;
reg  QCF ;
reg  QCG ;
reg  qch ;
reg  qci ;
reg  qcj ;
reg  QCL ;
reg  QCM ;
reg  qcn ;
reg  qcp ;
reg  qcq ;
reg  qcr ;
reg  qcs ;
reg  qct ;
reg  qcu ;
reg  QDA ;
reg  QDB ;
reg  QDC ;
reg  QDD ;
reg  QDE ;
reg  QDF ;
reg  qea ;
reg  qeb ;
reg  qec ;
reg  qed ;
reg  qee ;
reg  qef ;
reg  qeg ;
reg  qeh ;
reg  qfa ;
reg  qfb ;
reg  QFC ;
reg  qfg ;
reg  qfh ;
reg  qfi ;
reg  qfj ;
reg  qfk ;
reg  qfl ;
reg  qfm ;
reg  QFN ;
reg  QIA ;
reg  QIB ;
reg  QIC ;
reg  QID ;
reg  QIE ;
reg  QIF ;
reg  QIG ;
reg  QIH ;
reg  QII ;
reg  QIJ ;
reg  QIK ;
reg  QIL ;
reg  qja ;
reg  qjb ;
reg  qjc ;
reg  qka ;
reg  qkb ;
reg  qkc ;
reg  qla ;
reg  qlb ;
reg  qlc ;
reg  qma ;
reg  qmb ;
reg  qmc ;
reg  QNA ;
reg  QNB ;
reg  QNC ;
reg  QND ;
reg  QNE ;
reg  QNF ;
reg  qoa ;
reg  qob ;
reg  qoc ;
reg  qpa ;
reg  qpb ;
reg  qpc ;
reg  qpd ;
reg  qpe ;
reg  qpf ;
reg  qpg ;
reg  qph ;
reg  qpi ;
reg  qpj ;
reg  qpk ;
reg  qpl ;
reg  QQA ;
reg  qqb ;
reg  qqc ;
reg  qqd ;
reg  QUA ;
reg  QUB ;
reg  QUC ;
reg  QUD ;
reg  QVA ;
reg  QVB ;
reg  QVC ;
reg  QVD ;
reg  QVE ;
reg  QWA ;
reg  QWB ;
reg  QWC ;
reg  QXA ;
reg  QXB ;
reg  QXC ;
reg  QYA ;
reg  QYB ;
reg  QYC ;
reg  QYD ;
reg  QYE ;
reg  qza ;
reg  qzb ;
reg  qzc ;
reg  qzd ;
reg  qze ;
reg  RAA ;
reg  RAB ;
reg  RAC ;
reg  RAD ;
reg  RAE ;
reg  RAF ;
reg  RAG ;
reg  RAH ;
reg  RAI ;
reg  RAJ ;
reg  RAK ;
reg  RAL ;
reg  RAM ;
reg  RAN ;
reg  RAO ;
reg  RAP ;
reg  RBA ;
reg  RBB ;
reg  RBC ;
reg  RBD ;
reg  RBE ;
reg  RBF ;
reg  RBG ;
reg  RBH ;
reg  RBI ;
reg  RBJ ;
reg  RBK ;
reg  RBL ;
reg  RBM ;
reg  RBN ;
reg  RBO ;
reg  RBP ;
reg  rca ;
reg  rcb ;
reg  rcc ;
reg  rcd ;
reg  rce ;
reg  rcf ;
reg  rcg ;
reg  rch ;
reg  rci ;
reg  rcj ;
reg  rck ;
reg  rcl ;
reg  rcm ;
reg  rcn ;
reg  rco ;
reg  rcp ;
reg  rda ;
reg  rdb ;
reg  rdc ;
reg  rdd ;
reg  rde ;
reg  rdf ;
reg  rdg ;
reg  rdh ;
reg  RDI ;
reg  RDJ ;
reg  RDK ;
reg  RDL ;
reg  RDM ;
reg  RDN ;
reg  RDO ;
reg  RDP ;
reg  REA ;
reg  REB ;
reg  REC ;
reg  RED ;
reg  REE ;
reg  REFF ;
reg  REGG ;
reg  REH ;
reg  TAA ;
reg  TAB ;
reg  TAC ;
reg  TAD ;
reg  TAE ;
reg  TAF ;
reg  TAG ;
reg  TAH ;
reg  TAI ;
reg  TAJ ;
reg  TAK ;
reg  TAL ;
reg  TAM ;
reg  TAN ;
reg  TAO ;
reg  TAP ;
reg  TBA ;
reg  TBB ;
reg  TBC ;
reg  TBD ;
reg  TBE ;
reg  TBF ;
reg  TJA ;
reg  TJB ;
reg  TJC ;
reg  TJD ;
reg  TJE ;
reg  TJF ;
reg  tjg ;
reg  TKA ;
reg  TKB ;
reg  TKC ;
reg  TKD ;
reg  TLA ;
reg  TLB ;
reg  TLC ;
reg  TLD ;
reg  tle ;
reg  tlf ;
reg  tlg ;
reg  tlh ;
reg  TLM ;
reg  TLN ;
reg  TLO ;
reg  TLP ;
reg  TPA ;
reg  twa ;
reg  twe ;
wire  aaa ;
wire  aab ;
wire  aac ;
wire  aad ;
wire  aae ;
wire  aaf ;
wire  aag ;
wire  aah ;
wire  aai ;
wire  aaj ;
wire  aak ;
wire  aal ;
wire  aam ;
wire  aan ;
wire  aao ;
wire  aap ;
wire  aba ;
wire  abb ;
wire  abc ;
wire  abd ;
wire  abe ;
wire  abf ;
wire  abg ;
wire  abh ;
wire  abi ;
wire  abj ;
wire  abk ;
wire  abl ;
wire  abm ;
wire  abn ;
wire  abo ;
wire  abp ;
wire  aca ;
wire  acb ;
wire  acc ;
wire  acd ;
wire  ace ;
wire  acf ;
wire  acg ;
wire  ach ;
wire  aci ;
wire  acj ;
wire  ack ;
wire  acl ;
wire  acm ;
wire  acn ;
wire  aco ;
wire  acp ;
wire  ada ;
wire  adb ;
wire  adc ;
wire  add ;
wire  ade ;
wire  adf ;
wire  adg ;
wire  adh ;
wire  adi ;
wire  adj ;
wire  adk ;
wire  adl ;
wire  adm ;
wire  adn ;
wire  ado ;
wire  adp ;
wire  aea ;
wire  aeb ;
wire  aec ;
wire  aed ;
wire  aee ;
wire  aef ;
wire  aeg ;
wire  aeh ;
wire  aei ;
wire  aej ;
wire  aek ;
wire  ael ;
wire  aem ;
wire  aen ;
wire  aeo ;
wire  aep ;
wire  afa ;
wire  afb ;
wire  afc ;
wire  afd ;
wire  afe ;
wire  aff ;
wire  afg ;
wire  afh ;
wire  afi ;
wire  afj ;
wire  afk ;
wire  afl ;
wire  afm ;
wire  afn ;
wire  afo ;
wire  afp ;
wire  aga ;
wire  agb ;
wire  agc ;
wire  agd ;
wire  age ;
wire  agf ;
wire  agg ;
wire  agh ;
wire  agi ;
wire  agj ;
wire  agk ;
wire  agl ;
wire  agm ;
wire  agn ;
wire  ago ;
wire  agp ;
wire  aha ;
wire  ahb ;
wire  ahc ;
wire  ahd ;
wire  ahe ;
wire  ahf ;
wire  ahg ;
wire  ahh ;
wire  ahi ;
wire  ahj ;
wire  ahk ;
wire  ahl ;
wire  ahm ;
wire  ahn ;
wire  aho ;
wire  ahp ;
wire  aia ;
wire  aib ;
wire  aic ;
wire  aid ;
wire  aie ;
wire  aif ;
wire  aig ;
wire  aih ;
wire  aii ;
wire  aij ;
wire  aik ;
wire  ail ;
wire  aim ;
wire  ain ;
wire  aio ;
wire  aip ;
wire  aja ;
wire  ajb ;
wire  ajc ;
wire  ajd ;
wire  aje ;
wire  ajf ;
wire  ajg ;
wire  ajh ;
wire  aji ;
wire  ajj ;
wire  ajk ;
wire  ajl ;
wire  ajm ;
wire  ajn ;
wire  ajo ;
wire  ajp ;
wire  aka ;
wire  akb ;
wire  akc ;
wire  akd ;
wire  ake ;
wire  akf ;
wire  akg ;
wire  akh ;
wire  aki ;
wire  akj ;
wire  akk ;
wire  akl ;
wire  akm ;
wire  akn ;
wire  ako ;
wire  akp ;
wire  ala ;
wire  alb ;
wire  alc ;
wire  ald ;
wire  ale ;
wire  alf ;
wire  alg ;
wire  alh ;
wire  ali ;
wire  alj ;
wire  alk ;
wire  all ;
wire  alm ;
wire  aln ;
wire  alo ;
wire  alp ;
wire  ama ;
wire  amb ;
wire  amc ;
wire  amd ;
wire  ame ;
wire  amf ;
wire  amg ;
wire  amh ;
wire  ami ;
wire  amj ;
wire  amk ;
wire  aml ;
wire  amm ;
wire  amn ;
wire  amo ;
wire  amp ;
wire  ana ;
wire  anb ;
wire  anc ;
wire  andd ;
wire  ane ;
wire  anf ;
wire  ang ;
wire  anh ;
wire  ani ;
wire  anj ;
wire  ank ;
wire  anl ;
wire  anm ;
wire  ann ;
wire  ano ;
wire  anp ;
wire  aoa ;
wire  aob ;
wire  aoc ;
wire  aod ;
wire  aoe ;
wire  aof ;
wire  aog ;
wire  aoh ;
wire  aoi ;
wire  aoj ;
wire  aok ;
wire  aol ;
wire  aom ;
wire  aon ;
wire  aoo ;
wire  aop ;
wire  apa ;
wire  apb ;
wire  apc ;
wire  apd ;
wire  ape ;
wire  apf ;
wire  apg ;
wire  aph ;
wire  api ;
wire  apj ;
wire  apk ;
wire  apl ;
wire  apm ;
wire  apn ;
wire  apo ;
wire  app ;
wire  caa ;
wire  cab ;
wire  cac ;
wire  cad ;
wire  cba ;
wire  cbb ;
wire  cbc ;
wire  cbd ;
wire  cca ;
wire  ccb ;
wire  ccc ;
wire  ccd ;
wire  cda ;
wire  cdb ;
wire  cdc ;
wire  cdd ;
wire  cde ;
wire  cea ;
wire  ceb ;
wire  cec ;
wire  ced ;
wire  cfa ;
wire  cfb ;
wire  cfc ;
wire  cfd ;
wire  cga ;
wire  cgb ;
wire  cgc ;
wire  cgd ;
wire  cha ;
wire  chb ;
wire  chc ;
wire  chd ;
wire  eaa ;
wire  eab ;
wire  eac ;
wire  ead ;
wire  eae ;
wire  eaf ;
wire  eag ;
wire  eah ;
wire  eba ;
wire  ebb ;
wire  ebc ;
wire  ebd ;
wire  ebe ;
wire  ebf ;
wire  ebg ;
wire  ebh ;
wire  eca ;
wire  ecb ;
wire  ecc ;
wire  ecd ;
wire  ece ;
wire  ecf ;
wire  ecg ;
wire  ech ;
wire  eda ;
wire  edb ;
wire  edc ;
wire  edd ;
wire  ede ;
wire  edf ;
wire  edg ;
wire  edh ;
wire  eea ;
wire  eeb ;
wire  eec ;
wire  eed ;
wire  eee ;
wire  eef ;
wire  eeg ;
wire  eeh ;
wire  efa ;
wire  efb ;
wire  efc ;
wire  efd ;
wire  efe ;
wire  eff ;
wire  efg ;
wire  efh ;
wire  ega ;
wire  egb ;
wire  egc ;
wire  egd ;
wire  ege ;
wire  egf ;
wire  egg ;
wire  egh ;
wire  eha ;
wire  ehb ;
wire  ehc ;
wire  ehd ;
wire  ehe ;
wire  ehf ;
wire  ehg ;
wire  ehh ;
wire  EIA ;
wire  EIB ;
wire  EIC ;
wire  EID ;
wire  EIE ;
wire  EIF ;
wire  EIG ;
wire  EIH ;
wire  EJA ;
wire  EJB ;
wire  EJC ;
wire  EJD ;
wire  EJE ;
wire  EJF ;
wire  EJG ;
wire  EJH ;
wire  EKA ;
wire  EKB ;
wire  EKC ;
wire  EKD ;
wire  EKE ;
wire  EKF ;
wire  EKG ;
wire  EKH ;
wire  ELA ;
wire  ELB ;
wire  ELC ;
wire  ELD ;
wire  ELE ;
wire  ELF ;
wire  ELG ;
wire  ELH ;
wire  EMA ;
wire  EMB ;
wire  EMC ;
wire  EMD ;
wire  EME ;
wire  EMF ;
wire  EMG ;
wire  EMH ;
wire  ENA ;
wire  ENB ;
wire  ENC ;
wire  ENDD ;
wire  ENE ;
wire  ENF ;
wire  ENG ;
wire  ENH ;
wire  EOA ;
wire  EOB ;
wire  EOC ;
wire  EOD ;
wire  EOE ;
wire  EOF ;
wire  EOG ;
wire  EOH ;
wire  EPA ;
wire  EPB ;
wire  EPC ;
wire  EPD ;
wire  EPE ;
wire  EPF ;
wire  EPG ;
wire  EPH ;
wire  FAA ;
wire  FAB ;
wire  FAC ;
wire  FAD ;
wire  FAE ;
wire  FAF ;
wire  FAG ;
wire  FAH ;
wire  FAI ;
wire  FBA ;
wire  FBB ;
wire  FBC ;
wire  FBD ;
wire  FBE ;
wire  FBF ;
wire  FBG ;
wire  FBH ;
wire  FBI ;
wire  gab ;
wire  GAB ;
wire  gac ;
wire  GAC ;
wire  gad ;
wire  GAD ;
wire  gae ;
wire  GAE ;
wire  gbb ;
wire  GBB ;
wire  gbc ;
wire  GBC ;
wire  gbd ;
wire  GBD ;
wire  gbe ;
wire  GBE ;
wire  gcb ;
wire  GCB ;
wire  gcc ;
wire  GCC ;
wire  gcd ;
wire  GCD ;
wire  gce ;
wire  GCE ;
wire  gdb ;
wire  GDB ;
wire  gdc ;
wire  GDC ;
wire  gdd ;
wire  GDD ;
wire  gde ;
wire  GDE ;
wire  geb ;
wire  GEB ;
wire  gec ;
wire  GEC ;
wire  ged ;
wire  GED ;
wire  gee ;
wire  GEE ;
wire  gfb ;
wire  GFB ;
wire  gfc ;
wire  GFC ;
wire  gfd ;
wire  GFD ;
wire  gfe ;
wire  GFE ;
wire  ggb ;
wire  GGB ;
wire  ggc ;
wire  GGC ;
wire  ggd ;
wire  GGD ;
wire  gge ;
wire  GGE ;
wire  ghb ;
wire  GHB ;
wire  ghc ;
wire  GHC ;
wire  ghd ;
wire  GHD ;
wire  haa ;
wire  HAA ;
wire  hab ;
wire  HAB ;
wire  hac ;
wire  HAC ;
wire  had ;
wire  HAD ;
wire  hba ;
wire  HBA ;
wire  hbb ;
wire  HBB ;
wire  hbc ;
wire  HBC ;
wire  hbd ;
wire  HBD ;
wire  hca ;
wire  HCA ;
wire  hcb ;
wire  HCB ;
wire  hcc ;
wire  HCC ;
wire  hcd ;
wire  HCD ;
wire  hda ;
wire  HDA ;
wire  hdb ;
wire  HDB ;
wire  hdc ;
wire  HDC ;
wire  hdd ;
wire  HDD ;
wire  hea ;
wire  HEA ;
wire  heb ;
wire  HEB ;
wire  hec ;
wire  HEC ;
wire  hed ;
wire  HED ;
wire  hfa ;
wire  HFA ;
wire  hfb ;
wire  HFB ;
wire  hfc ;
wire  HFC ;
wire  hfd ;
wire  HFD ;
wire  hga ;
wire  HGA ;
wire  hgb ;
wire  HGB ;
wire  hgc ;
wire  HGC ;
wire  hgd ;
wire  HGD ;
wire  hha ;
wire  HHA ;
wire  hhb ;
wire  HHB ;
wire  hhc ;
wire  HHC ;
wire  hhd ;
wire  HHD ;
wire  iaa ;
wire  iab ;
wire  iac ;
wire  iad ;
wire  iae ;
wire  iaf ;
wire  iag ;
wire  iah ;
wire  ica ;
wire  icb ;
wire  icc ;
wire  icd ;
wire  ice ;
wire  icf ;
wire  icg ;
wire  ich ;
wire  iea ;
wire  ieb ;
wire  iec ;
wire  ied ;
wire  iee ;
wire  ief ;
wire  ieg ;
wire  ieh ;
wire  iga ;
wire  igb ;
wire  igc ;
wire  igd ;
wire  ige ;
wire  igf ;
wire  igg ;
wire  igh ;
wire  iia ;
wire  ija ;
wire  ika ;
wire  ila ;
wire  ipa ;
wire  iqa ;
wire  iqb ;
wire  iqc ;
wire  ira ;
wire  irb ;
wire  irc ;
wire  isa ;
wire  isb ;
wire  isc ;
wire  ita ;
wire  itb ;
wire  itc ;
wire  iua ;
wire  iub ;
wire  iuc ;
wire  iva ;
wire  ivb ;
wire  ivc ;
wire  iwa ;
wire  iwb ;
wire  iwc ;
wire  ixa ;
wire  ixb ;
wire  ixc ;
wire  iya ;
wire  izz ;
wire  jaa ;
wire  JAA ;
wire  jab ;
wire  JAB ;
wire  jac ;
wire  JAC ;
wire  jad ;
wire  JAD ;
wire  jae ;
wire  JAE ;
wire  jaf ;
wire  JAF ;
wire  jag ;
wire  JAG ;
wire  jah ;
wire  JAH ;
wire  jai ;
wire  JAI ;
wire  jaj ;
wire  JAJ ;
wire  jak ;
wire  JAK ;
wire  jal ;
wire  JAL ;
wire  jam ;
wire  JAM ;
wire  jan ;
wire  JAN ;
wire  jao ;
wire  JAO ;
wire  jap ;
wire  JAP ;
wire  jba ;
wire  JBA ;
wire  jbb ;
wire  JBB ;
wire  jbc ;
wire  JBC ;
wire  jbd ;
wire  JBD ;
wire  jbe ;
wire  JBE ;
wire  jbf ;
wire  JBF ;
wire  jbg ;
wire  JBG ;
wire  jbh ;
wire  JBH ;
wire  jbi ;
wire  JBI ;
wire  jbj ;
wire  JBJ ;
wire  jbk ;
wire  JBK ;
wire  jbl ;
wire  JBL ;
wire  jbm ;
wire  JBM ;
wire  jbn ;
wire  JBN ;
wire  jbo ;
wire  JBO ;
wire  jbp ;
wire  JBP ;
wire  jca ;
wire  JCA ;
wire  jcb ;
wire  JCB ;
wire  jcc ;
wire  JCC ;
wire  jcd ;
wire  JCD ;
wire  jce ;
wire  JCE ;
wire  jcf ;
wire  JCF ;
wire  jcg ;
wire  JCG ;
wire  jch ;
wire  JCH ;
wire  jci ;
wire  JCI ;
wire  jcj ;
wire  JCJ ;
wire  jck ;
wire  JCK ;
wire  jcl ;
wire  JCL ;
wire  jcm ;
wire  JCM ;
wire  jcn ;
wire  JCN ;
wire  jco ;
wire  JCO ;
wire  jcp ;
wire  JCP ;
wire  jda ;
wire  JDA ;
wire  jdb ;
wire  JDB ;
wire  jdc ;
wire  JDC ;
wire  jdd ;
wire  JDD ;
wire  jde ;
wire  JDE ;
wire  jdf ;
wire  JDF ;
wire  jdg ;
wire  JDG ;
wire  jdh ;
wire  JDH ;
wire  jdi ;
wire  JDI ;
wire  jdj ;
wire  JDJ ;
wire  jdk ;
wire  JDK ;
wire  jdl ;
wire  JDL ;
wire  jdm ;
wire  JDM ;
wire  jdn ;
wire  JDN ;
wire  jdo ;
wire  JDO ;
wire  jdp ;
wire  JDP ;
wire  jea ;
wire  JEA ;
wire  jeb ;
wire  JEB ;
wire  jec ;
wire  JEC ;
wire  jed ;
wire  JED ;
wire  jee ;
wire  JEE ;
wire  jef ;
wire  JEF ;
wire  jeg ;
wire  JEG ;
wire  jeh ;
wire  JEH ;
wire  jei ;
wire  JEI ;
wire  jej ;
wire  JEJ ;
wire  jek ;
wire  JEK ;
wire  jel ;
wire  JEL ;
wire  jem ;
wire  JEM ;
wire  jen ;
wire  JEN ;
wire  jeo ;
wire  JEO ;
wire  jep ;
wire  JEP ;
wire  jfa ;
wire  JFA ;
wire  jfb ;
wire  JFB ;
wire  jfc ;
wire  JFC ;
wire  jfd ;
wire  JFD ;
wire  jfe ;
wire  JFE ;
wire  jff ;
wire  JFF ;
wire  jfg ;
wire  JFG ;
wire  jfh ;
wire  JFH ;
wire  jfi ;
wire  JFI ;
wire  jfj ;
wire  JFJ ;
wire  jfk ;
wire  JFK ;
wire  jfl ;
wire  JFL ;
wire  jfm ;
wire  JFM ;
wire  jfn ;
wire  JFN ;
wire  jfo ;
wire  JFO ;
wire  jfp ;
wire  JFP ;
wire  jga ;
wire  JGA ;
wire  jgb ;
wire  JGB ;
wire  jgc ;
wire  JGC ;
wire  jgd ;
wire  JGD ;
wire  jge ;
wire  JGE ;
wire  jgf ;
wire  JGF ;
wire  jgg ;
wire  JGG ;
wire  jgh ;
wire  JGH ;
wire  jgi ;
wire  JGI ;
wire  jgj ;
wire  JGJ ;
wire  jgk ;
wire  JGK ;
wire  jgl ;
wire  JGL ;
wire  jgm ;
wire  JGM ;
wire  jgn ;
wire  JGN ;
wire  jgo ;
wire  JGO ;
wire  jgp ;
wire  JGP ;
wire  jha ;
wire  JHA ;
wire  jhb ;
wire  JHB ;
wire  jhc ;
wire  JHC ;
wire  jhd ;
wire  JHD ;
wire  jhe ;
wire  JHE ;
wire  jhf ;
wire  JHF ;
wire  jhg ;
wire  JHG ;
wire  jhh ;
wire  JHH ;
wire  jhi ;
wire  JHI ;
wire  jhj ;
wire  JHJ ;
wire  jhk ;
wire  JHK ;
wire  jhl ;
wire  JHL ;
wire  jhm ;
wire  JHM ;
wire  jhn ;
wire  JHN ;
wire  jho ;
wire  JHO ;
wire  jhp ;
wire  JHP ;
wire  kaa ;
wire  kab ;
wire  kac ;
wire  kad ;
wire  kba ;
wire  kbb ;
wire  kbc ;
wire  kbd ;
wire  kbe ;
wire  kbf ;
wire  kbg ;
wire  kbh ;
wire  kca ;
wire  kcb ;
wire  kcc ;
wire  kcd ;
wire  kce ;
wire  kcf ;
wire  kcg ;
wire  kch ;
wire  kda ;
wire  kdb ;
wire  kdc ;
wire  kdd ;
wire  kde ;
wire  kdf ;
wire  kdg ;
wire  kdh ;
wire  kea ;
wire  keb ;
wire  kec ;
wire  ked ;
wire  kee ;
wire  kef ;
wire  keg ;
wire  keh ;
wire  kfa ;
wire  kfb ;
wire  kfc ;
wire  kfd ;
wire  kfe ;
wire  kff ;
wire  kfg ;
wire  kfh ;
wire  kga ;
wire  kgb ;
wire  kgc ;
wire  kgd ;
wire  kge ;
wire  kgf ;
wire  kgg ;
wire  kgh ;
wire  kha ;
wire  khb ;
wire  khc ;
wire  khd ;
wire  khe ;
wire  khf ;
wire  khg ;
wire  khh ;
wire  MAA ;
wire  MAB ;
wire  MAC ;
wire  MAE ;
wire  MAF ;
wire  MAG ;
wire  naa ;
wire  nab ;
wire  nac ;
wire  nad ;
wire  nae ;
wire  naf ;
wire  nag ;
wire  nah ;
wire  nai ;
wire  naj ;
wire  nak ;
wire  nal ;
wire  nam ;
wire  nan ;
wire  nao ;
wire  nap ;
wire  nba ;
wire  nbb ;
wire  nbc ;
wire  nbd ;
wire  nbe ;
wire  nbf ;
wire  nbg ;
wire  nbh ;
wire  nbi ;
wire  nbj ;
wire  nbk ;
wire  nbl ;
wire  nbm ;
wire  nbn ;
wire  nbo ;
wire  nbp ;
wire  NCA ;
wire  NCB ;
wire  NCC ;
wire  NCD ;
wire  NCE ;
wire  NCF ;
wire  NCG ;
wire  NCH ;
wire  NCI ;
wire  NCJ ;
wire  NCK ;
wire  NCL ;
wire  NCM ;
wire  NCN ;
wire  NCO ;
wire  NCP ;
wire  NDA ;
wire  NDB ;
wire  NDC ;
wire  NDD ;
wire  NDE ;
wire  NDF ;
wire  NDG ;
wire  NDH ;
wire  NEA ;
wire  NEB ;
wire  NEC ;
wire  NED ;
wire  NEE ;
wire  NEF ;
wire  NEG ;
wire  NEH ;
wire  NEI ;
wire  NEJ ;
wire  NEK ;
wire  NEL ;
wire  NEM ;
wire  NEN ;
wire  NEO ;
wire  NEP ;
wire  NFA ;
wire  NFB ;
wire  NFC ;
wire  NFD ;
wire  NFE ;
wire  NFF ;
wire  NFG ;
wire  NFH ;
wire  nga ;
wire  ngb ;
wire  ngc ;
wire  ngd ;
wire  nge ;
wire  ngf ;
wire  ngg ;
wire  ngh ;
wire  NHA ;
wire  NHB ;
wire  NHC ;
wire  NHD ;
wire  NHE ;
wire  NHF ;
wire  NHG ;
wire  NHH ;
wire  oaa ;
wire  oab ;
wire  oac ;
wire  oad ;
wire  oae ;
wire  oaf ;
wire  oag ;
wire  oah ;
wire  oba ;
wire  obb ;
wire  obc ;
wire  obd ;
wire  obe ;
wire  obf ;
wire  obg ;
wire  obh ;
wire  oca ;
wire  ocb ;
wire  occ ;
wire  ocd ;
wire  oce ;
wire  ocf ;
wire  ocg ;
wire  och ;
wire  oda ;
wire  odb ;
wire  odc ;
wire  odd ;
wire  ode ;
wire  odf ;
wire  odg ;
wire  odh ;
wire  oka ;
wire  okb ;
wire  okc ;
wire  okd ;
wire  paa ;
wire  PAA ;
wire  pab ;
wire  PAB ;
wire  pac ;
wire  PAC ;
wire  pad ;
wire  PAD ;
wire  pae ;
wire  PAE ;
wire  paf ;
wire  PAF ;
wire  pag ;
wire  PAG ;
wire  pah ;
wire  PAH ;
wire  qaf ;
wire  qca ;
wire  qcc ;
wire  qcd ;
wire  qce ;
wire  qcf ;
wire  qcg ;
wire  QCH ;
wire  QCI ;
wire  QCJ ;
wire  qcl ;
wire  qcm ;
wire  QCN ;
wire  QCP ;
wire  QCQ ;
wire  QCR ;
wire  QCS ;
wire  QCT ;
wire  QCU ;
wire  qda ;
wire  qdb ;
wire  qdc ;
wire  qdd ;
wire  qde ;
wire  qdf ;
wire  QEA ;
wire  QEB ;
wire  QEC ;
wire  QED ;
wire  QEE ;
wire  QEF ;
wire  QEG ;
wire  QEH ;
wire  QFA ;
wire  QFB ;
wire  qfc ;
wire  QFG ;
wire  QFH ;
wire  QFI ;
wire  QFJ ;
wire  QFK ;
wire  QFL ;
wire  QFM ;
wire  qfn ;
wire  qhg ;
wire  QHG ;
wire  qhh ;
wire  QHH ;
wire  qhi ;
wire  QHI ;
wire  qia ;
wire  qib ;
wire  qic ;
wire  qid ;
wire  qie ;
wire  qif ;
wire  qig ;
wire  qih ;
wire  qii ;
wire  qij ;
wire  qik ;
wire  qil ;
wire  QJA ;
wire  QJB ;
wire  QJC ;
wire  QKA ;
wire  QKB ;
wire  QKC ;
wire  QLA ;
wire  QLB ;
wire  QLC ;
wire  QMA ;
wire  QMB ;
wire  QMC ;
wire  qna ;
wire  qnb ;
wire  qnc ;
wire  qnd ;
wire  qne ;
wire  qnf ;
wire  QOA ;
wire  QOB ;
wire  QOC ;
wire  QPA ;
wire  QPB ;
wire  QPC ;
wire  QPD ;
wire  QPE ;
wire  QPF ;
wire  QPG ;
wire  QPH ;
wire  QPI ;
wire  QPJ ;
wire  QPK ;
wire  QPL ;
wire  qqa ;
wire  QQB ;
wire  QQC ;
wire  QQD ;
wire  qua ;
wire  qub ;
wire  quc ;
wire  qud ;
wire  qva ;
wire  qvb ;
wire  qvc ;
wire  qvd ;
wire  qve ;
wire  qwa ;
wire  qwb ;
wire  qwc ;
wire  qxa ;
wire  qxb ;
wire  qxc ;
wire  qya ;
wire  qyb ;
wire  qyc ;
wire  qyd ;
wire  qye ;
wire  QZA ;
wire  QZB ;
wire  QZC ;
wire  QZD ;
wire  QZE ;
wire  raa ;
wire  rab ;
wire  rac ;
wire  rad ;
wire  rae ;
wire  raf ;
wire  rag ;
wire  rah ;
wire  rai ;
wire  raj ;
wire  rak ;
wire  ral ;
wire  ram ;
wire  ran ;
wire  rao ;
wire  rap ;
wire  rba ;
wire  rbb ;
wire  rbc ;
wire  rbd ;
wire  rbe ;
wire  rbf ;
wire  rbg ;
wire  rbh ;
wire  rbi ;
wire  rbj ;
wire  rbk ;
wire  rbl ;
wire  rbm ;
wire  rbn ;
wire  rbo ;
wire  rbp ;
wire  RCA ;
wire  RCB ;
wire  RCC ;
wire  RCD ;
wire  RCE ;
wire  RCF ;
wire  RCG ;
wire  RCH ;
wire  RCI ;
wire  RCJ ;
wire  RCK ;
wire  RCL ;
wire  RCM ;
wire  RCN ;
wire  RCO ;
wire  RCP ;
wire  RDA ;
wire  RDB ;
wire  RDC ;
wire  RDD ;
wire  RDE ;
wire  RDF ;
wire  RDG ;
wire  RDH ;
wire  rdi ;
wire  rdj ;
wire  rdk ;
wire  rdl ;
wire  rdm ;
wire  rdn ;
wire  rdo ;
wire  rdp ;
wire  rea ;
wire  reb ;
wire  rec ;
wire  red ;
wire  ree ;
wire  reff ;
wire  regg ;
wire  reh ;
wire  taa ;
wire  tab ;
wire  tac ;
wire  tad ;
wire  tae ;
wire  taf ;
wire  tag ;
wire  tah ;
wire  tai ;
wire  taj ;
wire  tak ;
wire  tal ;
wire  tam ;
wire  tan ;
wire  tao ;
wire  tap ;
wire  tba ;
wire  tbb ;
wire  tbc ;
wire  tbd ;
wire  tbe ;
wire  tbf ;
wire  tce ;
wire  TCE ;
wire  tcf ;
wire  TCF ;
wire  tde ;
wire  TDE ;
wire  tdf ;
wire  TDF ;
wire  tea ;
wire  TEA ;
wire  teb ;
wire  TEB ;
wire  tfe ;
wire  TFE ;
wire  tff ;
wire  TFF ;
wire  tja ;
wire  tjb ;
wire  tjc ;
wire  tjd ;
wire  tje ;
wire  tjf ;
wire  TJG ;
wire  tka ;
wire  tkb ;
wire  tkc ;
wire  tkd ;
wire  tla ;
wire  tlb ;
wire  tlc ;
wire  tld ;
wire  TLE ;
wire  TLF ;
wire  TLG ;
wire  TLH ;
wire  tlm ;
wire  tln ;
wire  tlo ;
wire  tlp ;
wire  tpa ;
wire  TWA ;
wire  TWE ;
wire  txa ;
wire  TXA ;
wire  txb ;
wire  TXB ;
wire  txc ;
wire  TXC ;
wire  txd ;
wire  TXD ;
wire  txe ;
wire  TXE ;
wire  txf ;
wire  TXF ;
wire  txg ;
wire  TXG ;
wire  txh ;
wire  TXH ;
wire  ZZI ;
wire  ZZO ;
assign ZZI = 1'b1;
assign ZZO = 1'b0;
assign GAB =  CAA  ; 
assign gab = ~GAB;  //complement 
assign GAC =  CAA & CAB  ; 
assign gac = ~GAC;  //complement 
assign caa = ~CAA;  //complement 
assign GAD =  CAA & CAB & CAC  ; 
assign gad = ~GAD;  //complement 
assign cab = ~CAB;  //complement 
assign kaa = ~KAA;  //complement 
assign GAE =  CAA & CAB & CAC & CAD  ; 
assign gae = ~GAE;  //complement 
assign kab = ~KAB;  //complement 
assign MAA = ~maa;  //complement 
assign keb = ~KEB;  //complement 
assign kef = ~KEF;  //complement 
assign kea = ~KEA;  //complement 
assign kee = ~KEE;  //complement 
assign GEE =  CEA & CEB & CEC & CED  ; 
assign gee = ~GEE;  //complement 
assign GED =  CEA & CEB & CEC  ; 
assign ged = ~GED;  //complement 
assign cea = ~CEA;  //complement 
assign MAE = ~mae;  //complement 
assign GEB =  CEA  ; 
assign geb = ~GEB;  //complement 
assign GEC =  CEA & CEB  ; 
assign gec = ~GEC;  //complement 
assign ceb = ~CEB;  //complement 
assign RCI = ~rci;  //complement 
assign RCJ = ~rcj;  //complement 
assign RDA = ~rda;  //complement 
assign RDB = ~rdb;  //complement 
assign aaa = ~AAA;  //complement 
assign aab = ~AAB;  //complement 
assign RCA = ~rca;  //complement 
assign RCB = ~rcb;  //complement 
assign aca = ~ACA;  //complement 
assign acb = ~ACB;  //complement 
assign eaa = ~EAA;  //complement 
assign eba = ~EBA;  //complement 
assign eca = ~ECA;  //complement 
assign eda = ~EDA;  //complement 
assign raa = ~RAA;  //complement 
assign rab = ~RAB;  //complement 
assign ama = ~AMA;  //complement 
assign amb = ~AMB;  //complement 
assign aea = ~AEA;  //complement 
assign aeb = ~AEB;  //complement 
assign akb = ~AKB;  //complement 
assign aga = ~AGA;  //complement 
assign agb = ~AGB;  //complement 
assign eea = ~EEA;  //complement 
assign efa = ~EFA;  //complement 
assign ega = ~EGA;  //complement 
assign eha = ~EHA;  //complement 
assign aia = ~AIA;  //complement 
assign aib = ~AIB;  //complement 
assign EIA = ~eia;  //complement 
assign EJA = ~eja;  //complement 
assign EKA = ~eka;  //complement 
assign ELA = ~ela;  //complement 
assign rba = ~RBA;  //complement 
assign rbb = ~RBB;  //complement 
assign aka = ~AKA;  //complement 
assign EMA = ~ema;  //complement 
assign ENA = ~ena;  //complement 
assign EOA = ~eoa;  //complement 
assign EPA = ~epa;  //complement 
assign aoa = ~AOA;  //complement 
assign aob = ~AOB;  //complement 
assign JAA =  AAA & EAA  |  ABA & EBA  |  ACA & ECA  |  ADA & EDA  ; 
assign jaa = ~JAA;  //complement 
assign JEA =  AAA & EAA  |  ABA & EBA  |  ACA & ECA  |  ADA & EDA  ; 
assign jea = ~JEA; //complement 
assign aba = ~ABA;  //complement 
assign abb = ~ABB;  //complement 
assign rdi = ~RDI;  //complement 
assign QJA = ~qja;  //complement 
assign QKA = ~qka;  //complement 
assign QLA = ~qla;  //complement 
assign QMA = ~qma;  //complement 
assign JAB =  AAB & EAA  |  ABB & EBA  |  ACB & ECA  |  ADB & EDA  ; 
assign jab = ~JAB;  //complement 
assign JEB =  AAB & EAA  |  ABB & EBA  |  ACB & ECA  |  ADB & EDA  ; 
assign jeb = ~JEB; //complement 
assign ada = ~ADA;  //complement 
assign adb = ~ADB;  //complement 
assign rdj = ~RDJ;  //complement 
assign qda = ~QDA;  //complement 
assign qdd = ~QDD;  //complement 
assign JBA =  AEA & EEA  |  AFA & EFA  |  AGA & EGA  |  AHA & EHA  ; 
assign jba = ~JBA;  //complement 
assign JFA =  AEA & EEA  |  AFA & EFA  |  AGA & EGA  |  AHA & EHA  ; 
assign jfa = ~JFA; //complement 
assign afa = ~AFA;  //complement 
assign afb = ~AFB;  //complement 
assign tpa = ~TPA;  //complement 
assign naa = ~NAA;  //complement 
assign JBB =  AEB & EEA  |  AFB & EFA  |  AGB & EGA  |  AHB & EHA  ; 
assign jbb = ~JBB;  //complement 
assign JFB =  AEB & EEA  |  AFB & EFA  |  AGB & EGA  |  AHB & EHA  ; 
assign jfb = ~JFB; //complement 
assign aha = ~AHA;  //complement 
assign ahb = ~AHB;  //complement 
assign rea = ~REA;  //complement 
assign reb = ~REB;  //complement 
assign NCI = ~nci;  //complement 
assign NEA = ~nea;  //complement 
assign nab = ~NAB;  //complement 
assign JCA =  AIA & EIA  |  AJA & EJA  |  AKA & EKA  |  ALA & ELA  ; 
assign jca = ~JCA;  //complement 
assign JGA =  AIA & EIA  |  AJA & EJA  |  AKA & EKA  |  ALA & ELA  ; 
assign jga = ~JGA; //complement 
assign aja = ~AJA;  //complement 
assign ajb = ~AJB;  //complement 
assign nba = ~NBA;  //complement 
assign JCB =  AIB & EIA  |  AJB & EJA  |  AKB & EKA  |  ALB & ELA  ; 
assign jcb = ~JCB;  //complement 
assign JGB =  AIB & EIA  |  AJB & EJA  |  AKB & EKA  |  ALB & ELA  ; 
assign jgb = ~JGB; //complement 
assign ala = ~ALA;  //complement 
assign alb = ~ALB;  //complement 
assign NCJ = ~ncj;  //complement 
assign NEB = ~neb;  //complement 
assign NHA = ~nha;  //complement 
assign NHB = ~nhb;  //complement 
assign nbb = ~NBB;  //complement 
assign JDA =  AMA & EMA  |  ANA & ENA  |  AOA & EOA  |  APA & EPA  ; 
assign jda = ~JDA;  //complement 
assign JHA =  AMA & EMA  |  ANA & ENA  |  AOA & EOA  |  APA & EPA  ; 
assign jha = ~JHA; //complement 
assign ana = ~ANA;  //complement 
assign anb = ~ANB;  //complement 
assign nga = ~NGA;  //complement 
assign oaa = ~OAA;  //complement 
assign oba = ~OBA;  //complement 
assign oca = ~OCA;  //complement 
assign oda = ~ODA;  //complement 
assign JDB =  AMB & EMA  |  ANB & ENA  |  AOB & EOA  |  APB & EPA  ; 
assign jdb = ~JDB;  //complement 
assign JHB =  AMB & EMA  |  ANB & ENA  |  AOB & EOA  |  APB & EPA  ; 
assign jhb = ~JHB; //complement 
assign apa = ~APA;  //complement 
assign apb = ~APB;  //complement 
assign oab = ~OAB;  //complement 
assign obb = ~OBB;  //complement 
assign ocb = ~OCB;  //complement 
assign odb = ~ODB;  //complement 
assign cac = ~CAC;  //complement 
assign cad = ~CAD;  //complement 
assign kac = ~KAC;  //complement 
assign HAA =  caa  ; 
assign haa = ~HAA;  //complement 
assign HAB =  cab  ; 
assign hab = ~HAB;  //complement 
assign HAC =  cac  ; 
assign hac = ~HAC;  //complement 
assign kad = ~KAD;  //complement 
assign HAD =  cad  ; 
assign had = ~HAD;  //complement  
assign ked = ~KED;  //complement 
assign keh = ~KEH;  //complement 
assign HED =  ced  ; 
assign hed = ~HED;  //complement  
assign kec = ~KEC;  //complement 
assign keg = ~KEG;  //complement 
assign HEA =  cea  ; 
assign hea = ~HEA;  //complement 
assign HEB =  ceb  ; 
assign heb = ~HEB;  //complement 
assign HEC =  cec  ; 
assign hec = ~HEC;  //complement 
assign pae =  TBF & QAF  ; 
assign PAE = ~pae;  //complement 
assign cec = ~CEC;  //complement 
assign ced = ~CED;  //complement 
assign RCK = ~rck;  //complement 
assign RCL = ~rcl;  //complement 
assign RDC = ~rdc;  //complement 
assign RDD = ~rdd;  //complement 
assign aac = ~AAC;  //complement 
assign aad = ~AAD;  //complement 
assign RCC = ~rcc;  //complement 
assign RCD = ~rcd;  //complement 
assign JAF =  AAF & EAC  |  ABF & EBC  |  ACF & ECC  |  ADF & EDC  ; 
assign jaf = ~JAF;  //complement 
assign acc = ~ACC;  //complement 
assign acd = ~ACD;  //complement 
assign eab = ~EAB;  //complement 
assign ebb = ~EBB;  //complement 
assign ecb = ~ECB;  //complement 
assign edb = ~EDB;  //complement 
assign rac = ~RAC;  //complement 
assign rad = ~RAD;  //complement 
assign amc = ~AMC;  //complement 
assign amd = ~AMD;  //complement 
assign aec = ~AEC;  //complement 
assign aed = ~AED;  //complement 
assign qnc = ~QNC;  //complement 
assign qnf = ~QNF;  //complement 
assign QPD = ~qpd;  //complement 
assign QPE = ~qpe;  //complement 
assign QPF = ~qpf;  //complement 
assign QPG = ~qpg;  //complement 
assign QOA = ~qoa;  //complement 
assign QOB = ~qob;  //complement 
assign QOC = ~qoc;  //complement 
assign agc = ~AGC;  //complement 
assign agd = ~AGD;  //complement 
assign eeb = ~EEB;  //complement 
assign efb = ~EFB;  //complement 
assign egb = ~EGB;  //complement 
assign ehb = ~EHB;  //complement 
assign QPH = ~qph;  //complement 
assign QPI = ~qpi;  //complement 
assign QPJ = ~qpj;  //complement 
assign QPK = ~qpk;  //complement 
assign QPA = ~qpa;  //complement 
assign QPB = ~qpb;  //complement 
assign QPC = ~qpc;  //complement 
assign QPL = ~qpl;  //complement 
assign aic = ~AIC;  //complement 
assign aid = ~AID;  //complement 
assign EIB = ~eib;  //complement 
assign EJB = ~ejb;  //complement 
assign EKB = ~ekb;  //complement 
assign ELB = ~elb;  //complement 
assign rbc = ~RBC;  //complement 
assign rbd = ~RBD;  //complement 
assign akc = ~AKC;  //complement 
assign akd = ~AKD;  //complement 
assign EMB = ~emb;  //complement 
assign ENB = ~enb;  //complement 
assign EOB = ~eob;  //complement 
assign EPB = ~epb;  //complement 
assign aoc = ~AOC;  //complement 
assign aod = ~AOD;  //complement 
assign JAC =  AAC & EAB  |  ABC & EBB  |  ACC & ECB  |  ADC & EDB  ; 
assign jac = ~JAC;  //complement 
assign JEC =  AAC & EAB  |  ABC & EBB  |  ACC & ECB  |  ADC & EDB  ; 
assign jec = ~JEC; //complement 
assign abc = ~ABC;  //complement 
assign abd = ~ABD;  //complement 
assign rdk = ~RDK;  //complement 
assign QJB = ~qjb;  //complement 
assign QKB = ~qkb;  //complement 
assign QLB = ~qlb;  //complement 
assign QMB = ~qmb;  //complement 
assign JAD =  AAD & EAB  |  ABD & EBB  |  ACD & ECB  |  ADD & EDB  ; 
assign jad = ~JAD;  //complement 
assign JED =  AAD & EAB  |  ABD & EBB  |  ACD & ECB  |  ADD & EDB  ; 
assign jed = ~JED; //complement 
assign JFC =  AAD & EAB  |  ABD & EBB  |  ACD & ECB  |  ADD & EDB  ; 
assign jfc = ~JFC;  //complement 
assign adc = ~ADC;  //complement 
assign add = ~ADD;  //complement 
assign rdl = ~RDL;  //complement 
assign qdb = ~QDB;  //complement 
assign qde = ~QDE;  //complement 
assign JBC =  AEC & EEB  |  AFC & EFB  |  AGC & EGB  |  AHC & EHB  ; 
assign jbc = ~JBC;  //complement 
assign afc = ~AFC;  //complement 
assign afd = ~AFD;  //complement 
assign nac = ~NAC;  //complement 
assign JBD =  AED & EEB  |  AFD & EFB  |  AGD & EGB  |  AHD & EHB  ; 
assign jbd = ~JBD;  //complement 
assign JFD =  AED & EEB  |  AFD & EFB  |  AGD & EGB  |  AHD & EHB  ; 
assign jfd = ~JFD; //complement 
assign ahc = ~AHC;  //complement 
assign ahd = ~AHD;  //complement 
assign rec = ~REC;  //complement 
assign red = ~RED;  //complement 
assign NCK = ~nck;  //complement 
assign NEC = ~nec;  //complement 
assign nad = ~NAD;  //complement 
assign JCC =  AIC & EIB  |  AJC & EJB  |  AKC & EKB  |  ALC & ELB  ; 
assign jcc = ~JCC;  //complement 
assign JGC =  AIC & EIB  |  AJC & EJB  |  AKC & EKB  |  ALC & ELB  ; 
assign jgc = ~JGC; //complement 
assign ajc = ~AJC;  //complement 
assign ajd = ~AJD;  //complement 
assign nbc = ~NBC;  //complement 
assign JCD =  AID & EIB  |  AJD & EJB  |  AKD & EKB  |  ALD & ELB  ; 
assign jcd = ~JCD;  //complement 
assign JGD =  AID & EIB  |  AJD & EJB  |  AKD & EKB  |  ALD & ELB  ; 
assign jgd = ~JGD; //complement 
assign alc = ~ALC;  //complement 
assign ald = ~ALD;  //complement 
assign NCL = ~ncl;  //complement 
assign NED = ~ned;  //complement 
assign NHC = ~nhc;  //complement 
assign NHD = ~nhd;  //complement 
assign nbd = ~NBD;  //complement 
assign JDC =  AMC & EMB  |  ANC & ENB  |  AOC & EOB  |  APC & EPB  ; 
assign jdc = ~JDC;  //complement 
assign JHC =  AMC & EMB  |  ANC & ENB  |  AOC & EOB  |  APC & EPB  ; 
assign jhc = ~JHC; //complement 
assign anc = ~ANC;  //complement 
assign andd = ~ANDD;  //complement 
assign ngb = ~NGB;  //complement 
assign oac = ~OAC;  //complement 
assign obc = ~OBC;  //complement 
assign occ = ~OCC;  //complement 
assign odc = ~ODC;  //complement 
assign JDD =  AMD & EMB  |  ANDD & ENB  |  AOD & EOB  |  APD & EPB  ; 
assign jdd = ~JDD;  //complement 
assign JHD =  AMD & EMB  |  ANDD & ENB  |  AOD & EOB  |  APD & EPB  ; 
assign jhd = ~JHD; //complement 
assign apc = ~APC;  //complement 
assign apd = ~APD;  //complement 
assign oad = ~OAD;  //complement 
assign obd = ~OBD;  //complement 
assign ocd = ~OCD;  //complement 
assign odd = ~ODD;  //complement 
assign GBB =  CBA  ; 
assign gbb = ~GBB;  //complement 
assign GBC =  CBA & CBB  ; 
assign gbc = ~GBC;  //complement 
assign cba = ~CBA;  //complement 
assign GBD =  CBA & CBB & CBC  ; 
assign gbd = ~GBD;  //complement 
assign cbb = ~CBB;  //complement 
assign kba = ~KBA;  //complement 
assign kbe = ~KBE;  //complement 
assign GBE =  CBA & CBB & CBC & CBD  ; 
assign gbe = ~GBE;  //complement 
assign paa =  TBE  ; 
assign PAA = ~paa;  //complement 
assign kbf = ~KBF;  //complement 
assign kbb = ~KBB;  //complement 
assign MAB = ~mab;  //complement 
assign kfb = ~KFB;  //complement 
assign kff = ~KFF;  //complement 
assign kfa = ~KFA;  //complement 
assign kfe = ~KFE;  //complement 
assign GFE =  CFA & CFB & CFC & CFD  ; 
assign gfe = ~GFE;  //complement 
assign GFD =  CFA & CFB & CFC  ; 
assign gfd = ~GFD;  //complement 
assign cfa = ~CFA;  //complement 
assign MAF = ~maf;  //complement 
assign GFB =  CFA  ; 
assign gfb = ~GFB;  //complement 
assign GFC =  CFA & CFB  ; 
assign gfc = ~GFC;  //complement 
assign cfb = ~CFB;  //complement 
assign RCM = ~rcm;  //complement 
assign RCN = ~rcn;  //complement 
assign RDE = ~rde;  //complement 
assign RDF = ~rdf;  //complement 
assign aae = ~AAE;  //complement 
assign aaf = ~AAF;  //complement 
assign qna = ~QNA;  //complement 
assign qnd = ~QND;  //complement 
assign RCE = ~rce;  //complement 
assign RCF = ~rcf;  //complement 
assign ace = ~ACE;  //complement 
assign acf = ~ACF;  //complement 
assign eac = ~EAC;  //complement 
assign ebc = ~EBC;  //complement 
assign ecc = ~ECC;  //complement 
assign edc = ~EDC;  //complement 
assign rae = ~RAE;  //complement 
assign raf = ~RAF;  //complement 
assign ame = ~AME;  //complement 
assign amf = ~AMF;  //complement 
assign aee = ~AEE;  //complement 
assign aef = ~AEF;  //complement 
assign qnb = ~QNB;  //complement 
assign qne = ~QNE;  //complement 
assign FAA = ~QDC & ~QDB & ~QDA & QCL ; 
assign FAB = ~QDC & ~QDB &  QDA & QCL ; 
assign FAC = ~QDC &  QDB & ~QDA & QCL ; 
assign FAD = ~QDC &  QDB &  QDA & QCL ; 
assign FAE =  QDC & ~QDB & ~QDA & QCL ; 
assign FAF =  QDC & ~QDB &  QDA & QCL ; 
assign FAG =  QDC &  QDB & ~QDA & QCL ; 
assign FAH =  QDC &  QDB &  QDA & QCL ; 
assign FAI = ZZI ; 
assign age = ~AGE;  //complement 
assign agf = ~AGF;  //complement 
assign eec = ~EEC;  //complement 
assign efc = ~EFC;  //complement 
assign egc = ~EGC;  //complement 
assign ehc = ~EHC;  //complement 
assign tla = ~TLA;  //complement 
assign TLE = ~tle;  //complement 
assign aie = ~AIE;  //complement 
assign aif = ~AIF;  //complement 
assign EIC = ~eic;  //complement 
assign EJC = ~ejc;  //complement 
assign EKC = ~ekc;  //complement 
assign ELC = ~elc;  //complement 
assign rbe = ~RBE;  //complement 
assign rbf = ~RBF;  //complement 
assign ake = ~AKE;  //complement 
assign akf = ~AKF;  //complement 
assign tlm = ~TLM;  //complement 
assign qia = ~QIA;  //complement 
assign qie = ~QIE;  //complement 
assign qii = ~QII;  //complement 
assign EMC = ~emc;  //complement 
assign ENC = ~enc;  //complement 
assign EOC = ~eoc;  //complement 
assign EPC = ~epc;  //complement 
assign qua = ~QUA;  //complement 
assign qub = ~QUB;  //complement 
assign quc = ~QUC;  //complement 
assign TWA = ~twa;  //complement 
assign aoe = ~AOE;  //complement 
assign aof = ~AOF;  //complement 
assign qud = ~QUD;  //complement 
assign tja = ~TJA;  //complement 
assign tka = ~TKA;  //complement 
assign JAE =  AAE & EAC  |  ABE & EBC  |  ACE & ECC  |  ADE & EDC  ; 
assign jae = ~JAE;  //complement 
assign JEE =  AAE & EAC  |  ABE & EBC  |  ACE & ECC  |  ADE & EDC  ; 
assign jee = ~JEE; //complement 
assign abe = ~ABE;  //complement 
assign abf = ~ABF;  //complement 
assign rdm = ~RDM;  //complement 
assign QJC = ~qjc;  //complement 
assign QKC = ~qkc;  //complement 
assign QLC = ~qlc;  //complement 
assign QMC = ~qmc;  //complement 
assign JEF =  AAF & EAC  |  ABF & EBC  |  ACF & ECC  |  ADF & EDC  ; 
assign jef = ~JEF;  //complement 
assign ade = ~ADE;  //complement 
assign adf = ~ADF;  //complement 
assign rdn = ~RDN;  //complement 
assign qdc = ~QDC;  //complement 
assign qdf = ~QDF;  //complement 
assign JBE =  AEE & EEC  |  AFE & EFC  |  AGE & EGC  |  AHE & EHC  ; 
assign jbe = ~JBE;  //complement 
assign JFE =  AEE & EEC  |  AFE & EFC  |  AGE & EGC  |  AHE & EHC  ; 
assign jfe = ~JFE; //complement 
assign afe = ~AFE;  //complement 
assign aff = ~AFF;  //complement 
assign oag = ~OAG;  //complement 
assign obg = ~OBG;  //complement 
assign ocg = ~OCG;  //complement 
assign odg = ~ODG;  //complement 
assign nae = ~NAE;  //complement 
assign JBF =  AEF & EEC  |  AFF & EFC  |  AGF & EGC  |  AHF & EHC  ; 
assign jbf = ~JBF;  //complement 
assign JFF =  AEF & EEC  |  AFF & EFC  |  AGF & EGC  |  AHF & EHC  ; 
assign jff = ~JFF; //complement 
assign ahe = ~AHE;  //complement 
assign ahf = ~AHF;  //complement 
assign ree = ~REE;  //complement 
assign reff = ~REFF;  //complement 
assign NCM = ~ncm;  //complement 
assign NEE = ~nee;  //complement 
assign naf = ~NAF;  //complement 
assign JCE =  AIE & EIC  |  AJE & EJC  |  AKE & EKC  |  ALE & ELC  ; 
assign jce = ~JCE;  //complement 
assign JGE =  AIE & EIC  |  AJE & EJC  |  AKE & EKC  |  ALE & ELC  ; 
assign jge = ~JGE; //complement 
assign aje = ~AJE;  //complement 
assign ajf = ~AJF;  //complement 
assign oah = ~OAH;  //complement 
assign obh = ~OBH;  //complement 
assign och = ~OCH;  //complement 
assign odh = ~ODH;  //complement 
assign nbe = ~NBE;  //complement 
assign JCF =  AIF & EIC  |  AJF & EJC  |  AKF & EKC  |  ALF & ELC  ; 
assign jcf = ~JCF;  //complement 
assign JGF =  AIF & EIC  |  AJF & EJC  |  AKF & EKC  |  ALF & ELC  ; 
assign jgf = ~JGF; //complement 
assign ale = ~ALE;  //complement 
assign alf = ~ALF;  //complement 
assign NCN = ~ncn;  //complement 
assign NEF = ~nef;  //complement 
assign NHE = ~nhe;  //complement 
assign NHF = ~nhf;  //complement 
assign nbf = ~NBF;  //complement 
assign JDE =  AME & EMC  |  ANE & ENC  |  AOE & EOC  |  APE & EPC  ; 
assign jde = ~JDE;  //complement 
assign JHE =  AME & EMC  |  ANE & ENC  |  AOE & EOC  |  APE & EPC  ; 
assign jhe = ~JHE; //complement 
assign ane = ~ANE;  //complement 
assign anf = ~ANF;  //complement 
assign ngc = ~NGC;  //complement 
assign oae = ~OAE;  //complement 
assign obe = ~OBE;  //complement 
assign oce = ~OCE;  //complement 
assign ode = ~ODE;  //complement 
assign JDF =  AMF & EMC  |  ANF & ENC  |  AOF & EOC  |  APF & EPC  ; 
assign jdf = ~JDF;  //complement 
assign JHF =  AMF & EMC  |  ANF & ENC  |  AOF & EOC  |  APF & EPC  ; 
assign jhf = ~JHF; //complement 
assign ape = ~APE;  //complement 
assign apf = ~APF;  //complement 
assign QZA = ~qza;  //complement 
assign QZB = ~qzb;  //complement 
assign QZC = ~qzc;  //complement 
assign QZD = ~qzd;  //complement 
assign oaf = ~OAF;  //complement 
assign obf = ~OBF;  //complement 
assign ocf = ~OCF;  //complement 
assign odf = ~ODF;  //complement 
assign cbc = ~CBC;  //complement 
assign cbd = ~CBD;  //complement 
assign kbc = ~KBC;  //complement 
assign kbg = ~KBG;  //complement 
assign HBA =  cba  ; 
assign hba = ~HBA;  //complement 
assign HBB =  cbb  ; 
assign hbb = ~HBB;  //complement 
assign HBC =  cbc  ; 
assign hbc = ~HBC;  //complement 
assign pab =  TBE & MAA  ; 
assign PAB = ~pab;  //complement 
assign kbd = ~KBD;  //complement 
assign kbh = ~KBH;  //complement 
assign HBD =  cbd  ; 
assign hbd = ~HBD;  //complement  
assign kfd = ~KFD;  //complement 
assign kfh = ~KFH;  //complement 
assign HFD =  cfd  ; 
assign hfd = ~HFD;  //complement  
assign kfc = ~KFC;  //complement 
assign kfg = ~KFG;  //complement 
assign HFA =  cfa  ; 
assign hfa = ~HFA;  //complement 
assign HFB =  cfb  ; 
assign hfb = ~HFB;  //complement 
assign HFC =  cfc  ; 
assign hfc = ~HFC;  //complement 
assign paf =  TBF & QAF & MAE  ; 
assign PAF = ~paf;  //complement 
assign cfc = ~CFC;  //complement 
assign cfd = ~CFD;  //complement 
assign NHG = ~nhg;  //complement 
assign NHH = ~nhh;  //complement 
assign aag = ~AAG;  //complement 
assign aah = ~AAH;  //complement 
assign taa = ~TAA;  //complement 
assign tab = ~TAB;  //complement 
assign tac = ~TAC;  //complement 
assign tad = ~TAD;  //complement 
assign RCO = ~rco;  //complement 
assign RCP = ~rcp;  //complement 
assign RDG = ~rdg;  //complement 
assign RDH = ~rdh;  //complement 
assign acg = ~ACG;  //complement 
assign ach = ~ACH;  //complement 
assign ead = ~EAD;  //complement 
assign ebd = ~EBD;  //complement 
assign ecd = ~ECD;  //complement 
assign edd = ~EDD;  //complement 
assign rag = ~RAG;  //complement 
assign rah = ~RAH;  //complement 
assign amg = ~AMG;  //complement 
assign amh = ~AMH;  //complement 
assign aeg = ~AEG;  //complement 
assign aeh = ~AEH;  //complement 
assign tae = ~TAE;  //complement 
assign taf = ~TAF;  //complement 
assign tag = ~TAG;  //complement 
assign tah = ~TAH;  //complement 
assign NEG = ~neg;  //complement 
assign NEH = ~neh;  //complement 
assign RCG = ~rcg;  //complement 
assign RCH = ~rch;  //complement 
assign agg = ~AGG;  //complement 
assign agh = ~AGH;  //complement 
assign eed = ~EED;  //complement 
assign efd = ~EFD;  //complement 
assign egd = ~EGD;  //complement 
assign ehd = ~EHD;  //complement 
assign FBA = ~QDF & ~QDE & ~QDD & QCM ; 
assign FBB = ~QDF & ~QDE &  QDD & QCM ; 
assign FBC = ~QDF &  QDE & ~QDD & QCM ; 
assign FBD = ~QDF &  QDE &  QDD & QCM ; 
assign FBE =  QDF & ~QDE & ~QDD & QCM ; 
assign FBF =  QDF & ~QDE &  QDD & QCM ; 
assign FBG =  QDF &  QDE & ~QDD & QCM ; 
assign FBH =  QDF &  QDE &  QDD & QCM ; 
assign FBI = ZZI ; 
assign aig = ~AIG;  //complement 
assign aih = ~AIH;  //complement 
assign EID = ~eid;  //complement 
assign EJD = ~ejd;  //complement 
assign EKD = ~ekd;  //complement 
assign ELD = ~eld;  //complement 
assign rbg = ~RBG;  //complement 
assign rbh = ~RBH;  //complement 
assign akg = ~AKG;  //complement 
assign akh = ~AKH;  //complement 
assign tai = ~TAI;  //complement 
assign taj = ~TAJ;  //complement 
assign tak = ~TAK;  //complement 
assign tal = ~TAL;  //complement 
assign EMD = ~emd;  //complement 
assign ENDD = ~endd;  //complement 
assign EOD = ~eod;  //complement 
assign EPD = ~epd;  //complement 
assign aog = ~AOG;  //complement 
assign aoh = ~AOH;  //complement 
assign tam = ~TAM;  //complement 
assign tan = ~TAN;  //complement 
assign tao = ~TAO;  //complement 
assign tap = ~TAP;  //complement 
assign JAG =  AAG & EAD  |  ABG & EBD  |  ACG & ECD  |  ADG & EDD  ; 
assign jag = ~JAG;  //complement 
assign JEG =  AAG & EAD  |  ABG & EBD  |  ACG & ECD  |  ADG & EDD  ; 
assign jeg = ~JEG; //complement 
assign abg = ~ABG;  //complement 
assign abh = ~ABH;  //complement 
assign rdo = ~RDO;  //complement 
assign oka = ~OKA;  //complement 
assign JAH =  AAH & EAD  |  ABH & EBD  |  ACH & ECD  |  ADH & EDD  ; 
assign jah = ~JAH;  //complement 
assign JEH =  AAH & EAD  |  ABH & EBD  |  ACH & ECD  |  ADH & EDD  ; 
assign jeh = ~JEH; //complement 
assign adg = ~ADG;  //complement 
assign adh = ~ADH;  //complement 
assign rdp = ~RDP;  //complement 
assign tje = ~TJE;  //complement 
assign tjf = ~TJF;  //complement 
assign TJG = ~tjg;  //complement 
assign JBG =  AEG & EED  |  AFG & EFD  |  AGG & EGD  |  AHG & EHD  ; 
assign jbg = ~JBG;  //complement 
assign JFG =  AEG & EED  |  AFG & EFD  |  AGG & EGD  |  AHG & EHD  ; 
assign jfg = ~JFG; //complement 
assign afg = ~AFG;  //complement 
assign afh = ~AFH;  //complement 
assign nag = ~NAG;  //complement 
assign JBH =  AEH & EED  |  AFH & EFD  |  AGH & EGD  |  AHH & EHD  ; 
assign jbh = ~JBH;  //complement 
assign JFH =  AEH & EED  |  AFH & EFD  |  AGH & EGD  |  AHH & EHD  ; 
assign jfh = ~JFH; //complement 
assign ahg = ~AHG;  //complement 
assign ahh = ~AHH;  //complement 
assign regg = ~REGG;  //complement 
assign reh = ~REH;  //complement 
assign NCO = ~nco;  //complement 
assign NCP = ~ncp;  //complement 
assign nah = ~NAH;  //complement 
assign JCG =  AIG & EID  |  AJG & EJD  |  AKG & EKD  |  ALG & ELD  ; 
assign jcg = ~JCG;  //complement 
assign JGG =  AIG & EID  |  AJG & EJD  |  AKG & EKD  |  ALG & ELD  ; 
assign jgg = ~JGG; //complement 
assign ajg = ~AJG;  //complement 
assign ajh = ~AJH;  //complement 
assign nbg = ~NBG;  //complement 
assign JCH =  AIH & EID  |  AJH & EJD  |  AKH & EKD  |  ALH & ELD  ; 
assign jch = ~JCH;  //complement 
assign JGH =  AIH & EID  |  AJH & EJD  |  AKH & EKD  |  ALH & ELD  ; 
assign jgh = ~JGH; //complement 
assign alg = ~ALG;  //complement 
assign alh = ~ALH;  //complement 
assign nbh = ~NBH;  //complement 
assign JDG =  AMG & EMD  |  ANG & ENDD |  AOG & EOD  |  APG & EPD  ; 
assign jdg = ~JDG;  //complement 
assign JHG =  AMG & EMD  |  ANG & ENDD |  AOG & EOD  |  APG & EPD  ; 
assign jhg = ~JHG; //complement 
assign ang = ~ANG;  //complement 
assign anh = ~ANH;  //complement 
assign ngd = ~NGD;  //complement 
assign qhh =  qie & qif & qig & qih  ; 
assign QHH = ~qhh;  //complement  
assign qhi =  qie & qif & qig & qih  ; 
assign QHI = ~qhi;  //complement 
assign JDH =  AMH & EMD  |  ANH & ENDD |  AOH & EOD  |  APH & EPD  ; 
assign jdh = ~JDH;  //complement 
assign JHH =  AMH & EMD  |  ANH & ENDD |  AOH & EOD  |  APH & EPD  ; 
assign jhh = ~JHH; //complement 
assign apg = ~APG;  //complement 
assign aph = ~APH;  //complement 
assign GCB =  CCA  ; 
assign gcb = ~GCB;  //complement 
assign GCC =  CCA & CCB  ; 
assign gcc = ~GCC;  //complement 
assign cca = ~CCA;  //complement 
assign GCD =  CCA & CCB & CCC  ; 
assign gcd = ~GCD;  //complement 
assign ccb = ~CCB;  //complement 
assign kca = ~KCA;  //complement 
assign kce = ~KCE;  //complement 
assign GCE =  CCA & CCB & CCC & CCD  ; 
assign gce = ~GCE;  //complement 
assign tbe = ~TBE;  //complement 
assign tbf = ~TBF;  //complement 
assign kcb = ~KCB;  //complement 
assign kcf = ~KCF;  //complement 
assign MAC = ~mac;  //complement 
assign kgb = ~KGB;  //complement 
assign kgf = ~KGF;  //complement 
assign kga = ~KGA;  //complement 
assign kge = ~KGE;  //complement 
assign GGE =  CGA & CGB & CGC & CGD  ; 
assign gge = ~GGE;  //complement 
assign GGD =  CGA & CGB & CGC  ; 
assign ggd = ~GGD;  //complement 
assign cga = ~CGA;  //complement 
assign MAG = ~mag;  //complement 
assign GGB =  CGA  ; 
assign ggb = ~GGB;  //complement 
assign GGC =  CGA & CGB  ; 
assign ggc = ~GGC;  //complement 
assign cgb = ~CGB;  //complement 
assign aai = ~AAI;  //complement 
assign aaj = ~AAJ;  //complement 
assign QCQ = ~qcq;  //complement 
assign QFM = ~qfm;  //complement 
assign aci = ~ACI;  //complement 
assign acj = ~ACJ;  //complement 
assign eae = ~EAE;  //complement 
assign ebe = ~EBE;  //complement 
assign ece = ~ECE;  //complement 
assign ede = ~EDE;  //complement 
assign rai = ~RAI;  //complement 
assign raj = ~RAJ;  //complement 
assign ami = ~AMI;  //complement 
assign amj = ~AMJ;  //complement 
assign aei = ~AEI;  //complement 
assign aej = ~AEJ;  //complement 
assign tba = ~TBA;  //complement 
assign tbb = ~TBB;  //complement 
assign tbc = ~TBC;  //complement 
assign tbd = ~TBD;  //complement 
assign QFG = ~qfg;  //complement 
assign QFH = ~qfh;  //complement 
assign QFI = ~qfi;  //complement 
assign QFJ = ~qfj;  //complement 
assign QCS = ~qcs;  //complement 
assign QCT = ~qct;  //complement 
assign QFK = ~qfk;  //complement 
assign QFL = ~qfl;  //complement 
assign agi = ~AGI;  //complement 
assign agj = ~AGJ;  //complement 
assign eee = ~EEE;  //complement 
assign efe = ~EFE;  //complement 
assign ege = ~EGE;  //complement 
assign ehe = ~EHE;  //complement 
assign QCR = ~qcr;  //complement 
assign QCU = ~qcu;  //complement 
assign qfn = ~QFN;  //complement 
assign aii = ~AII;  //complement 
assign aij = ~AIJ;  //complement 
assign EIE = ~eie;  //complement 
assign EJE = ~eje;  //complement 
assign EKE = ~eke;  //complement 
assign ELE = ~ele;  //complement 
assign rbi = ~RBI;  //complement 
assign rbj = ~RBJ;  //complement 
assign TXA =  QCQ  ; 
assign txa = ~TXA;  //complement 
assign TXC =  QCS  ; 
assign txc = ~TXC;  //complement 
assign TXE =  QCQ  ; 
assign txe = ~TXE;  //complement 
assign aki = ~AKI;  //complement 
assign akj = ~AKJ;  //complement 
assign qca = ~QCA;  //complement 
assign QFA = ~qfa;  //complement 
assign EME = ~eme;  //complement 
assign ENE = ~ene;  //complement 
assign EOE = ~eoe;  //complement 
assign EPE = ~epe;  //complement 
assign TXB =  QCR  ; 
assign txb = ~TXB;  //complement 
assign TXF =  QCU  ; 
assign txf = ~TXF;  //complement 
assign aoi = ~AOI;  //complement 
assign aoj = ~AOJ;  //complement 
assign TXD =  QCT  ; 
assign txd = ~TXD;  //complement 
assign TXG =  QCS  ; 
assign txg = ~TXG;  //complement 
assign TXH =  QCT  ; 
assign txh = ~TXH;  //complement 
assign JAI =  AAI & EAE  |  ABI & EBE  |  ACI & ECE  |  ADI & EDE  ; 
assign jai = ~JAI;  //complement 
assign JEI =  AAI & EAE  |  ABI & EBE  |  ACI & ECE  |  ADI & EDE  ; 
assign jei = ~JEI; //complement 
assign abi = ~ABI;  //complement 
assign abj = ~ABJ;  //complement 
assign QEA = ~qea;  //complement 
assign QEB = ~qeb;  //complement 
assign JAJ =  AAJ & EAE  |  ABJ & EBE  |  ACJ & ECE  |  ADJ & EDE  ; 
assign jaj = ~JAJ;  //complement 
assign JEJ =  AAJ & EAE  |  ABJ & EBE  |  ACJ & ECE  |  ADJ & EDE  ; 
assign jej = ~JEJ; //complement 
assign adi = ~ADI;  //complement 
assign adj = ~ADJ;  //complement 
assign okb = ~OKB;  //complement 
assign JBI =  AEI & EEE  |  AFI & EFE  |  AGI & EGE  |  AHI & EHE  ; 
assign jbi = ~JBI;  //complement 
assign JFI =  AEI & EEE  |  AFI & EFE  |  AGI & EGE  |  AHI & EHE  ; 
assign jfi = ~JFI; //complement 
assign afi = ~AFI;  //complement 
assign afj = ~AFJ;  //complement 
assign NCA = ~nca;  //complement 
assign QZE = ~qze;  //complement 
assign nai = ~NAI;  //complement 
assign JBJ =  AEJ & EEE  |  AFJ & EFE  |  AGJ & EGE  |  AHJ & EHE  ; 
assign jbj = ~JBJ;  //complement 
assign JFJ =  AEJ & EEE  |  AFJ & EFE  |  AGJ & EGE  |  AHJ & EHE  ; 
assign jfj = ~JFJ; //complement 
assign ahi = ~AHI;  //complement 
assign ahj = ~AHJ;  //complement 
assign NCB = ~ncb;  //complement 
assign NDA = ~nda;  //complement 
assign NDB = ~ndb;  //complement 
assign NEI = ~nei;  //complement 
assign naj = ~NAJ;  //complement 
assign JCI =  AII & EIE  |  AJI & EJE  |  AKI & EKE  |  ALI & ELE  ; 
assign jci = ~JCI;  //complement 
assign JGI =  AII & EIE  |  AJI & EJE  |  AKI & EKE  |  ALI & ELE  ; 
assign jgi = ~JGI; //complement 
assign aji = ~AJI;  //complement 
assign ajj = ~AJJ;  //complement 
assign NEJ = ~nej;  //complement 
assign NFA = ~nfa;  //complement 
assign NFB = ~nfb;  //complement 
assign nbi = ~NBI;  //complement 
assign JCJ =  AIJ & EIE  |  AJJ & EJE  |  AKJ & EKE  |  ALJ & ELE  ; 
assign jcj = ~JCJ;  //complement 
assign JGJ =  AIJ & EIE  |  AJJ & EJE  |  AKJ & EKE  |  ALJ & ELE  ; 
assign jgj = ~JGJ; //complement 
assign ali = ~ALI;  //complement 
assign alj = ~ALJ;  //complement 
assign qhg =  qie & qif & qig & qih  ; 
assign QHG = ~qhg;  //complement  
assign nbj = ~NBJ;  //complement 
assign JDI =  AMI & EME  |  ANI & ENE  |  AOI & EOE  |  API & EPE  ; 
assign jdi = ~JDI;  //complement 
assign JHI =  AMI & EME  |  ANI & ENE  |  AOI & EOE  |  API & EPE  ; 
assign jhi = ~JHI; //complement 
assign ani = ~ANI;  //complement 
assign anj = ~ANJ;  //complement 
assign nge = ~NGE;  //complement 
assign qib = ~QIB;  //complement 
assign qif = ~QIF;  //complement 
assign qij = ~QIJ;  //complement 
assign JDJ =  AMJ & EME  |  ANJ & ENE  |  AOJ & EOE  |  APJ & EPE  ; 
assign jdj = ~JDJ;  //complement 
assign JHJ =  AMJ & EME  |  ANJ & ENE  |  AOJ & EOE  |  APJ & EPE  ; 
assign jhj = ~JHJ; //complement 
assign api = ~API;  //complement 
assign apj = ~APJ;  //complement 
assign qic = ~QIC;  //complement 
assign qig = ~QIG;  //complement 
assign qik = ~QIK;  //complement 
assign ccc = ~CCC;  //complement 
assign ccd = ~CCD;  //complement 
assign kcc = ~KCC;  //complement 
assign kcg = ~KCG;  //complement 
assign HCA =  cca  ; 
assign hca = ~HCA;  //complement 
assign HCB =  ccb  ; 
assign hcb = ~HCB;  //complement 
assign HCC =  ccc  ; 
assign hcc = ~HCC;  //complement 
assign pac =  TBE & MAA & MAB  ; 
assign PAC = ~pac;  //complement 
assign kcd = ~KCD;  //complement 
assign kch = ~KCH;  //complement 
assign HCD =  ccd  ; 
assign hcd = ~HCD;  //complement  
assign kgd = ~KGD;  //complement 
assign kgh = ~KGH;  //complement 
assign HGD =  cgd  ; 
assign hgd = ~HGD;  //complement  
assign kgc = ~KGC;  //complement 
assign kgg = ~KGG;  //complement 
assign HGA =  cga  ; 
assign hga = ~HGA;  //complement 
assign HGB =  cgb  ; 
assign hgb = ~HGB;  //complement 
assign HGC =  cgc  ; 
assign hgc = ~HGC;  //complement 
assign pag =  TBF & QAF & MAE & MAF  ; 
assign PAG = ~pag;  //complement 
assign cgc = ~CGC;  //complement 
assign cgd = ~CGD;  //complement 
assign aak = ~AAK;  //complement 
assign aal = ~AAL;  //complement 
assign ack = ~ACK;  //complement 
assign acl = ~ACL;  //complement 
assign eaf = ~EAF;  //complement 
assign ebf = ~EBF;  //complement 
assign ecf = ~ECF;  //complement 
assign edf = ~EDF;  //complement 
assign rak = ~RAK;  //complement 
assign ral = ~RAL;  //complement 
assign amk = ~AMK;  //complement 
assign aml = ~AML;  //complement 
assign aek = ~AEK;  //complement 
assign ael = ~AEL;  //complement 
assign TCE = TLM; 
assign tce = ~TCE; //complement 
assign TCF = TLM; 
assign tcf = ~TCF;  //complement 
assign TDE = TLN; 
assign tde = ~TDE;  //complement 
assign TDF = TLN; 
assign tdf = ~TDF;  //complement 
assign agk = ~AGK;  //complement 
assign agl = ~AGL;  //complement 
assign eef = ~EEF;  //complement 
assign eff = ~EFF;  //complement 
assign egf = ~EGF;  //complement 
assign ehf = ~EHF;  //complement 
assign QCP = ~qcp;  //complement 
assign qcc = ~QCC;  //complement 
assign qcd = ~QCD;  //complement 
assign aik = ~AIK;  //complement 
assign ail = ~AIL;  //complement 
assign EIF = ~eif;  //complement 
assign EJF = ~ejf;  //complement 
assign EKF = ~ekf;  //complement 
assign ELF = ~elf;  //complement 
assign rbk = ~RBK;  //complement 
assign rbl = ~RBL;  //complement 
assign akk = ~AKK;  //complement 
assign akl = ~AKL;  //complement 
assign qfc = ~QFC;  //complement 
assign qcg = ~QCG;  //complement 
assign EMF = ~emf;  //complement 
assign ENF = ~enf;  //complement 
assign EOF = ~eof;  //complement 
assign EPF = ~epf;  //complement 
assign aok = ~AOK;  //complement 
assign aol = ~AOL;  //complement 
assign QCH = ~qch;  //complement 
assign QFB = ~qfb;  //complement 
assign JAK =  AAK & EAF  |  ABK & EBF  |  ACK & ECF  |  ADK & EDF  ; 
assign jak = ~JAK;  //complement 
assign JEK =  AAK & EAF  |  ABK & EBF  |  ACK & ECF  |  ADK & EDF  ; 
assign jek = ~JEK; //complement 
assign abk = ~ABK;  //complement 
assign abl = ~ABL;  //complement 
assign QEC = ~qec;  //complement 
assign QED = ~qed;  //complement 
assign JAL =  AAL & EAF  |  ABL & EBF  |  ACL & ECF  |  ADL & EDF  ; 
assign jal = ~JAL;  //complement 
assign JEL =  AAL & EAF  |  ABL & EBF  |  ACL & ECF  |  ADL & EDF  ; 
assign jel = ~JEL; //complement 
assign adk = ~ADK;  //complement 
assign adl = ~ADL;  //complement 
assign JBK =  AEK & EEF  |  AFK & EFF  |  AGK & EGF  |  AHK & EHF  ; 
assign jbk = ~JBK;  //complement 
assign JFK =  AEK & EEF  |  AFK & EFF  |  AGK & EGF  |  AHK & EHF  ; 
assign jfk = ~JFK; //complement 
assign afk = ~AFK;  //complement 
assign afl = ~AFL;  //complement 
assign okc = ~OKC;  //complement 
assign nak = ~NAK;  //complement 
assign JBL =  AEL & EEF  |  AFL & EFF  |  AGL & EGF  |  AHL & EHF  ; 
assign jbl = ~JBL;  //complement 
assign JFL =  AEL & EEF  |  AFL & EFF  |  AGL & EGF  |  AHL & EHF  ; 
assign jfl = ~JFL; //complement 
assign ahk = ~AHK;  //complement 
assign ahl = ~AHL;  //complement 
assign NCC = ~ncc;  //complement 
assign NCD = ~ncd;  //complement 
assign NDC = ~ndc;  //complement 
assign NDD = ~ndd;  //complement 
assign nal = ~NAL;  //complement 
assign JCK =  AIK & EIF  |  AJK & EJF  |  AKK & EKF  |  ALK & ELF  ; 
assign jck = ~JCK;  //complement 
assign JGK =  AIK & EIF  |  AJK & EJF  |  AKK & EKF  |  ALK & ELF  ; 
assign jgk = ~JGK; //complement 
assign ajk = ~AJK;  //complement 
assign ajl = ~AJL;  //complement 
assign okd = ~OKD;  //complement 
assign nbk = ~NBK;  //complement 
assign JCL =  AIL & EIF  |  AJL & EJF  |  AKL & EKF  |  ALL & ELF  ; 
assign jcl = ~JCL;  //complement 
assign JGL =  AIL & EIF  |  AJL & EJF  |  AKL & EKF  |  ALL & ELF  ; 
assign jgl = ~JGL; //complement 
assign alk = ~ALK;  //complement 
assign all = ~ALL;  //complement 
assign NEK = ~nek;  //complement 
assign NEL = ~nel;  //complement 
assign NFC = ~nfc;  //complement 
assign NFD = ~nfd;  //complement 
assign nbl = ~NBL;  //complement 
assign JDK =  AMK & EMF  |  ANK & ENF  |  AOK & EOF  |  APK & EPF  ; 
assign jdk = ~JDK;  //complement 
assign JHK =  AMK & EMF  |  ANK & ENF  |  AOK & EOF  |  APK & EPF  ; 
assign jhk = ~JHK; //complement 
assign ank = ~ANK;  //complement 
assign anl = ~ANL;  //complement 
assign ngf = ~NGF;  //complement 
assign qid = ~QID;  //complement 
assign qih = ~QIH;  //complement 
assign qil = ~QIL;  //complement 
assign JDL =  AML & EMF  |  ANL & ENF  |  AOL & EOF  |  APL & EPF  ; 
assign jdl = ~JDL;  //complement 
assign JHL =  AML & EMF  |  ANL & ENF  |  AOL & EOF  |  APL & EPF  ; 
assign jhl = ~JHL; //complement 
assign apk = ~APK;  //complement 
assign apl = ~APL;  //complement 
assign TWE = ~twe;  //complement 
assign GDB =  CDA  ; 
assign gdb = ~GDB;  //complement 
assign GDC =  CDA & CDB  ; 
assign gdc = ~GDC;  //complement 
assign cda = ~CDA;  //complement 
assign cde = ~CDE;  //complement 
assign GDD =  CDA & CDB & CDC  ; 
assign gdd = ~GDD;  //complement 
assign cdb = ~CDB;  //complement 
assign kda = ~KDA;  //complement 
assign kde = ~KDE;  //complement 
assign GDE =  CDE & CDB & CDC & CDD  ; 
assign gde = ~GDE;  //complement 
assign kdb = ~KDB;  //complement 
assign kdf = ~KDF;  //complement 
assign khb = ~KHB;  //complement 
assign khf = ~KHF;  //complement 
assign qaf = ~QAF;  //complement 
assign kha = ~KHA;  //complement 
assign khe = ~KHE;  //complement 
assign GHD =  CHA & CHB & CHC  ; 
assign ghd = ~GHD;  //complement 
assign cha = ~CHA;  //complement 
assign GHB =  CHA  ; 
assign ghb = ~GHB;  //complement 
assign GHC =  CHA & CHB  ; 
assign ghc = ~GHC;  //complement 
assign chb = ~CHB;  //complement 
assign aam = ~AAM;  //complement 
assign aan = ~AAN;  //complement 
assign acm = ~ACM;  //complement 
assign acn = ~ACN;  //complement 
assign eag = ~EAG;  //complement 
assign ebg = ~EBG;  //complement 
assign ecg = ~ECG;  //complement 
assign edg = ~EDG;  //complement 
assign ram = ~RAM;  //complement 
assign ran = ~RAN;  //complement 
assign amm = ~AMM;  //complement 
assign amn = ~AMN;  //complement 
assign aem = ~AEM;  //complement 
assign aen = ~AEN;  //complement 
assign agm = ~AGM;  //complement 
assign agn = ~AGN;  //complement 
assign eeg = ~EEG;  //complement 
assign efg = ~EFG;  //complement 
assign egg = ~EGG;  //complement 
assign ehg = ~EHG;  //complement 
assign aim = ~AIM;  //complement 
assign ain = ~AIN;  //complement 
assign EIG = ~eig;  //complement 
assign EJG = ~ejg;  //complement 
assign EKG = ~ekg;  //complement 
assign ELG = ~elg;  //complement 
assign rbm = ~RBM;  //complement 
assign rbn = ~RBN;  //complement 
assign akm = ~AKM;  //complement 
assign akn = ~AKN;  //complement 
assign tln = ~TLN;  //complement 
assign tlo = ~TLO;  //complement 
assign EMG = ~emg;  //complement 
assign ENG = ~eng;  //complement 
assign EOG = ~eog;  //complement 
assign EPG = ~epg;  //complement 
assign aon = ~AON;  //complement 
assign aom = ~AOM;  //complement 
assign qce = ~QCE;  //complement 
assign qcf = ~QCF;  //complement 
assign JAM =  AAM & EAG  |  ABM & EBG  |  ACM & ECG  |  ADM & EDG  ; 
assign jam = ~JAM;  //complement 
assign JEM =  AAM & EAG  |  ABM & EBG  |  ACM & ECG  |  ADM & EDG  ; 
assign jem = ~JEM; //complement 
assign abm = ~ABM;  //complement 
assign abn = ~ABN;  //complement 
assign tlb = ~TLB;  //complement 
assign QEE = ~qee;  //complement 
assign QEF = ~qef;  //complement 
assign JAN =  AAN & EAG  |  ABN & EBG  |  ACN & ECG  |  ADN & EDG  ; 
assign jan = ~JAN;  //complement 
assign JEN =  AAN & EAG  |  ABN & EBG  |  ACN & ECG  |  ADN & EDG  ; 
assign jen = ~JEN; //complement 
assign adm = ~ADM;  //complement 
assign adn = ~ADN;  //complement 
assign TLF = ~tlf;  //complement 
assign TEA = TLO; 
assign tea = ~TEA; //complement 
assign TEB = TLO; 
assign teb = ~TEB;  //complement 
assign JBM =  AEM & EEG  |  AFM & EFG  |  AGM & EGG  |  AHM & EHG  ; 
assign jbm = ~JBM;  //complement 
assign JFM =  AEM & EEG  |  AFM & EFG  |  AGM & EGG  |  AHM & EHG  ; 
assign jfm = ~JFM; //complement 
assign afm = ~AFM;  //complement 
assign afn = ~AFN;  //complement 
assign tjb = ~TJB;  //complement 
assign tkb = ~TKB;  //complement 
assign nam = ~NAM;  //complement 
assign JBN =  AEN & EEG  |  AFN & EFG  |  AGN & EGG  |  AHN & EHG  ; 
assign jbn = ~JBN;  //complement 
assign JFN =  AEN & EEG  |  AFN & EFG  |  AGN & EGG  |  AHN & EHG  ; 
assign jfn = ~JFN; //complement 
assign ahm = ~AHM;  //complement 
assign ahn = ~AHN;  //complement 
assign NCE = ~nce;  //complement 
assign NCF = ~ncf;  //complement 
assign NDE = ~nde;  //complement 
assign NDF = ~ndf;  //complement 
assign nan = ~NAN;  //complement 
assign JCM =  AIM & EIG  |  AJM & EJG  |  AKM & EKG  |  ALM & ELG  ; 
assign jcm = ~JCM;  //complement 
assign JGM =  AIM & EIG  |  AJM & EJG  |  AKM & EKG  |  ALM & ELG  ; 
assign jgm = ~JGM; //complement 
assign ajm = ~AJM;  //complement 
assign ajn = ~AJN;  //complement 
assign TFE = TLP; 
assign tfe = ~TFE; //complement 
assign TFF = TLP; 
assign tff = ~TFF;  //complement 
assign nbm = ~NBM;  //complement 
assign JCN =  AIN & EIG  |  AJN & EJG  |  AKN & EKG  |  ALN & ELG  ; 
assign jcn = ~JCN;  //complement 
assign JGN =  AIN & EIG  |  AJN & EJG  |  AKN & EKG  |  ALN & ELG  ; 
assign jgn = ~JGN; //complement 
assign alm = ~ALM;  //complement 
assign aln = ~ALN;  //complement 
assign NEM = ~nem;  //complement 
assign NEN = ~nen;  //complement 
assign NFE = ~nfe;  //complement 
assign NFF = ~nff;  //complement 
assign nbn = ~NBN;  //complement 
assign JDM =  AMM & EMG  |  ANM & ENG  |  AOM & EOG  |  APM & EPG  ; 
assign jdm = ~JDM;  //complement 
assign JHM =  AMM & EMG  |  ANM & ENG  |  AOM & EOG  |  APM & EPG  ; 
assign jhm = ~JHM; //complement 
assign anm = ~ANM;  //complement 
assign ann = ~ANN;  //complement 
assign ngg = ~NGG;  //complement 
assign QCI = ~qci;  //complement 
assign QCJ = ~qcj;  //complement 
assign QCN = ~qcn;  //complement 
assign JDN =  AMN & EMG  |  ANN & ENG  |  AON & EOG  |  APN & EPG  ; 
assign jdn = ~JDN;  //complement 
assign JHN =  AMN & EMG  |  ANN & ENG  |  AON & EOG  |  APN & EPG  ; 
assign jhn = ~JHN; //complement 
assign apm = ~APM;  //complement 
assign apn = ~APN;  //complement 
assign qcl = ~QCL;  //complement 
assign qcm = ~QCM;  //complement 
assign cdc = ~CDC;  //complement 
assign cdd = ~CDD;  //complement 
assign kdc = ~KDC;  //complement 
assign kdg = ~KDG;  //complement 
assign HDA =  cda  ; 
assign hda = ~HDA;  //complement 
assign HDB =  cdb  ; 
assign hdb = ~HDB;  //complement 
assign HDC =  cdc  ; 
assign hdc = ~HDC;  //complement 
assign pad =  TBE & MAA & MAB & MAC  ; 
assign PAD = ~pad;  //complement 
assign kdd = ~KDD;  //complement 
assign kdh = ~KDH;  //complement 
assign HDD =  cdd  ; 
assign hdd = ~HDD;  //complement  
assign chc = ~CHC;  //complement 
assign khd = ~KHD;  //complement 
assign khh = ~KHH;  //complement 
assign HHD =  chd  ; 
assign hhd = ~HHD;  //complement  
assign khc = ~KHC;  //complement 
assign khg = ~KHG;  //complement 
assign HHA =  cha  ; 
assign hha = ~HHA;  //complement 
assign HHB =  chb  ; 
assign hhb = ~HHB;  //complement 
assign HHC =  chc  ; 
assign hhc = ~HHC;  //complement 
assign pah =  TBF & QAF & MAE & MAF & MAG  ; 
assign PAH = ~pah;  //complement 
assign chd = ~CHD;  //complement 
assign qyd = ~QYD;  //complement 
assign aao = ~AAO;  //complement 
assign aap = ~AAP;  //complement 
assign qyb = ~QYB;  //complement 
assign qyc = ~QYC;  //complement 
assign qye = ~QYE;  //complement 
assign aco = ~ACO;  //complement 
assign acp = ~ACP;  //complement 
assign eah = ~EAH;  //complement 
assign ebh = ~EBH;  //complement 
assign ech = ~ECH;  //complement 
assign edh = ~EDH;  //complement 
assign rao = ~RAO;  //complement 
assign rap = ~RAP;  //complement 
assign amo = ~AMO;  //complement 
assign amp = ~AMP;  //complement 
assign aeo = ~AEO;  //complement 
assign tlc = ~TLC;  //complement 
assign qya = ~QYA;  //complement 
assign ago = ~AGO;  //complement 
assign agp = ~AGP;  //complement 
assign eeh = ~EEH;  //complement 
assign efh = ~EFH;  //complement 
assign egh = ~EGH;  //complement 
assign ehh = ~EHH;  //complement 
assign aio = ~AIO;  //complement 
assign aip = ~AIP;  //complement 
assign EIH = ~eih;  //complement 
assign EJH = ~ejh;  //complement 
assign EKH = ~ekh;  //complement 
assign ELH = ~elh;  //complement 
assign rbo = ~RBO;  //complement 
assign rbp = ~RBP;  //complement 
assign ako = ~AKO;  //complement 
assign akp = ~AKP;  //complement 
assign aep = ~AEP;  //complement 
assign tlp = ~TLP;  //complement 
assign EMH = ~emh;  //complement 
assign ENH = ~enh;  //complement 
assign EOH = ~eoh;  //complement 
assign EPH = ~eph;  //complement 
assign aoo = ~AOO;  //complement 
assign aop = ~AOP;  //complement 
assign tld = ~TLD;  //complement 
assign JAO =  AAO & EAH  |  ABO & EBH  |  ACO & ECH  |  ADO & EDH  ; 
assign jao = ~JAO;  //complement 
assign JEO =  AAO & EAH  |  ABO & EBH  |  ACO & ECH  |  ADO & EDH  ; 
assign jeo = ~JEO; //complement 
assign abo = ~ABO;  //complement 
assign abp = ~ABP;  //complement 
assign TLG = ~tlg;  //complement 
assign QEG = ~qeg;  //complement 
assign QEH = ~qeh;  //complement 
assign JAP =  AAP & EAH  |  ABP & EBH  |  ACP & ECH  |  ADP & EDH  ; 
assign jap = ~JAP;  //complement 
assign JEP =  AAP & EAH  |  ABP & EBH  |  ACP & ECH  |  ADP & EDH  ; 
assign jep = ~JEP; //complement 
assign ado = ~ADO;  //complement 
assign adp = ~ADP;  //complement 
assign qve = ~QVE;  //complement 
assign qwa = ~QWA;  //complement 
assign qwb = ~QWB;  //complement 
assign qwc = ~QWC;  //complement 
assign qva = ~QVA;  //complement 
assign qvb = ~QVB;  //complement 
assign qvc = ~QVC;  //complement 
assign qvd = ~QVD;  //complement 
assign JBO =  AEO & EEH  |  AFO & EFH  |  AGO & EGH  |  AHO & EHH  ; 
assign jbo = ~JBO;  //complement 
assign JFO =  AEO & EEH  |  AFO & EFH  |  AGO & EGH  |  AHO & EHH  ; 
assign jfo = ~JFO; //complement 
assign afo = ~AFO;  //complement 
assign afp = ~AFP;  //complement 
assign tjc = ~TJC;  //complement 
assign tkc = ~TKC;  //complement 
assign nao = ~NAO;  //complement 
assign JBP =  AEP & EEH  |  AFP & EFH  |  AGP & EGH  |  AHP & EHH  ; 
assign jbp = ~JBP;  //complement 
assign JFP =  AEP & EEH  |  AFP & EFH  |  AGP & EGH  |  AHP & EHH  ; 
assign jfp = ~JFP; //complement 
assign aho = ~AHO;  //complement 
assign ahp = ~AHP;  //complement 
assign NCG = ~ncg;  //complement 
assign NCH = ~nch;  //complement 
assign NDG = ~ndg;  //complement 
assign NDH = ~ndh;  //complement 
assign nap = ~NAP;  //complement 
assign JCO =  AIO & EIH  |  AJO & EJH  |  AKO & EKH  |  ALO & ELH  ; 
assign jco = ~JCO;  //complement 
assign JGO =  AIO & EIH  |  AJO & EJH  |  AKO & EKH  |  ALO & ELH  ; 
assign jgo = ~JGO; //complement 
assign ajo = ~AJO;  //complement 
assign ajp = ~AJP;  //complement 
assign NEO = ~neo;  //complement 
assign NEP = ~nep;  //complement 
assign NFG = ~nfg;  //complement 
assign NFH = ~nfh;  //complement 
assign nbo = ~NBO;  //complement 
assign JCP =  AIP & EIH  |  AJP & EJH  |  AKP & EKH  |  ALP & ELH  ; 
assign jcp = ~JCP;  //complement 
assign JGP =  AIP & EIH  |  AJP & EJH  |  AKP & EKH  |  ALP & ELH  ; 
assign jgp = ~JGP; //complement 
assign alo = ~ALO;  //complement 
assign alp = ~ALP;  //complement 
assign tjd = ~TJD;  //complement 
assign tkd = ~TKD;  //complement 
assign nbp = ~NBP;  //complement 
assign JDO =  AMO & EMH  |  ANO & ENH  |  AOO & EOH  |  APO & EPH  ; 
assign jdo = ~JDO;  //complement 
assign JHO =  AMO & EMH  |  ANO & ENH  |  AOO & EOH  |  APO & EPH  ; 
assign jho = ~JHO; //complement 
assign ano = ~ANO;  //complement 
assign anp = ~ANP;  //complement 
assign ngh = ~NGH;  //complement 
assign qqa = ~QQA;  //complement 
assign qxa = ~QXA;  //complement 
assign qxb = ~QXB;  //complement 
assign qxc = ~QXC;  //complement 
assign JDP =  AMP & EMH  |  ANP & ENH  |  AOP & EOH  |  APP & EPH  ; 
assign jdp = ~JDP;  //complement 
assign JHP =  AMP & EMH  |  ANP & ENH  |  AOP & EOH  |  APP & EPH  ; 
assign jhp = ~JHP; //complement 
assign apo = ~APO;  //complement 
assign app = ~APP;  //complement 
assign TLH = ~tlh;  //complement 
assign QQB = ~qqb;  //complement 
assign QQC = ~qqc;  //complement 
assign QQD = ~qqd;  //complement 
assign iaa = ~IAA; //complement 
assign iab = ~IAB; //complement 
assign iac = ~IAC; //complement 
assign iad = ~IAD; //complement 
assign iae = ~IAE; //complement 
assign iaf = ~IAF; //complement 
assign iag = ~IAG; //complement 
assign iah = ~IAH; //complement 
assign ica = ~ICA; //complement 
assign icb = ~ICB; //complement 
assign icc = ~ICC; //complement 
assign icd = ~ICD; //complement 
assign ice = ~ICE; //complement 
assign icf = ~ICF; //complement 
assign icg = ~ICG; //complement 
assign ich = ~ICH; //complement 
assign iea = ~IEA; //complement 
assign ieb = ~IEB; //complement 
assign iec = ~IEC; //complement 
assign ied = ~IED; //complement 
assign iee = ~IEE; //complement 
assign ief = ~IEF; //complement 
assign ieg = ~IEG; //complement 
assign ieh = ~IEH; //complement 
assign iga = ~IGA; //complement 
assign igb = ~IGB; //complement 
assign igc = ~IGC; //complement 
assign igd = ~IGD; //complement 
assign ige = ~IGE; //complement 
assign igf = ~IGF; //complement 
assign igg = ~IGG; //complement 
assign igh = ~IGH; //complement 
assign iia = ~IIA; //complement 
assign ija = ~IJA; //complement 
assign ika = ~IKA; //complement 
assign ila = ~ILA; //complement 
assign ipa = ~IPA; //complement 
assign iqa = ~IQA; //complement 
assign iqb = ~IQB; //complement 
assign iqc = ~IQC; //complement 
assign ira = ~IRA; //complement 
assign irb = ~IRB; //complement 
assign irc = ~IRC; //complement 
assign isa = ~ISA; //complement 
assign isb = ~ISB; //complement 
assign isc = ~ISC; //complement 
assign ita = ~ITA; //complement 
assign itb = ~ITB; //complement 
assign itc = ~ITC; //complement 
assign iua = ~IUA; //complement 
assign iub = ~IUB; //complement 
assign iuc = ~IUC; //complement 
assign iva = ~IVA; //complement 
assign ivb = ~IVB; //complement 
assign ivc = ~IVC; //complement 
assign iwa = ~IWA; //complement 
assign iwb = ~IWB; //complement 
assign iwc = ~IWC; //complement 
assign ixa = ~IXA; //complement 
assign ixb = ~IXB; //complement 
assign ixc = ~IXC; //complement 
assign iya = ~IYA; //complement 
assign izz = ~IZZ; //complement 
always@(posedge IZZ )
   begin 
 CAA <=  JAA  |  JBA  ; 
 CAB <=  JAB  |  JBB  ; 
 KAA <=  HAA  ; 
 KAB <=  gab & hab  |  GAB & HAB  ; 
 maa <= gae ; 
 KEB <=  geb & heb  |  GEB & HEB  ; 
 KEF <=  TBD & heb  ; 
 KEA <=  HEA & hea  ; 
 KEE <=  TBC & hea  ; 
 CEA <=  JCA  |  JDA  ; 
 mae <= gee ; 
 CEB <=  JCB  |  JDB  ; 
 rci <= rda ; 
 rcj <= rdb ; 
 rda <= rdi ; 
 rdb <= rdj ; 
 AAA <=  RAA & TAA  |  RCA & TAA  |  AAA & taa  ; 
 AAB <=  RAB & TAA  |  RCB & TAA  |  AAB & taa  ; 
 rca <= rci ; 
 rcb <= rcj ; 
 ACA <=  RAA & TAC  |  RCA & TAC  |  ACA & tac  ; 
 ACB <=  RAB & TAC  |  RCB & TAC  |  ACB & tac  ; 
 EAA <= QEA ; 
 EBA <= QEB ; 
 ECA <= QEC ; 
 EDA <= QED ; 
 RAA <=  KAA & paa  ; 
 RAB <=  KAB & paa  ; 
 AMA <=  RBA & TAM  |  RDA & TAM  |  AMA & tam  ; 
 AMB <=  RBB & TAM  |  RDB & TAM  |  AMB & tam  ; 
 AEA <=  RAA & TAE  |  RCA & TAE  |  AEA & tae  ; 
 AEB <=  RAB & TAE  |  RCB & TAE  |  AEB & tae  ; 
 AKB <=  RBB & TAK  |  RDB & TAK  |  AKB & tak  ; 
 AGA <=  RAA & TAG  |  RCA & TAG  |  AGA & tag  ; 
 AGB <=  RAB & TAG  |  RCB & TAG  |  AGB & tag  ; 
 EEA <= QEE ; 
 EFA <= QEF ; 
 EGA <= QEG ; 
 EHA <= QEH ; 
 AIA <=  RBA & TAI  |  RDA & TAI  |  AIA & tai  ; 
 AIB <=  RBB & TAI  |  RDB & TAI  |  AIB & tai  ; 
 eia <= qea ; 
 eja <= qeb ; 
 eka <= qec ; 
 ela <= qed ; 
 RBA <=  KEA & pae  |  KEE & PAE  ; 
 RBB <=  KEB & pae  |  KEF & PAE  ; 
 AKA <=  RBA & TAK  |  RDA & TAK  |  AKA & tak  ; 
 ema <= qee ; 
 ena <= qef ; 
 eoa <= QEG ; 
 epa <= QEH ; 
 AOA <=  RBA & TAO  |  RDA & TAO  |  AOA & tao  ; 
 AOB <=  RBB & TAO  |  RDB & TAO  |  AOB & tao  ; 
 ABA <=  RAA & TAB  |  RCA & TAB  |  ABA & tab  ; 
 ABB <=  RAB & TAB  |  RCB & TAB  |  ABB & tab  ; 
 RDI <=  REA & TCE  |  ICA & TDE  |  IEA & TEA  |  IGA & TFE  ; 
 qja <= iga ; 
 qka <= ira ; 
 qla <= isa ; 
 qma <= ita ; 
 ADA <=  RAA & TAD  |  RCA & TAD  |  ADA & tad  ; 
 ADB <=  RAB & TAD  |  RCB & TAD  |  ADB & tad  ; 
 RDJ <=  REB & TCF  |  ICB & TDF  |  IEB & TEB  |  IGB & TFF  ; 
 QDA <= QPD & QYD |  QPJ & qyd ; 
 QDD <= QPD & QYD |  QPJ & qyd ; 
 AFA <=  RAA & TAF  |  RCA & TAF  |  AFA & taf  ; 
 AFB <=  RAB & TAF  |  RCB & TAF  |  AFB & taf  ; 
 TPA <= TJE ; 
 NAA <=  JEA  |  JFA  ; 
 AHA <=  RAA & TAH  |  RCA & TAH  |  AHA & tah  ; 
 AHB <=  RAB & TAH  |  RCB & TAH  |  AHB & tah  ; 
 REA <= IAA ; 
 REB <= IAB ; 
 nci <= nba ; 
 nea <= nci ; 
 NAB <=  JEB  |  JFB  ; 
 AJA <=  RBA & TAJ  |  RDA & TAJ  |  AJA & taj  ; 
 AJB <=  RBB & TAJ  |  RDB & TAJ  |  AJB & taj  ; 
 NBA <=  JGA  |  JHA  ; 
 ALA <=  RBA & TAL  |  RDA & TAL  |  ALA & tal  ; 
 ALB <=  RBB & TAL  |  RDB & TAL  |  ALB & tal  ; 
 ncj <= nbb ; 
 neb <= ncj ; 
 nha <= nga ; 
 nhb <= ngb ; 
 NBB <=  JGB  |  JHB  ; 
 ANA <=  RBA & TAN  |  RDA & TAN  |  AMA & tan  ; 
 ANB <=  RBB & TAN  |  RDB & TAN  |  ANB & tan  ; 
 NGA <=  TXA & NAA  |  TXB & NCA  |  TXC & NEA  |  TXD & NFA  ; 
 OAA <= NHA ; 
 OBA <= NGA ; 
 OCA <= NGA ; 
 ODA <= NGA ; 
 APA <=  RBA & TAP  |  RDA & TAP  |  APA & tap  ; 
 APB <=  RBB & TAP  |  RDB & TAP  |  APB & tap  ; 
 OAB <= NHB ; 
 OBB <= NGB ; 
 OCB <= NGB ; 
 ODB <= NGB ; 
 CAC <=  JAC  |  JBC  ; 
 CAD <=  JAD  |  JBD  ; 
 KAC <=  gac & hac  |  GAC & HAC  ; 
 KAD <=  gad & had  |  GAD & HAD  ; 
 KED <=  ged & hed  |  GED & HED  ; 
 KEH <=  TBD & hed  ; 
 KEC <=  gec & hec  |  GEC & HEC  ; 
 KEG <=  TBC & hec  ; 
 CEC <=  JCC  |  JDC  ; 
 CED <=  JCD  |  JDD  ; 
 rck <= rdc ; 
 rcl <= rdd ; 
 rdc <= rdk ; 
 rdd <= rdl ; 
 AAC <=  RAC & TAA  |  RCC & TAA  |  AAC & taa  ; 
 AAD <=  RAD & TAA  |  RCD & TAA  |  AAD & taa  ; 
 rcc <= rck ; 
 rcd <= rcl ; 
 ACC <=  RAC & TAC  |  RCC & TAC  |  ACC & tac  ; 
 ACD <=  RAD & TAC  |  RCD & TAC  |  ACD & tac  ; 
 EAB <= QEA ; 
 EBB <= QEB ; 
 ECB <= QEC ; 
 EDB <= QED ; 
 RAC <=  KAC & paa  ; 
 RAD <=  KAD & paa  ; 
 AMC <=  RBC & TAM  |  RDC & TAM  |  AMC & tam  ; 
 AMD <=  RBD & TAM  |  RDD & TAM  |  AMD & tam  ; 
 AEC <=  RAC & TAE  |  RCC & TAE  |  AEC & tae  ; 
 AED <=  RAD & TAE  |  RCD & TAE  |  AED & tae  ; 
 QNC <=  QJC & TKA  |  QKC & TKB  |  QLC & TKC  |  QMC & TKD  ; 
 QNF <=  QJC & TKA  |  QKC & TKB  |  QLC & TKC  |  QMC & TKD  ; 
 qpd <= qpa ; 
 qpe <= qpb ; 
 qpf <= qpc ; 
 qpg <= qpd ; 
 qoa <= qnd ; 
 qob <= qne ; 
 qoc <= qnf ; 
 AGC <=  RAC & TAG  |  RCC & TAG  |  AGC & tag  ; 
 AGD <=  RAD & TAG  |  RCD & TAG  |  AGD & tag  ; 
 EEB <= QEE ; 
 EFB <= QEF ; 
 EGB <= QEG ; 
 EHB <= QEH ; 
 qph <= qpe ; 
 qpi <= qpf ; 
 qpj <= qpg ; 
 qpk <= qph ; 
 qpa <= qoa ; 
 qpb <= qob ; 
 qpc <= qoc ; 
 qpl <= qpi ; 
 AIC <=  RBC & TAI  |  RDC & TAI  |  AIC & tai  ; 
 AID <=  RBD & TAI  |  RDD & TAI  |  AID & tai  ; 
 eib <= qea ; 
 ejb <= qeb ; 
 ekb <= qec ; 
 elb <= qed ; 
 RBC <=  KEC & pae  |  KEG & PAE  ; 
 RBD <=  KED & pae  |  KEH & PAE  ; 
 AKC <=  RBC & TAK  |  RDC & TAK  |  AKC & tak  ; 
 AKD <=  RBD & TAK  |  RDD & TAK  |  AKD & tak  ; 
 emb <= qee ; 
 enb <= qef ; 
 eob <= QEG ; 
 epb <= QEH ; 
 AOC <=  RBC & TAO  |  RDC & TAO  |  AOC & tao  ; 
 AOD <=  RBD & TAO  |  RDD & TAO  |  AOD & tao  ; 
 ABC <=  RAC & TAB  |  RCC & TAB  |  ABC & tab  ; 
 ABD <=  RAD & TAB  |  RCD & TAB  |  ABD & tab  ; 
 RDK <=  REC & TCE  |  ICC & TDE  |  IEC & TEA  |  IGC & TFE  ; 
 qjb <= igb ; 
 qkb <= irb ; 
 qlb <= isb ; 
 qmb <= itb ; 
 ADC <=  RAC & TAD  |  RCC & TAD  |  ADC & tad  ; 
 ADD <=  RAD & TAD  |  RCD & TAD  |  ADD & tad  ; 
 RDL <=  RED & TCF  |  ICD & TDF  |  IED & TEB  |  IGD & TFF  ; 
 QDB <= QPE & QYD |  QPK & qyd ; 
 QDE <= QPE & QYD |  QPK & qyd ; 
 AFC <=  RAC & TAF  |  RCC & TAF  |  AFC & taf  ; 
 AFD <=  RAD & TAF  |  RCD & TAF  |  AFD & taf  ; 
 NAC <=  JEC  |  JFC  ; 
 AHC <=  RAC & TAH  |  RCC & TAH  |  AHC & tah  ; 
 AHD <=  RAD & TAH  |  RCD & TAH  |  AHD & tah  ; 
 REC <= IAC ; 
 RED <= IAD ; 
 nck <= nbc ; 
 nec <= nck ; 
 NAD <=  JED  |  JFD  ; 
 AJC <=  RBC & TAJ  |  RDC & TAJ  |  AJC & taj  ; 
 AJD <=  RBD & TAJ  |  RDD & TAJ  |  AJD & taj  ; 
 NBC <=  JGC  |  JHC  ; 
 ALC <=  RBC & TAL  |  RDC & TAL  |  ALC & tal  ; 
 ALD <=  RBD & TAL  |  RDD & TAL  |  ALD & tal  ; 
 ncl <= nbd ; 
 ned <= ncl ; 
 nhc <= ngc ; 
 nhd <= ngd ; 
 NBD <=  JGD  |  JHD  ; 
 ANC <=  RBC & TAN  |  RDC & TAN  |  ANC & tan  ; 
 ANDD <=  RBD & TAN  |  RDD & TAN  |  ANDD & tan  ; 
 NGB <=  TXA & NAB  |  TXB & NCB  |  TXC & NEB  |  TXD & NFB  ; 
 OAC <= NHC ; 
 OBC <= NGC ; 
 OCC <= NGC ; 
 ODC <= NGC ; 
 APC <=  RBC & TAP  |  RDC & TAP  |  APC & tap  ; 
 APD <=  RBD & TAP  |  RDD & TAP  |  APD & tap  ; 
 OAD <= NHD ; 
 OBD <= NGD ; 
 OCD <= NGD ; 
 ODD <= NGD ; 
 CBA <=  JAE  |  JBE  ; 
 CBB <=  JAF  |  JBF  ; 
 KBA <=  HBA & hba  ; 
 KBE <=  TBA & hba  ; 
 KBF <=  TBB & hbb  ; 
 KBB <=  gbb & hbb  |  GBB & HBB  ; 
 mab <= gbe ; 
 KFB <=  gfb & hfb  |  GFB & HFB  ; 
 KFF <=  TBD & hfb  ; 
 KFA <=  HFA & hfa  ; 
 KFE <=  TBC & hfa  ; 
 CFA <=  JCE  |  JDE  ; 
 maf <= gfe ; 
 CFB <=  JCF  |  JDF  ; 
 rcm <= rde ; 
 rcn <= rdf ; 
 rde <= rdm ; 
 rdf <= rdn ; 
 AAE <=  RAE & TAA  |  RCE & TAA  |  AAE & taa  ; 
 AAF <=  RAF & TAA  |  RCF & TAA  |  AAF & taa  ; 
 QNA <=  QJA & TKA  |  QKA & TKB  |  QLA & TKC  |  QMA & TKD  ; 
 QND <=  QJA & TKA  |  QKA & TKB  |  QLA & TKC  |  QMA & TKD  ; 
 rce <= rcm ; 
 rcf <= rcn ; 
 ACE <=  RAE & TAC  |  RCE & TAC  |  ACE & tac  ; 
 ACF <=  RAF & TAC  |  RCF & TAC  |  ACF & tac  ; 
 EAC <= QEA ; 
 EBC <= QEB ; 
 ECC <= QEC ; 
 EDC <= QED ; 
 RAE <=  KBA & pab  |  KBE & PAB  ; 
 RAF <=  KBB & pab  |  KBF & PAB  ; 
 AME <=  RBE & TAM  |  RDE & TAM  |  AME & tam  ; 
 AMF <=  RBF & TAM  |  RDF & TAM  |  AMF & tam  ; 
 AEE <=  RAE & TAE  |  RCE & TAE  |  AEE & tae  ; 
 AEF <=  RAF & TAE  |  RCF & TAE  |  AEF & tae  ; 
 QNB <=  QJB & TKA  |  QKB & TKB  |  QLB & TKC  |  QMB & TKD  ; 
 QNE <=  QJB & TKA  |  QKB & TKB  |  QLB & TKC  |  QMB & TKD  ; 
 AGE <=  RAE & TAG  |  RCE & TAG  |  AGE & tag  ; 
 AGF <=  RAF & TAG  |  RCF & TAG  |  AGF & tag  ; 
 EEC <= QEE ; 
 EFC <= QEF ; 
 EGC <= QEG ; 
 EHC <= QEH ; 
 TLA <= QUA & quc |  ZZO & QUC ; 
 tle <= tla ; 
 AIE <=  RBE & TAI  |  RDE & TAI  |  AIE & tai  ; 
 AIF <=  RBF & TAI  |  RDF & TAI  |  AIF & tai  ; 
 eic <= qea ; 
 ejc <= qeb ; 
 ekc <= qec ; 
 elc <= qed ; 
 RBE <=  KFA & paf  |  KFE & PAF  ; 
 RBF <=  KFB & paf  |  KFF & PAF  ; 
 AKE <=  RBE & TAK  |  RDE & TAK  |  AKE & tak  ; 
 AKF <=  RBF & TAK  |  RDF & TAK  |  AKF & tak  ; 
 TLM <=  TLM & qcn  |  TLE  ; 
 QIA <=  QQA & qhh & IIA  |  QIA & twa  ; 
 QIE <=  QQA & qhh & IIA  |  QIA & twa  ; 
 QII <=  QQA & qhh & IIA  |  QIA & twa  ; 
 emc <= qee ; 
 enc <= qef ; 
 eoc <= QEG ; 
 epc <= QEH ; 
 QUA <= IUA ; 
 QUB <= IUB ; 
 QUC <= IUC ; 
 twa <= qfn ; 
 AOE <=  RBE & TAO  |  RDE & TAO  |  AOE & tao  ; 
 AOF <=  RBF & TAO  |  RDF & TAO  |  AOF & tao  ; 
 QUD <= IUC ; 
 TJA <= QII ; 
 TKA <= QII ; 
 ABE <=  RAE & TAB  |  RCE & TAB  |  ABE & tab  ; 
 ABF <=  RAF & TAB  |  RCF & TAB  |  ABF & tab  ; 
 RDM <=  REE & TCE  |  ICE & TDE  |  IEE & TEA  |  IGE & TFE  ; 
 qjc <= igc ; 
 qkc <= irc ; 
 qlc <= isc ; 
 qmc <= itc ; 
 ADE <=  RAE & TAD  |  RCE & TAD  |  ADE & tad  ; 
 ADF <=  RAF & TAD  |  RCF & TAD  |  ADF & tad  ; 
 RDN <=  REFF & TCF  |  ICF & TDF  |  IEF & TEB  |  IGF & TFF  ; 
 QDC <= QPF & QYD |  QPL & qyd ; 
 QDF <= QPF & QYD |  QPL & qyd ; 
 AFE <=  RAE & TAF  |  RCE & TAF  |  AFE & taf  ; 
 AFF <=  RAF & TAF  |  RCF & TAF  |  AFF & taf  ; 
 OAG <= NHG ; 
 OBG <= NGG ; 
 OCG <= NGG ; 
 ODG <= NGG ; 
 NAE <=  JEE  |  JFE  ; 
 AHE <=  RAE & TAH  |  RCE & TAH  |  AHE & tah  ; 
 AHF <=  RAF & TAH  |  RCF & TAH  |  AHF & tah  ; 
 REE <= IAE ; 
 REFF <= IAF ; 
 ncm <= nbe ; 
 nee <= ncm ; 
 NAF <=  JEF  |  JFF  ; 
 AJE <=  RBE & TAJ  |  RDE & TAJ  |  AJE & taj  ; 
 AJF <=  RBF & TAJ  |  RDF & TAJ  |  AJF & taj  ; 
 OAH <= NHH ; 
 OBH <= NGH ; 
 OCH <= NGH ; 
 ODH <= NGH ; 
 NBE <=  JGE  |  JHE  ; 
 ALE <=  RBE & TAL  |  RDE & TAL  |  ALE & tal  ; 
 ALF <=  RBF & TAL  |  RDF & TAL  |  ALF & tal  ; 
 ncn <= nbf ; 
 nef <= ncn ; 
 nhe <= nge ; 
 nhf <= ngf ; 
 NBF <=  JGF  |  JHF  ; 
 ANE <=  RBE & TAN  |  RDE & TAN  |  ANE & tan  ; 
 ANF <=  RBF & TAN  |  RDF & TAN  |  ANF & tan  ; 
 NGC <=  TXA & NAC  |  TXB & NCC  |  TXC & NEC  |  TXD & NFC  ; 
 OAE <= NHE ; 
 OBE <= NGE ; 
 OCE <= NGE ; 
 ODE <= NGE ; 
 APE <=  RBE & TAP  |  RDE & TAP  |  APE & tap  ; 
 APF <=  RBF & TAP  |  RDF & TAP  |  APF & tap  ; 
 qza <= qia ; 
 qzb <= qib ; 
 qzc <= qic ; 
 qzd <= qid ; 
 OAF <= NHF ; 
 OBF <= NGF ; 
 OCF <= NGF ; 
 ODF <= NGF ; 
 CBC <=  JAG  |  JBG  ; 
 CBD <=  JAH  |  JBH  ; 
 KBC <=  gbc & hbc  |  GBC & HBC  ; 
 KBG <=  TBA & hbc  ; 
 KBD <=  gbd & hbd  |  GBD & HBD  ; 
 KBH <=  TBB & hbd  ; 
 KFD <=  gfd & hfd  |  GFD & HFD  ; 
 KFH <=  TBD & hfd  ; 
 KFC <=  gfc & hfc  |  GFC & HFC  ; 
 KFG <=  TBC & hfc  ; 
 CFC <=  JCG  |  JDG  ; 
 CFD <=  JCH  |  JDH  ; 
 nhg <= ngg ; 
 nhh <= ngh ; 
 AAG <=  RAG & TAA  |  RCG & TAA  |  AAG & taa  ; 
 AAH <=  RAH & TAA  |  RCH & TAA  |  AAH & taa  ; 
 TAA <= FAA ; 
 TAB <= FAB ; 
 TAC <= FAC ; 
 TAD <= FAD ; 
 rco <= rdg ; 
 rcp <= rdh ; 
 rdg <= rdo ; 
 rdh <= rdp ; 
 ACG <=  RAG & TAC  |  RCG & TAC  |  ACG & tac  ; 
 ACH <=  RAH & TAC  |  RCH & TAC  |  ACH & tac  ; 
 EAD <= QEA ; 
 EBD <= QEB ; 
 ECD <= QEC ; 
 EDD <= QED ; 
 RAG <=  KBC & pab  |  KBG & PAB  ; 
 RAH <=  KBD & pab  |  KBH & PAB  ; 
 AMG <=  RBG & TAM  |  RDG & TAM  |  AMG & tam  ; 
 AMH <=  RBH & TAM  |  RDH & TAM  |  AMH & tam  ; 
 AEG <=  RAG & TAE  |  RCG & TAE  |  AEG & tae  ; 
 AEH <=  RAH & TAE  |  RCH & TAE  |  AEH & tae  ; 
 TAE <= FAE ; 
 TAF <= FAF ; 
 TAG <= FAG ; 
 TAH <= FAH ; 
 neg <= nco ; 
 neh <= ncp ; 
 rcg <= rco ; 
 rch <= rcp ; 
 AGG <=  RAG & TAG  |  RCG & TAG  |  AGG & tag  ; 
 AGH <=  RAH & TAG  |  RCH & TAG  |  AGH & tag  ; 
 EED <= QEE ; 
 EFD <= QEF ; 
 EGD <= QEG ; 
 EHD <= QEH ; 
 AIG <=  RBG & TAI  |  RDG & TAI  |  AIG & tai  ; 
 AIH <=  RBH & TAI  |  RDH & TAI  |  AIH & tai  ; 
 eid <= qea ; 
 ejd <= qeb ; 
 ekd <= qec ; 
 eld <= qed ; 
 RBG <=  KFC & paf  |  KFG & PAF  ; 
 RBH <=  KFD & paf  |  KFH & PAF  ; 
 AKG <=  RBG & TAK  |  RDG & TAK  |  AKG & tak  ; 
 AKH <=  RBH & TAK  |  RDH & TAK  |  AKH & tak  ; 
 TAI <= FBA ; 
 TAJ <= FBB ; 
 TAK <= FBC ; 
 TAL <= FBD ; 
 emd <= qee ; 
 endd <= qef ; 
 eod <= QEG ; 
 epd <= QEH ; 
 AOG <=  RBG & TAO  |  RDG & TAO  |  AOG & tao  ; 
 AOH <=  RBH & TAO  |  RDH & TAO  |  AOH & tao  ; 
 TAM <= FBE ; 
 TAN <= FBF ; 
 TAO <= FBG ; 
 TAP <= FBH ; 
 ABG <=  RAG & TAB  |  RCG & TAB  |  ABG & tab  ; 
 ABH <=  RAH & TAB  |  RCH & TAB  |  ABH & tab  ; 
 RDO <=  REGG & TCE  |  ICG & TDE  |  IEG & TEA  |  IGG & TFE  ; 
 OKA <= QIA & qza |  ZZO & QZA ; 
 ADG <=  RAG & TAD  |  RCG & TAD  |  ADG & tad  ; 
 ADH <=  RAH & TAD  |  RCH & TAD  |  ADH & tad  ; 
 RDP <=  REH & TCF  |  ICH & TDF  |  IEH & TEB  |  IGH & TFF  ; 
 TJE <= QYB ; 
 TJF <= QYB ; 
 tjg <= qyc ; 
 AFG <=  RAG & TAF  |  RCG & TAF  |  AFG & taf  ; 
 AFH <=  RAH & TAF  |  RCH & TAF  |  AFH & taf  ; 
 NAG <=  JEG  |  JFG  ; 
 AHG <=  RAG & TAH  |  RCG & TAH  |  AHG & tah  ; 
 AHH <=  RAH & TAH  |  RCH & TAH  |  AHH & tah  ; 
 REGG <= IAG ; 
 REH <= IAH ; 
 nco <= nbg ; 
 ncp <= nbh ; 
 NAH <=  JEH  |  JFH  ; 
 AJG <=  RBG & TAJ  |  RDG & TAJ  |  AJG & taj  ; 
 AJH <=  RBH & TAJ  |  RDH & TAJ  |  AJH & taj  ; 
 NBG <=  JGG  |  JHG  ; 
 ALG <=  RBG & TAL  |  RDG & TAL  |  ALG & tal  ; 
 ALH <=  RBH & TAL  |  RDH & TAL  |  ALH & tal  ; 
 NBH <=  JGH  |  JHH  ; 
 ANG <=  RBG & TAN  |  RDG & TAN  |  ANG & tan  ; 
 ANH <=  RBH & TAN  |  RDH & TAN  |  ANH & tan  ; 
 NGD <=  TXA & NAD  |  TXB & NCD  |  TXC & NED  |  TXD & NFD  ; 
 APG <=  RBG & TAP  |  RDG & TAP  |  APG & tap  ; 
 APH <=  RBH & TAP  |  RDH & TAP  |  APH & tap  ; 
 CCA <=  JAI  |  JBI  ; 
 CCB <=  JAJ  |  JBJ  ; 
 KCA <=  HCA & hca  ; 
 KCE <=  TBA & hca  ; 
 TBE <= TJG ; 
 TBF <= TJG ; 
 KCB <=  gcb & hcb  |  GCB & HCB  ; 
 KCF <=  TBB & hcb  ; 
 mac <= gce ; 
 KGB <=  ggb & hgb  |  GGB & HGB  ; 
 KGF <=  TBD & hgb  ; 
 KGA <=  HGA & hga  ; 
 KGE <=  TBC & hga  ; 
 CGA <=  JCI  |  JDI  ; 
 mag <= gge ; 
 CGB <=  JCJ  |  JDJ  ; 
 AAI <=  RAI & TAA  |  RCI & TAA  |  AAI & taa  ; 
 AAJ <=  RAJ & TAA  |  RCJ & TAA  |  AAJ & taa  ; 
 qcq <= qcp ; 
 qfm <= qfl ; 
 ACI <=  RAI & TAC  |  RCE & TAC  |  ACI & tac  ; 
 ACJ <=  RAJ & TAC  |  RCJ & TAC  |  ACJ & tac  ; 
 EAE <= QEA ; 
 EBE <= QEB ; 
 ECE <= QEC ; 
 EDE <= QED ; 
 RAI <=  KCA & pac  |  KCE & PAC  ; 
 RAJ <=  KCB & pac  |  KCF & PAC  ; 
 AMI <=  RBI & TAM  |  RDI & TAM  |  AMI & tam  ; 
 AMJ <=  RBJ & TAM  |  RDJ & TAM  |  AMJ & tam  ; 
 AEI <=  RAI & TAE  |  RCI & TAE  |  AEI & tae  ; 
 AEJ <=  RAJ & TAE  |  RCJ & TAE  |  AEJ & tae  ; 
 TBA <= TJF ; 
 TBB <= TJF ; 
 TBC <= TJF ; 
 TBD <= TJF ; 
 qfg <= qfc ; 
 qfh <= qfg ; 
 qfi <= qfh ; 
 qfj <= qfi ; 
 qcs <= qcr ; 
 qct <= qcs ; 
 qfk <= qfj ; 
 qfl <= qfk ; 
 AGI <=  RAI & TAG  |  RCI & TAG  |  AGI & tag  ; 
 AGJ <=  RAJ & TAG  |  RCJ & TAG  |  AGJ & tag  ; 
 EEE <= QEE ; 
 EFE <= QEF ; 
 EGE <= QEG ; 
 EHE <= QEH ; 
 qcr <= qcq ; 
 qcu <= qcq ; 
 QFN <=  QFM  |  QZE  ; 
 AII <=  RBI & TAI  |  RDI & TAI  |  AII & tai  ; 
 AIJ <=  RBJ & TAI  |  RDJ & TAI  |  AIJ & tai  ; 
 eie <= qea ; 
 eje <= qeb ; 
 eke <= qec ; 
 ele <= qed ; 
 RBI <=  KGA & pag  |  KGE & PAG  ; 
 RBJ <=  KGB & pag  |  KGF & PAG  ; 
 AKI <=  RBI & TAK  |  RDI & TAK  |  AKI & tak  ; 
 AKJ <=  RBJ & TAK  |  RDJ & TAK  |  AKJ & tak  ; 
 QCA <=  TLA  |  TLB  |  TLC  |  TLD  ; 
 qfa <=  qii & qij & qik & qil  ; 
 eme <= qee ; 
 ene <= qef ; 
 eoe <= QEG ; 
 epe <= QEH ; 
 AOI <=  RBI & TAO  |  RDI & TAO  |  AOI & tao  ; 
 AOJ <=  RBJ & TAO  |  RDJ & TAO  |  AOJ & tao  ; 
 ABI <=  RAI & TAB  |  RCI & TAB  |  ABI & tab  ; 
 ABJ <=  RAJ & TAB  |  RCJ & TAB  |  ABJ & tab  ; 
 qea <=  QNC  |  QNB  |  QNA  ; 
 qeb <=  QNC  |  QNB  |  qna  ; 
 ADI <=  RAI & TAD  |  RCI & TAD  |  ADI & tad  ; 
 ADJ <=  RAJ & TAD  |  RCJ & TAD  |  ADJ & tad  ; 
 OKB <= QIB & qzb |  ZZO & QZB ; 
 AFI <=  RAI & TAF  |  RCI & TAF  |  AFI & taf  ; 
 AFJ <=  RAJ & TAF  |  RCJ & TAF  |  AFJ & taf  ; 
 nca <= nai ; 
 qze <= iya ; 
 NAI <=  JEI  |  JFI  ; 
 AHI <=  RAI & TAH  |  RCI & TAH  |  AHI & tah  ; 
 AHJ <=  RAJ & TAH  |  RCJ & TAH  |  AHJ & tah  ; 
 ncb <= naj ; 
 nda <= nbi ; 
 ndb <= nbj ; 
 nei <= nda ; 
 NAJ <=  JEJ  |  JFJ  ; 
 AJI <=  RBI & TAJ  |  RDI & TAJ  |  AJI & taj  ; 
 AJJ <=  RBJ & TAJ  |  RDJ & TAJ  |  AJJ & taj  ; 
 nej <= ndb ; 
 nfa <= nei ; 
 nfb <= nej ; 
 NBI <=  JGI  |  JHI  ; 
 ALI <=  RBI & TAL  |  RDI & TAL  |  ALI & tal  ; 
 ALJ <=  RBJ & TAL  |  RDJ & TAL  |  ALJ & tal  ; 
 NBJ <=  JGJ  |  JHJ  ; 
 ANI <=  RBI & TAN  |  RDI & TAN  |  ANI & tan  ; 
 ANJ <=  RBJ & TAN  |  RDJ & TAN  |  ANJ & tan  ; 
 NGE <=  TXE & NAE  |  TXF & NCE  |  TXG & NEE  |  TXH & NFE  ; 
 QIB <=  QQB & qhi & IJA  |  QIB & twe  ; 
 QIF <=  QQB & qhi & IJA  |  QIB & twe  ; 
 QIJ <=  QQB & qhi & IJA  |  QIB & twe  ; 
 API <=  RBI & TAP  |  RDI & TAP  |  API & tap  ; 
 APJ <=  RBJ & TAP  |  RDJ & TAP  |  APJ & tap  ; 
 QIC <=  QQC & qhg & IKA  |  QIC & twe  ; 
 QIG <=  QQC & qhg & IKA  |  QIC & twe  ; 
 QIK <=  QQC & qhg & IKA  |  QIC & twe  ; 
 CCC <=  JAK  |  JBK  ; 
 CCD <=  JAL  |  JBL  ; 
 KCC <=  gcc & hcc  |  GCC & HCC  ; 
 KCG <=  TBA & hcc  ; 
 KCD <=  gcd & hcd  |  GCD & HCD  ; 
 KCH <=  TBB & hcd  ; 
 KGD <=  ggd & hgd  |  GGD & HGD  ; 
 KGH <=  TBD & hgd  ; 
 KGC <=  ggc & hgc  |  GGC & HGC  ; 
 KGG <=  TBC & hgc  ; 
 CGC <=  JCK  |  JDK  ; 
 CGD <=  JCL  |  JDL  ; 
 AAK <=  RAK & TAA  |  RCK & TAA  |  AAK & taa  ; 
 AAL <=  RAL & TAA  |  RCL & TAA  |  AAL & taa  ; 
 ACK <=  RAK & TAC  |  RCK & TAC  |  ACK & tac  ; 
 ACL <=  RAL & TAC  |  RCL & TAC  |  ACL & tac  ; 
 EAF <= QEA ; 
 EBF <= QEB ; 
 ECF <= QEC ; 
 EDF <= QED ; 
 RAK <=  KCC & pac  |  KCG & PAC  ; 
 RAL <=  KCD & pac  |  KCH & PAC  ; 
 AMK <=  RBK & TAM  |  RDK & TAM  |  AMK & tam  ; 
 AML <=  RBL & TAM  |  RDL & TAM  |  AML & tam  ; 
 AEK <=  RAK & TAE  |  RCK & TAE  |  AEK & tae  ; 
 AEL <=  RAL & TAE  |  RCL & TAE  |  AEL & tae  ; 
 AGK <=  RAK & TAG  |  RCK & TAG  |  AGK & tag  ; 
 AGL <=  RAL & TAG  |  RCL & TAG  |  AGL & tag  ; 
 EEF <= QEE ; 
 EFF <= QEF ; 
 EGF <= QEG ; 
 EHF <= QEH ; 
 qcp <= qcg ; 
 QCC <=  QUA & QUD  ; 
 QCD <=  QVA & QUD  ; 
 AIK <=  RBK & TAI  |  RDK & TAI  |  AIK & tai  ; 
 AIL <=  RBL & TAI  |  RDL & TAI  |  AIL & tai  ; 
 eif <= qea ; 
 ejf <= qeb ; 
 ekf <= qec ; 
 elf <= qed ; 
 RBK <=  KGC & pag  |  KGG & PAG  ; 
 RBL <=  KGD & pag  |  KGH & PAG  ; 
 AKK <=  RBK & TAK  |  RDK & TAK  |  AKK & tak  ; 
 AKL <=  RBL & TAK  |  RDL & TAK  |  AKL & tak  ; 
 QFC <= qfb & QFA ; 
 QCG <=  QCC  |  QCD  |  QCE  |  QCF  ; 
 emf <= qee ; 
 enf <= qef ; 
 eof <= QEG ; 
 epf <= QEH ; 
 AOK <=  RBK & TAO  |  RDK & TAO  |  AOK & tao  ; 
 AOL <=  RBL & TAO  |  RDL & TAO  |  AOL & tao  ; 
 qch <= qca ; 
 qfb <= qfa ; 
 ABK <=  RAK & TAB  |  RCK & TAB  |  ABK & tab  ; 
 ABL <=  RAL & TAB  |  RCL & TAB  |  ABL & tab  ; 
 qec <=  QNC  |  qnb  |  QNA  ; 
 qed <=  QNC  |  qnb  |  qna  ; 
 ADK <=  RAK & TAD  |  RCK & TAD  |  ADK & tad  ; 
 ADL <=  RAL & TAD  |  RCL & TAD  |  ADL & tad  ; 
 AFK <=  RAK & TAF  |  RCK & TAF  |  AFK & taf  ; 
 AFL <=  RAL & TAF  |  RCL & TAF  |  AFL & taf  ; 
 OKC <= QIC & qzc |  ZZO & QZC ; 
 NAK <=  JEK  |  JFK  ; 
 AHK <=  RAK & TAH  |  RCK & TAH  |  AHK & tah  ; 
 AHL <=  RAL & TAH  |  RCL & TAH  |  AHL & tah  ; 
 ncc <= nak ; 
 ncd <= nal ; 
 ndc <= nbk ; 
 ndd <= nbl ; 
 NAL <=  JEL  |  JFL  ; 
 AJK <=  RBK & TAJ  |  RDK & TAJ  |  AJK & taj  ; 
 AJL <=  RBL & TAJ  |  RDL & TAJ  |  AJL & taj  ; 
 OKD <= QID & qzd |  ZZO & QZD ; 
 NBK <=  JGK  |  JHK  ; 
 ALK <=  RBK & TAL  |  RDK & TAL  |  ALK & tal  ; 
 ALL <=  RBL & TAL  |  RDL & TAL  |  ALL & tal  ; 
 nek <= ndc ; 
 nel <= ndd ; 
 nfc <= nek ; 
 nfd <= nel ; 
 NBL <=  JGL  |  JHL  ; 
 ANK <=  RBK & TAN  |  RDK & TAN  |  ANK & tan  ; 
 ANL <=  RBL & TAN  |  RDL & TAN  |  ANL & tan  ; 
 NGF <=  TXE & NAF  |  TXF & NCF  |  TXG & NEF  |  TXH & NFF  ; 
 QID <=  QQD & qhg & ILA  |  QID & twe  ; 
 QIH <=  QQD & qhg & ILA  |  QID & twe  ; 
 QIL <=  QQD & qhg & ILA  |  QID & twe  ; 
 APK <=  RBK & TAP  |  RDK & TAP  |  APK & tap  ; 
 APL <=  RBL & TAP  |  RDL & TAP  |  APL & tap  ; 
 twe <= qfn ; 
 CDA <=  JAM  |  JBM  ; 
 CDE <=  JAM  |  JBM  ; 
 CDB <=  JAN  |  JBN  ; 
 KDA <=  HDA & hda  ; 
 KDE <=  TBA & hda  ; 
 KDB <=  gdb & hdb  |  GDB & HDB  ; 
 KDF <=  TBB & hdb  ; 
 KHB <=  ghb & hhb  |  GHB & HHB  ; 
 KHF <=  TBD & hhb  ; 
 QAF <=  GAE & GBE & GCE & GDE  ; 
 KHA <=  HHA & hha  ; 
 KHE <=  TBC & hha  ; 
 CHA <=  JCM  |  JDM  ; 
 CHB <=  JCN  |  JDN  ; 
 AAM <=  RAM & TAA  |  RCM & TAA  |  AAM & taa  ; 
 AAN <=  RAN & TAA  |  RCN & TAA  |  AAN & taa  ; 
 ACM <=  RAM & TAC  |  RCM & TAC  |  ACM & tac  ; 
 ACN <=  RAN & TAC  |  RCN & TAC  |  ACN & tac  ; 
 EAG <= QEA ; 
 EBG <= QEB ; 
 ECG <= QEC ; 
 EDG <= QED ; 
 RAM <=  KDA & pad  |  KDE & PAD  ; 
 RAN <=  KDB & pad  |  KDF & PAD  ; 
 AMM <=  RBM & TAM  |  RDM & TAM  |  AMM & tam  ; 
 AMN <=  RBN & TAM  |  RDN & TAM  |  AMN & tam  ; 
 AEM <=  RAM & TAE  |  RCM & TAE  |  AEM & tae  ; 
 AEN <=  RAN & TAE  |  RCN & TAE  |  AEN & tae  ; 
 AGM <=  RAM & TAG  |  RCM & TAG  |  AGM & tag  ; 
 AGN <=  RAN & TAG  |  RCN & TAG  |  AGN & tag  ; 
 EEG <= QEE ; 
 EFG <= QEF ; 
 EGG <= QEG ; 
 EHG <= QEH ; 
 AIM <=  RBM & TAI  |  RDM & TAI  |  AIM & tai  ; 
 AIN <=  RBN & TAI  |  RDN & TAI  |  AIN & tai  ; 
 eig <= qea ; 
 ejg <= qeb ; 
 ekg <= qec ; 
 elg <= qed ; 
 RBM <=  KHA & pah  |  KHE & PAH  ; 
 RBN <=  KHB & pah  |  KHF & PAH  ; 
 AKM <=  RBM & TAK  |  RDM & TAK  |  AKM & tak  ; 
 AKN <=  RBN & TAK  |  RDN & TAK  |  AKN & tak  ; 
 TLN <=  TLN & qcn  |  TLF  ; 
 TLO <=  TLO & qcn  |  TLG  ; 
 emg <= qee ; 
 eng <= qef ; 
 eog <= QEG ; 
 epg <= QEH ; 
 AON <=  RBN & TAO  |  RDN & TAO  |  AON & tao  ; 
 AOM <=  RBM & TAO  |  RDM & TAO  |  AOM & tao  ; 
 QCE <=  QWA & QWC  ; 
 QCF <=  QXA & QWC  ; 
 ABM <=  RAM & TAB  |  RCM & TAB  |  ABM & tab  ; 
 ABN <=  RAN & TAB  |  RCN & TAB  |  ABN & tab  ; 
 TLB <= QVD & qve |  ZZO & QVE ; 
 qee <=  qnc  |  QNB  |  QNA  ; 
 qef <=  qnc  |  QNB  |  qna  ; 
 ADM <=  RAM & TAD  |  RCM & TAD  |  ADM & tad  ; 
 ADN <=  RAN & TAD  |  RCN & TAD  |  ADN & tad  ; 
 tlf <= tlb ; 
 AFM <=  RAM & TAF  |  RCM & TAF  |  AFM & taf  ; 
 AFN <=  RAN & TAF  |  RCM & TAF  |  AFN & taf  ; 
 TJB <= QIJ ; 
 TKB <= QIJ ; 
 NAM <=  JEM  |  JFM  ; 
 AHM <=  RAM & TAH  |  RCM & TAH  |  AHM & tah  ; 
 AHN <=  RAN & TAH  |  RCN & TAH  |  AHN & tah  ; 
 nce <= nam ; 
 ncf <= nan ; 
 nde <= nbm ; 
 ndf <= nbn ; 
 NAN <=  JEN  |  JFN  ; 
 AJM <=  RBM & TAJ  |  RDM & TAJ  |  AJM & taj  ; 
 AJN <=  RBN & TAJ  |  RDN & TAJ  |  AJN & taj  ; 
 NBM <=  JGM  |  JHM  ; 
 ALM <=  RBM & TAL  |  RDM & TAL  |  ALM & tal  ; 
 ALN <=  RBN & TAL  |  RDN & TAL  |  ALN & tal  ; 
 nem <= nde ; 
 nen <= ndf ; 
 nfe <= nem ; 
 nff <= nen ; 
 NBN <=  JGN  |  JHN  ; 
 ANM <=  RBM & TAN  |  RDM & TAN  |  ANM & tan  ; 
 ANN <=  RBN & TAN  |  RDN & TAN  |  ANN & tan  ; 
 NGG <=  TXE & NAG  |  TXF & NCG  |  TXG & NEG  |  TXH & NFG  ; 
 qci <= qch ; 
 qcj <= qci ; 
 qcn <= qcj ; 
 APM <=  RBM & TAP  |  RDM & TAP  |  APM & tap  ; 
 APN <=  RBN & TAP  |  RDN & TAP  |  APN & tap  ; 
 QCL <=  QCJ  |  TPA  ; 
 QCM <=  QCJ  |  TPA  ; 
 CDC <=  JAO  |  JBO  ; 
 CDD <=  JAP  |  JBP  ; 
 KDC <=  gdc & hdc  |  GDC & HDC  ; 
 KDG <=  TBA & hdc  ; 
 KDD <=  gdd & hdd  |  GDD & HDD  ; 
 KDH <=  TBB & hdd  ; 
 CHC <=  JCO  |  JDO  ; 
 KHD <=  ghd & hhd  |  GHD & HHD  ; 
 KHH <=  TBD & hhd  ; 
 KHC <=  ghc & hhc  |  GHC & HHC  ; 
 KHG <=  TBC & hhc  ; 
 CHD <=  JCP  |  JDP  ; 
 QYD <= QYC ; 
 AAO <=  RAO & TAA  |  RCO & TAA  |  AAO & taa  ; 
 AAP <=  RAP & TAA  |  RCP & TAA  |  AAP & taa  ; 
 QYB <=  QYA & QYE  ; 
 QYC <=  QYB & QYE  ; 
 QYE <=  QUA & QUC  |  QVA & QVC  |  QWA & QWC  |  QXA & QXC  ; 
 ACO <=  RAO & TAC  |  RCO & TAC  |  ACO & tac  ; 
 ACP <=  RAP & TAC  |  RCP & TAC  |  ACP & tac  ; 
 EAH <= QEA ; 
 EBH <= QEB ; 
 ECH <= QEC ; 
 EDH <= QED ; 
 RAO <=  KDC & pad  |  KDG & PAD  ; 
 RAP <=  KDD & pad  |  KDH & PAD  ; 
 AMO <=  RBO & TAM  |  RDO & TAM  |  AMO & tam  ; 
 AMP <=  RBP & TAM  |  RDP & TAM  |  AMP & tam  ; 
 AEO <=  RAO & TAE  |  RCO & TAE  |  AEO & tae  ; 
 TLC <= QWA & qwc |  ZZO & QWC ; 
 QYA <=  QUA & QUB  |  QVA & QVB  |  QWA & QWB  |  QXA & QXB  ; 
 AGO <=  RAO & TAG  |  RCO & TAG  |  AGO & tag  ; 
 AGP <=  RAP & TAG  |  RCP & TAG  |  AGP & tag  ; 
 EEH <= QEE ; 
 EFH <= QEF ; 
 EGH <= QEG ; 
 EHH <= QEH ; 
 AIO <=  RBO & TAI  |  RDO & TAI  |  AIO & tai  ; 
 AIP <=  RBP & TAI  |  RDP & TAI  |  AIP & tai  ; 
 eih <= qea ; 
 ejh <= qeb ; 
 ekh <= qec ; 
 elh <= qed ; 
 RBO <=  KHC & pah  |  KHG & PAH  ; 
 RBP <=  KHD & pah  |  KHH & PAH  ; 
 AKO <=  RBO & TAK  |  RDO & TAK  |  AKO & tak  ; 
 AKP <=  RBP & TAK  |  RDP & TAK  |  AKP & tak  ; 
 AEP <=  RAP & TAE  |  RCP & TAE  |  AEP & tae  ; 
 TLP <=  TLP & TAE  |  TLH & TAE  ; 
 emh <= qee ; 
 enh <= qef ; 
 eoh <= QEG ; 
 eph <= QEH ; 
 AOO <=  RBO & TAO  |  RDO & TAO  |  AOO & tao  ; 
 AOP <=  RBP & TAO  |  RDP & TAO  |  AOP & tao  ; 
 TLD <= QXA & qxc |  ZZO & QXC ; 
 ABO <=  RAO & TAB  |  RCO & TAB  |  ABO & tab  ; 
 ABP <=  RAP & TAB  |  RCP & TAB  |  ABP & tab  ; 
 tlg <= tlc ; 
 qeg <=  qnc  |  qnb  |  QNA  ; 
 qeh <=  qnc  |  qnb  |  qna  ; 
 ADO <=  RAO & TAD  |  RCO & TAD  |  ADO & tad  ; 
 ADP <=  RAP & TAD  |  RCP & TAD  |  ADP & tad  ; 
 QVE <= IVB ; 
 QWA <= IWA ; 
 QWB <= IWB ; 
 QWC <= IWC ; 
 QVA <= IVA ; 
 QVB <= IVB ; 
 QVC <= IVC ; 
 QVD <= IVA ; 
 AFO <=  RAO & TAF  |  RCO & TAF  |  AFO & taf  ; 
 AFP <=  RAP & TAF  |  RCP & TAF  |  AFP & taf  ; 
 TJC <= QIK ; 
 TKC <= QIK ; 
 NAO <=  JEO  |  JFO  ; 
 AHO <=  RAO & TAH  |  RCO & TAH  |  AHO & tah  ; 
 AHP <=  RAP & TAH  |  RCP & TAH  |  AHP & tah  ; 
 ncg <= nao ; 
 nch <= nap ; 
 ndg <= nbo ; 
 ndh <= nbp ; 
 NAP <=  JEP  |  JFP  ; 
 AJO <=  RBO & TAJ  |  RDO & TAJ  |  AJO & taj  ; 
 AJP <=  RBP & TAJ  |  RDP & TAJ  |  AJP & taj  ; 
 neo <= ndg ; 
 nep <= ndh ; 
 nfg <= neo ; 
 nfh <= nep ; 
 NBO <=  JGO  |  JHO  ; 
 ALO <=  RBO & TAL  |  RDO & TAL  |  ALO & tal  ; 
 ALP <=  RBP & TAL  |  RDP & TAL  |  ALP & tal  ; 
 TJD <= QIL ; 
 TKD <= QIL ; 
 NBP <=  JGP  |  JHP  ; 
 ANO <=  RBO & TAN  |  RDO & TAN  |  ANO & tan  ; 
 ANP <=  RBP & TAN  |  RDP & TAN  |  ANP & tan  ; 
 NGH <=  TXE & NAH  |  TXF & NCH  |  TXG & NEH  |  TXH & NFH  ; 
 QQA <= ipa ; 
 QXA <= IXA ; 
 QXB <= IXB ; 
 QXC <= IXC ; 
 APO <=  RBO & TAP  |  RDO & TAP  |  APO & tap  ; 
 APP <=  RBP & TAP  |  RDP & TAP  |  APP & tap  ; 
 tlh <= tld ; 
 qqb <= qqa ; 
 qqc <= qqb ; 
 qqd <= qqc ; 
 end 
endmodule;
