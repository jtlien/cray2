module mc( IZZ,
 IAL, 
 IAM, 
 IAN, 
 IAO, 
 IAP, 
 IBA, 
 IBB, 
 IBC, 
 IBD, 
 IBE, 
 IBF, 
 IBG, 
 IBH, 
 IBI, 
 IBJ, 
 IBK, 
 IBL, 
 IBM, 
 IBN, 
 IBO, 
 IBP, 
 ICA, 
 ICB, 
 ICC, 
 ICD, 
 ICE, 
 ICF, 
 ICG, 
 ICH, 
 ICI, 
 ICJ, 
 ICK, 
 ICL, 
 ICM, 
 ICN, 
 ICO, 
 ICP, 
 IDL, 
 IDM, 
 IDN, 
 IDO, 
 IDP, 
 IEA, 
 IEB, 
 IEC, 
 IED, 
 IEE, 
 IEF, 
 IEG, 
 IEH, 
 IEI, 
 IEJ, 
 IEK, 
 IEL, 
 IEM, 
 IEN, 
 IEO, 
 IEP, 
 IFA, 
 IFB, 
 IFC, 
 IFD, 
 IFE, 
 IFFF , 
 IFG, 
 IFH, 
 IFI, 
 IFJ, 
 IFK, 
 IFL, 
 IFM, 
 IFN, 
 IFO, 
 IFP, 
 IGA, 
 IGB, 
 IGC, 
 IGD, 
 IGE, 
 IGF, 
 IGG, 
 IGH, 
 IGI, 
 IGJ, 
 ILA, 
 ILB, 
 ILC, 
 ILD, 
 ILE, 
 ILF, 
 ILG, 
 ILH, 
 ILI, 
 ILJ, 
 ILK, 
 ILL, 
 ILM, 
 IMA, 
 IMB, 
 IMC, 
 IMD, 
 IME, 
 IMF, 
 IMG, 
 IMH, 
 IMI, 
 IMJ, 
 IMK, 
 IML, 
 INA, 
 INB, 
 INC, 
 IND, 
 INE, 
 INF, 
 IOA, 
 IOB, 
 IQC, 
 IQD, 
 IQE, 
 IQF, 
 IQG, 
 IQH, 
 IRA, 
 IRB, 
 IRC, 
 OGA, 
 OGB, 
 OGC, 
 OGD, 
 OGE, 
 OGF, 
 OGG, 
 OGH, 
 OGI, 
 OHA, 
 OHB, 
 OHC, 
 OHD, 
 OHE, 
 OHF, 
 OIE, 
 OIF, 
 OKA, 
 OKB, 
 OKC, 
 OLC, 
 OMA, 
 OMB, 
 OPA, 
 OPB, 
 OPC, 
 OPD, 
 OPE, 
 OPF, 
 OPG, 
 OPI, 
 OPK, 
 OPM, 
 OPO, 
 OPQ, 
 OPS, 
 OPU, 
 OQA, 
 OQC, 
 OQG, 
 OQI, 
 OQK, 
 OQM, 
 OQO, 
 OQQ, 
 OQS, 
OQU ); 
    
 input IZZ; 
 input IAL; 
 input IAM; 
 input IAN; 
 input IAO; 
 input IAP; 
 input IBA; 
 input IBB; 
 input IBC; 
 input IBD; 
 input IBE; 
 input IBF; 
 input IBG; 
 input IBH; 
 input IBI; 
 input IBJ; 
 input IBK; 
 input IBL; 
 input IBM; 
 input IBN; 
 input IBO; 
 input IBP; 
 input ICA; 
 input ICB; 
 input ICC; 
 input ICD; 
 input ICE; 
 input ICF; 
 input ICG; 
 input ICH; 
 input ICI; 
 input ICJ; 
 input ICK; 
 input ICL; 
 input ICM; 
 input ICN; 
 input ICO; 
 input ICP; 
 input IDL; 
 input IDM; 
 input IDN; 
 input IDO; 
 input IDP; 
 input IEA; 
 input IEB; 
 input IEC; 
 input IED; 
 input IEE; 
 input IEF; 
 input IEG; 
 input IEH; 
 input IEI; 
 input IEJ; 
 input IEK; 
 input IEL; 
 input IEM; 
 input IEN; 
 input IEO; 
 input IEP; 
 input IFA; 
 input IFB; 
 input IFC; 
 input IFD; 
 input IFE; 
 input IFFF ; 
 input IFG; 
 input IFH; 
 input IFI; 
 input IFJ; 
 input IFK; 
 input IFL; 
 input IFM; 
 input IFN; 
 input IFO; 
 input IFP; 
 input IGA; 
 input IGB; 
 input IGC; 
 input IGD; 
 input IGE; 
 input IGF; 
 input IGG; 
 input IGH; 
 input IGI; 
 input IGJ; 
 input ILA; 
 input ILB; 
 input ILC; 
 input ILD; 
 input ILE; 
 input ILF; 
 input ILG; 
 input ILH; 
 input ILI; 
 input ILJ; 
 input ILK; 
 input ILL; 
 input ILM; 
 input IMA; 
 input IMB; 
 input IMC; 
 input IMD; 
 input IME; 
 input IMF; 
 input IMG; 
 input IMH; 
 input IMI; 
 input IMJ; 
 input IMK; 
 input IML; 
 input INA; 
 input INB; 
 input INC; 
 input IND; 
 input INE; 
 input INF; 
 input IOA; 
 input IOB; 
 input IQC; 
 input IQD; 
 input IQE; 
 input IQF; 
 input IQG; 
 input IQH; 
 input IRA; 
 input IRB; 
 input IRC; 
 output OGA; 
 output OGB; 
 output OGC; 
 output OGD; 
 output OGE; 
 output OGF; 
 output OGG; 
 output OGH; 
 output OGI; 
 output OHA; 
 output OHB; 
 output OHC; 
 output OHD; 
 output OHE; 
 output OHF; 
 output OIE; 
 output OIF; 
 output OKA; 
 output OKB; 
 output OKC; 
 output OLC; 
 output OMA; 
 output OMB; 
 output OPA; 
 output OPB; 
 output OPC; 
 output OPD; 
 output OPE; 
 output OPF; 
 output OPG; 
 output OPI; 
 output OPK; 
 output OPM; 
 output OPO; 
 output OPQ; 
 output OPS; 
 output OPU; 
 output OQA; 
 output OQC; 
 output OQG; 
 output OQI; 
 output OQK; 
 output OQM; 
 output OQO; 
 output OQQ; 
 output OQS; 
 output OQU; 
  
  
reg  CAL ;
reg  CAM ;
reg  CAN ;
reg  CAO ;
reg  CAP ;
reg  CBA ;
reg  CBB ;
reg  CBC ;
reg  CBD ;
reg  CBE ;
reg  CBF ;
reg  CBG ;
reg  CBH ;
reg  CBI ;
reg  CBJ ;
reg  CBK ;
reg  CBL ;
reg  CBM ;
reg  CBN ;
reg  CBO ;
reg  CBP ;
reg  CCA ;
reg  CCB ;
reg  CCC ;
reg  CCD ;
reg  CCE ;
reg  CCF ;
reg  CCG ;
reg  CCH ;
reg  CCI ;
reg  CCJ ;
reg  CCK ;
reg  CCL ;
reg  CCM ;
reg  CCN ;
reg  CCO ;
reg  CCP ;
reg  CDP ;
reg  CEA ;
reg  CEB ;
reg  CEC ;
reg  CED ;
reg  CEE ;
reg  CEF ;
reg  CEG ;
reg  CEH ;
reg  CEI ;
reg  CEJ ;
reg  CEK ;
reg  CEL ;
reg  CEM ;
reg  CEN ;
reg  CEO ;
reg  CEP ;
reg  CFA ;
reg  CFB ;
reg  CFC ;
reg  CFD ;
reg  CFE ;
reg  CFF ;
reg  CFG ;
reg  CFH ;
reg  CFI ;
reg  CFJ ;
reg  CFK ;
reg  CFL ;
reg  CFM ;
reg  CFN ;
reg  CFO ;
reg  CFP ;
reg  cgn ;
reg  cgo ;
reg  cgp ;
reg  cha ;
reg  chb ;
reg  chc ;
reg  chd ;
reg  che ;
reg  chf ;
reg  chg ;
reg  chh ;
reg  chi ;
reg  chj ;
reg  chk ;
reg  chl ;
reg  chm ;
reg  chn ;
reg  cho ;
reg  chp ;
reg  cia ;
reg  cib ;
reg  cic ;
reg  cid ;
reg  cie ;
reg  cif ;
reg  cig ;
reg  cih ;
reg  cii ;
reg  cij ;
reg  cik ;
reg  cil ;
reg  cim ;
reg  cin ;
reg  cio ;
reg  cip ;
reg  cki ;
reg  ckj ;
reg  ckk ;
reg  ckl ;
reg  ckm ;
reg  ckn ;
reg  cko ;
reg  ckp ;
reg  cla ;
reg  clb ;
reg  clc ;
reg  cld ;
reg  DAL ;
reg  DAM ;
reg  DAN ;
reg  DAO ;
reg  DAP ;
reg  DBA ;
reg  DBB ;
reg  DBC ;
reg  DBD ;
reg  DBE ;
reg  DBF ;
reg  DBG ;
reg  DBH ;
reg  DBI ;
reg  DBJ ;
reg  DBK ;
reg  DBL ;
reg  DBM ;
reg  DBN ;
reg  DBO ;
reg  DBP ;
reg  DCA ;
reg  DCB ;
reg  DCC ;
reg  DCD ;
reg  DCE ;
reg  DCF ;
reg  DCG ;
reg  DCH ;
reg  DCI ;
reg  DCJ ;
reg  DCK ;
reg  DCL ;
reg  DCM ;
reg  DCN ;
reg  DCO ;
reg  DCP ;
reg  DDO ;
reg  DDP ;
reg  DEA ;
reg  DEB ;
reg  DEC ;
reg  DED ;
reg  DEE ;
reg  DEF ;
reg  DEG ;
reg  DEH ;
reg  DEI ;
reg  DEJ ;
reg  DEK ;
reg  DEL ;
reg  DEM ;
reg  DEN ;
reg  DEO ;
reg  DEP ;
reg  DFA ;
reg  DFB ;
reg  DFC ;
reg  DFD ;
reg  DFE ;
reg  DFF ;
reg  DFG ;
reg  DFH ;
reg  DFI ;
reg  DFJ ;
reg  DFK ;
reg  DFL ;
reg  DFM ;
reg  DFN ;
reg  DFO ;
reg  DFP ;
reg  dha ;
reg  dhb ;
reg  dhc ;
reg  dhd ;
reg  dhe ;
reg  dhf ;
reg  dhg ;
reg  dhh ;
reg  dhi ;
reg  dhj ;
reg  dhk ;
reg  dhl ;
reg  dhm ;
reg  dhn ;
reg  dho ;
reg  dhp ;
reg  dia ;
reg  dib ;
reg  dic ;
reg  did ;
reg  die ;
reg  dif ;
reg  dig ;
reg  dih ;
reg  dii ;
reg  dij ;
reg  dik ;
reg  dil ;
reg  dim ;
reg  din ;
reg  dio ;
reg  dip ;
reg  FAA ;
reg  FAB ;
reg  FAC ;
reg  FAD ;
reg  FAE ;
reg  FAF ;
reg  FAG ;
reg  FAH ;
reg  FAI ;
reg  FAJ ;
reg  FAK ;
reg  FAL ;
reg  FAM ;
reg  FAN ;
reg  fba ;
reg  fbb ;
reg  fbc ;
reg  fbd ;
reg  fbe ;
reg  fbf ;
reg  fbg ;
reg  fbh ;
reg  fbi ;
reg  fbj ;
reg  fbk ;
reg  fbl ;
reg  FCA ;
reg  FCB ;
reg  FCC ;
reg  FCD ;
reg  FCE ;
reg  FCF ;
reg  FCG ;
reg  FCH ;
reg  FCI ;
reg  FCJ ;
reg  FCK ;
reg  FCL ;
reg  FCM ;
reg  fda ;
reg  fdb ;
reg  fdc ;
reg  fdd ;
reg  fde ;
reg  fdf ;
reg  fdg ;
reg  fdh ;
reg  fdi ;
reg  fdj ;
reg  fdk ;
reg  fdl ;
reg  FEA ;
reg  FEB ;
reg  FEC ;
reg  FED ;
reg  FEE ;
reg  FEF ;
reg  FEG ;
reg  FEH ;
reg  FEI ;
reg  FEJ ;
reg  FEK ;
reg  FEL ;
reg  ffa ;
reg  ffb ;
reg  ffc ;
reg  ffd ;
reg  ffe ;
reg  fff ;
reg  ffg ;
reg  ffh ;
reg  ffi ;
reg  ffj ;
reg  ffk ;
reg  ffl ;
reg  FGA ;
reg  FGB ;
reg  FGC ;
reg  FGD ;
reg  FGE ;
reg  FGF ;
reg  FGG ;
reg  FGH ;
reg  FGI ;
reg  FGJ ;
reg  FGK ;
reg  FGL ;
reg  FGM ;
reg  fha ;
reg  fhb ;
reg  fhc ;
reg  fhd ;
reg  fhe ;
reg  fhf ;
reg  fhg ;
reg  fhh ;
reg  fhi ;
reg  fhj ;
reg  fhk ;
reg  FIA ;
reg  FIB ;
reg  FIC ;
reg  FID ;
reg  FIE ;
reg  FIF ;
reg  FIG ;
reg  FIH ;
reg  FII ;
reg  FIJ ;
reg  FIK ;
reg  FIL ;
reg  fja ;
reg  fjb ;
reg  fjc ;
reg  fjd ;
reg  fje ;
reg  fjf ;
reg  fjg ;
reg  fjh ;
reg  fji ;
reg  fjj ;
reg  fjk ;
reg  FKA ;
reg  FKB ;
reg  FKC ;
reg  FKD ;
reg  FKE ;
reg  FKF ;
reg  FKG ;
reg  FKH ;
reg  FKI ;
reg  FKJ ;
reg  FKK ;
reg  fla ;
reg  flb ;
reg  flc ;
reg  fld ;
reg  fle ;
reg  flf ;
reg  flg ;
reg  flh ;
reg  fli ;
reg  flj ;
reg  flk ;
reg  FMA ;
reg  FMB ;
reg  FMC ;
reg  FMD ;
reg  FME ;
reg  FMF ;
reg  FMG ;
reg  FMH ;
reg  FMI ;
reg  FMJ ;
reg  FMK ;
reg  FML ;
reg  fna ;
reg  fnb ;
reg  fnc ;
reg  fnd ;
reg  fne ;
reg  fnf ;
reg  fng ;
reg  fnh ;
reg  fni ;
reg  fnj ;
reg  FOA ;
reg  FOB ;
reg  FOC ;
reg  FOD ;
reg  FOE ;
reg  FOF ;
reg  FOG ;
reg  FOH ;
reg  FOI ;
reg  FOJ ;
reg  FOK ;
reg  fpa ;
reg  fpb ;
reg  fpc ;
reg  fpd ;
reg  fpe ;
reg  fpf ;
reg  fpg ;
reg  fph ;
reg  fpi ;
reg  fpj ;
reg  FQA ;
reg  FQB ;
reg  FQC ;
reg  FQD ;
reg  FQE ;
reg  FQF ;
reg  FQG ;
reg  FQH ;
reg  FQI ;
reg  FQJ ;
reg  fra ;
reg  frb ;
reg  frc ;
reg  frd ;
reg  fre ;
reg  frf ;
reg  frg ;
reg  frh ;
reg  fri ;
reg  frj ;
reg  FSA ;
reg  FSB ;
reg  FSC ;
reg  FSD ;
reg  FSE ;
reg  FSF ;
reg  FSG ;
reg  FSH ;
reg  FSI ;
reg  FSJ ;
reg  FSK ;
reg  fta ;
reg  ftb ;
reg  ftc ;
reg  ftd ;
reg  fte ;
reg  ftf ;
reg  ftg ;
reg  fth ;
reg  fti ;
reg  FUA ;
reg  FUB ;
reg  FUC ;
reg  FUD ;
reg  FUE ;
reg  FUF ;
reg  FUG ;
reg  FUH ;
reg  FUI ;
reg  FUJ ;
reg  HAA ;
reg  HAB ;
reg  HAC ;
reg  HAD ;
reg  HAE ;
reg  HAF ;
reg  HAG ;
reg  hba ;
reg  hbb ;
reg  hbc ;
reg  hbd ;
reg  hbe ;
reg  hbf ;
reg  HCA ;
reg  HCB ;
reg  HCC ;
reg  HCD ;
reg  HCE ;
reg  hda ;
reg  hdb ;
reg  hdc ;
reg  hdd ;
reg  HEA ;
reg  HEB ;
reg  HEC ;
reg  HED ;
reg  HEE ;
reg  HEF ;
reg  hfa ;
reg  hfb ;
reg  hfc ;
reg  hfd ;
reg  hfe ;
reg  HGA ;
reg  HGB ;
reg  HGC ;
reg  HGD ;
reg  HGE ;
reg  HGF ;
reg  HGG ;
reg  hha ;
reg  hhb ;
reg  hhc ;
reg  hhd ;
reg  hhe ;
reg  HIA ;
reg  HIB ;
reg  HIC ;
reg  HID ;
reg  HIE ;
reg  HIF ;
reg  HIG ;
reg  hja ;
reg  hjb ;
reg  hjc ;
reg  hjd ;
reg  hje ;
reg  HKA ;
reg  HKB ;
reg  HKC ;
reg  HKD ;
reg  HKE ;
reg  hla ;
reg  hlb ;
reg  hlc ;
reg  hld ;
reg  hle ;
reg  HMA ;
reg  HMB ;
reg  HMC ;
reg  HMD ;
reg  HME ;
reg  HMF ;
reg  hna ;
reg  hnb ;
reg  hnc ;
reg  hnd ;
reg  hne ;
reg  HOA ;
reg  HOB ;
reg  HOC ;
reg  HOD ;
reg  HOE ;
reg  HOF ;
reg  hpa ;
reg  hpb ;
reg  hpc ;
reg  hpd ;
reg  HQA ;
reg  HQB ;
reg  HQC ;
reg  HQD ;
reg  HQE ;
reg  hra ;
reg  hrb ;
reg  hrc ;
reg  hrd ;
reg  hre ;
reg  HSA ;
reg  HSB ;
reg  HSC ;
reg  HSD ;
reg  HSE ;
reg  hta ;
reg  htb ;
reg  htc ;
reg  htd ;
reg  HUA ;
reg  HUB ;
reg  HUC ;
reg  HUD ;
reg  HUE ;
reg  HUF ;
reg  KAA ;
reg  KAB ;
reg  KAC ;
reg  KAD ;
reg  KAE ;
reg  kba ;
reg  kbb ;
reg  kbc ;
reg  kbd ;
reg  KCA ;
reg  KCB ;
reg  KCC ;
reg  kda ;
reg  kdb ;
reg  kdc ;
reg  KEA ;
reg  KEB ;
reg  KEC ;
reg  kfa ;
reg  kfb ;
reg  KGA ;
reg  KGB ;
reg  KGC ;
reg  kha ;
reg  khb ;
reg  KIA ;
reg  KIB ;
reg  KIC ;
reg  KID ;
reg  kja ;
reg  kjb ;
reg  KKA ;
reg  KKB ;
reg  KKC ;
reg  KKD ;
reg  kla ;
reg  klb ;
reg  KMA ;
reg  KMB ;
reg  KMC ;
reg  KMD ;
reg  kna ;
reg  knb ;
reg  KOA ;
reg  KOB ;
reg  KOC ;
reg  KOD ;
reg  kpa ;
reg  kpb ;
reg  KQA ;
reg  KQB ;
reg  kra ;
reg  krb ;
reg  KSA ;
reg  KSB ;
reg  KSC ;
reg  kta ;
reg  ktb ;
reg  KUA ;
reg  KUB ;
reg  KUC ;
reg  MAA ;
reg  MAB ;
reg  MAC ;
reg  MAD ;
reg  mba ;
reg  mbb ;
reg  MCA ;
reg  MCB ;
reg  MCC ;
reg  mda ;
reg  MEA ;
reg  MEB ;
reg  mfa ;
reg  MGA ;
reg  MGB ;
reg  MGC ;
reg  mha ;
reg  MIA ;
reg  mja ;
reg  MKA ;
reg  MKB ;
reg  mla ;
reg  MMA ;
reg  MMB ;
reg  mna ;
reg  MOA ;
reg  MOB ;
reg  mpa ;
reg  MQA ;
reg  MQB ;
reg  mra ;
reg  MSA ;
reg  MSB ;
reg  mta ;
reg  MUA ;
reg  MUB ;
reg  oga ;
reg  ogb ;
reg  ogc ;
reg  ogd ;
reg  oge ;
reg  ogf ;
reg  ogg ;
reg  ogh ;
reg  ogi ;
reg  oha ;
reg  ohb ;
reg  ohc ;
reg  ohd ;
reg  OHE ;
reg  OHF ;
reg  oie ;
reg  oif ;
reg  oka ;
reg  okb ;
reg  OKC ;
reg  olc ;
reg  oma ;
reg  OMB ;
reg  OPA ;
reg  OPB ;
reg  OPC ;
reg  OPD ;
reg  OPE ;
reg  OPF ;
reg  OPG ;
reg  OPI ;
reg  OPK ;
reg  OPM ;
reg  OPO ;
reg  OPQ ;
reg  OPS ;
reg  OPU ;
reg  oqa ;
reg  oqc ;
reg  oqg ;
reg  oqi ;
reg  oqk ;
reg  oqm ;
reg  oqo ;
reg  oqq ;
reg  oqs ;
reg  oqu ;
reg  QIC ;
reg  QID ;
reg  QIE ;
reg  QIF ;
reg  QIG ;
reg  QIH ;
reg  QJA ;
reg  QJB ;
reg  QJC ;
reg  TAA ;
reg  TAB ;
wire  cal ;
wire  cam ;
wire  can ;
wire  cao ;
wire  cap ;
wire  cba ;
wire  cbb ;
wire  cbc ;
wire  cbd ;
wire  cbe ;
wire  cbf ;
wire  cbg ;
wire  cbh ;
wire  cbi ;
wire  cbj ;
wire  cbk ;
wire  cbl ;
wire  cbm ;
wire  cbn ;
wire  cbo ;
wire  cbp ;
wire  cca ;
wire  ccb ;
wire  ccc ;
wire  ccd ;
wire  cce ;
wire  ccf ;
wire  ccg ;
wire  cch ;
wire  cci ;
wire  ccj ;
wire  cck ;
wire  ccl ;
wire  ccm ;
wire  ccn ;
wire  cco ;
wire  ccp ;
wire  cdp ;
wire  cea ;
wire  ceb ;
wire  cec ;
wire  ced ;
wire  cee ;
wire  cef ;
wire  ceg ;
wire  ceh ;
wire  cei ;
wire  cej ;
wire  cek ;
wire  cel ;
wire  cem ;
wire  cen ;
wire  ceo ;
wire  cep ;
wire  cfa ;
wire  cfb ;
wire  cfc ;
wire  cfd ;
wire  cfe ;
wire  cff ;
wire  cfg ;
wire  cfh ;
wire  cfi ;
wire  cfj ;
wire  cfk ;
wire  cfl ;
wire  cfm ;
wire  cfn ;
wire  cfo ;
wire  cfp ;
wire  CGN ;
wire  CGO ;
wire  CGP ;
wire  CHA ;
wire  CHB ;
wire  CHC ;
wire  CHD ;
wire  CHE ;
wire  CHF ;
wire  CHG ;
wire  CHH ;
wire  CHI ;
wire  CHJ ;
wire  CHK ;
wire  CHL ;
wire  CHM ;
wire  CHN ;
wire  CHO ;
wire  CHP ;
wire  CIA ;
wire  CIB ;
wire  CIC ;
wire  CID ;
wire  CIE ;
wire  CIF ;
wire  CIG ;
wire  CIH ;
wire  CII ;
wire  CIJ ;
wire  CIK ;
wire  CIL ;
wire  CIM ;
wire  CIN ;
wire  CIO ;
wire  CIP ;
wire  CKI ;
wire  CKJ ;
wire  CKK ;
wire  CKL ;
wire  CKM ;
wire  CKN ;
wire  CKO ;
wire  CKP ;
wire  CLA ;
wire  CLB ;
wire  CLC ;
wire  CLD ;
wire  dal ;
wire  dam ;
wire  dan ;
wire  dao ;
wire  dap ;
wire  dba ;
wire  dbb ;
wire  dbc ;
wire  dbd ;
wire  dbe ;
wire  dbf ;
wire  dbg ;
wire  dbh ;
wire  dbi ;
wire  dbj ;
wire  dbk ;
wire  dbl ;
wire  dbm ;
wire  dbn ;
wire  dbo ;
wire  dbp ;
wire  dca ;
wire  dcb ;
wire  dcc ;
wire  dcd ;
wire  dce ;
wire  dcf ;
wire  dcg ;
wire  dch ;
wire  dci ;
wire  dcj ;
wire  dck ;
wire  dcl ;
wire  dcm ;
wire  dcn ;
wire  dco ;
wire  dcp ;
wire  ddo ;
wire  ddp ;
wire  dea ;
wire  deb ;
wire  dec ;
wire  ded ;
wire  dee ;
wire  def ;
wire  deg ;
wire  deh ;
wire  dei ;
wire  dej ;
wire  dek ;
wire  del ;
wire  dem ;
wire  den ;
wire  deo ;
wire  dep ;
wire  dfa ;
wire  dfb ;
wire  dfc ;
wire  dfd ;
wire  dfe ;
wire  dff ;
wire  dfg ;
wire  dfh ;
wire  dfi ;
wire  dfj ;
wire  dfk ;
wire  dfl ;
wire  dfm ;
wire  dfn ;
wire  dfo ;
wire  dfp ;
wire  DHA ;
wire  DHB ;
wire  DHC ;
wire  DHD ;
wire  DHE ;
wire  DHF ;
wire  DHG ;
wire  DHH ;
wire  DHI ;
wire  DHJ ;
wire  DHK ;
wire  DHL ;
wire  DHM ;
wire  DHN ;
wire  DHO ;
wire  DHP ;
wire  DIA ;
wire  DIB ;
wire  DIC ;
wire  DID ;
wire  DIE ;
wire  DIF ;
wire  DIG ;
wire  DIH ;
wire  DII ;
wire  DIJ ;
wire  DIK ;
wire  DIL ;
wire  DIM ;
wire  DIN ;
wire  DIO ;
wire  DIP ;
wire  eal ;
wire  EAL ;
wire  eam ;
wire  EAM ;
wire  ean ;
wire  EAN ;
wire  eao ;
wire  EAO ;
wire  eap ;
wire  EAP ;
wire  eaq ;
wire  EAQ ;
wire  ear ;
wire  EAR ;
wire  eas ;
wire  EAS ;
wire  eat ;
wire  EAT ;
wire  eau ;
wire  EAU ;
wire  eav ;
wire  EAV ;
wire  eaw ;
wire  EAW ;
wire  eax ;
wire  EAX ;
wire  eba ;
wire  EBA ;
wire  ebb ;
wire  EBB ;
wire  ebc ;
wire  EBC ;
wire  ebd ;
wire  EBD ;
wire  ebe ;
wire  EBE ;
wire  ebf ;
wire  EBF ;
wire  ebg ;
wire  EBG ;
wire  ebh ;
wire  EBH ;
wire  ebi ;
wire  EBI ;
wire  ebj ;
wire  EBJ ;
wire  ebk ;
wire  EBK ;
wire  ebl ;
wire  EBL ;
wire  ebm ;
wire  EBM ;
wire  ebn ;
wire  EBN ;
wire  ebo ;
wire  EBO ;
wire  ebp ;
wire  EBP ;
wire  ebq ;
wire  EBQ ;
wire  ebr ;
wire  EBR ;
wire  ebs ;
wire  EBS ;
wire  ebt ;
wire  EBT ;
wire  ebu ;
wire  EBU ;
wire  ebv ;
wire  EBV ;
wire  ebw ;
wire  EBW ;
wire  ebx ;
wire  EBX ;
wire  ecm ;
wire  ECM ;
wire  ecn ;
wire  ECN ;
wire  eco ;
wire  ECO ;
wire  ecp ;
wire  ECP ;
wire  ecq ;
wire  ECQ ;
wire  ecr ;
wire  ECR ;
wire  ecs ;
wire  ECS ;
wire  ect ;
wire  ECT ;
wire  ecu ;
wire  ECU ;
wire  ecv ;
wire  ECV ;
wire  ecw ;
wire  ECW ;
wire  ecx ;
wire  ECX ;
wire  eda ;
wire  EDA ;
wire  edb ;
wire  EDB ;
wire  edc ;
wire  EDC ;
wire  edd ;
wire  EDD ;
wire  ede ;
wire  EDE ;
wire  edf ;
wire  EDF ;
wire  edg ;
wire  EDG ;
wire  edh ;
wire  EDH ;
wire  edi ;
wire  EDI ;
wire  edj ;
wire  EDJ ;
wire  edk ;
wire  EDK ;
wire  edl ;
wire  EDL ;
wire  edm ;
wire  EDM ;
wire  edn ;
wire  EDN ;
wire  edo ;
wire  EDO ;
wire  edp ;
wire  EDP ;
wire  edq ;
wire  EDQ ;
wire  edr ;
wire  EDR ;
wire  eds ;
wire  EDS ;
wire  edt ;
wire  EDT ;
wire  edu ;
wire  EDU ;
wire  edv ;
wire  EDV ;
wire  edw ;
wire  EDW ;
wire  edx ;
wire  EDX ;
wire  een ;
wire  EEN ;
wire  eeo ;
wire  EEO ;
wire  eep ;
wire  EEP ;
wire  eeq ;
wire  EEQ ;
wire  eer ;
wire  EER ;
wire  ees ;
wire  EES ;
wire  eet ;
wire  EET ;
wire  eeu ;
wire  EEU ;
wire  eev ;
wire  EEV ;
wire  eew ;
wire  EEW ;
wire  eex ;
wire  EEX ;
wire  efa ;
wire  EFA ;
wire  efb ;
wire  EFB ;
wire  efc ;
wire  EFC ;
wire  efd ;
wire  EFD ;
wire  efe ;
wire  EFE ;
wire  eff ;
wire  EFF ;
wire  efg ;
wire  EFG ;
wire  efh ;
wire  EFH ;
wire  efi ;
wire  EFI ;
wire  efj ;
wire  EFJ ;
wire  efk ;
wire  EFK ;
wire  efl ;
wire  EFL ;
wire  efm ;
wire  EFM ;
wire  efn ;
wire  EFN ;
wire  efo ;
wire  EFO ;
wire  efp ;
wire  EFP ;
wire  efq ;
wire  EFQ ;
wire  efr ;
wire  EFR ;
wire  efs ;
wire  EFS ;
wire  eft ;
wire  EFT ;
wire  efu ;
wire  EFU ;
wire  efv ;
wire  EFV ;
wire  efw ;
wire  EFW ;
wire  efx ;
wire  EFX ;
wire  ego ;
wire  EGO ;
wire  egp ;
wire  EGP ;
wire  egq ;
wire  EGQ ;
wire  egr ;
wire  EGR ;
wire  egs ;
wire  EGS ;
wire  egt ;
wire  EGT ;
wire  egu ;
wire  EGU ;
wire  egv ;
wire  EGV ;
wire  egw ;
wire  EGW ;
wire  egx ;
wire  EGX ;
wire  eha ;
wire  EHA ;
wire  ehb ;
wire  EHB ;
wire  ehc ;
wire  EHC ;
wire  ehd ;
wire  EHD ;
wire  ehe ;
wire  EHE ;
wire  ehf ;
wire  EHF ;
wire  ehg ;
wire  EHG ;
wire  ehh ;
wire  EHH ;
wire  ehi ;
wire  EHI ;
wire  ehj ;
wire  EHJ ;
wire  ehk ;
wire  EHK ;
wire  ehl ;
wire  EHL ;
wire  ehm ;
wire  EHM ;
wire  ehn ;
wire  EHN ;
wire  eho ;
wire  EHO ;
wire  ehp ;
wire  EHP ;
wire  ehq ;
wire  EHQ ;
wire  ehr ;
wire  EHR ;
wire  ehs ;
wire  EHS ;
wire  eht ;
wire  EHT ;
wire  ehu ;
wire  EHU ;
wire  ehv ;
wire  EHV ;
wire  ehw ;
wire  EHW ;
wire  ehx ;
wire  EHX ;
wire  eip ;
wire  EIP ;
wire  eiq ;
wire  EIQ ;
wire  eir ;
wire  EIR ;
wire  eis ;
wire  EIS ;
wire  eit ;
wire  EIT ;
wire  eiu ;
wire  EIU ;
wire  eiv ;
wire  EIV ;
wire  eiw ;
wire  EIW ;
wire  eix ;
wire  EIX ;
wire  eja ;
wire  EJA ;
wire  ejb ;
wire  EJB ;
wire  ejc ;
wire  EJC ;
wire  ejd ;
wire  EJD ;
wire  eje ;
wire  EJE ;
wire  ejf ;
wire  EJF ;
wire  ejg ;
wire  EJG ;
wire  ejh ;
wire  EJH ;
wire  eji ;
wire  EJI ;
wire  ejj ;
wire  EJJ ;
wire  ejk ;
wire  EJK ;
wire  ejl ;
wire  EJL ;
wire  ejm ;
wire  EJM ;
wire  ejn ;
wire  EJN ;
wire  ejo ;
wire  EJO ;
wire  ejp ;
wire  EJP ;
wire  ejq ;
wire  EJQ ;
wire  ejr ;
wire  EJR ;
wire  ejs ;
wire  EJS ;
wire  ejt ;
wire  EJT ;
wire  eju ;
wire  EJU ;
wire  ejv ;
wire  EJV ;
wire  ejw ;
wire  EJW ;
wire  ejx ;
wire  EJX ;
wire  ekq ;
wire  EKQ ;
wire  ekr ;
wire  EKR ;
wire  eks ;
wire  EKS ;
wire  ekt ;
wire  EKT ;
wire  eku ;
wire  EKU ;
wire  ekv ;
wire  EKV ;
wire  ekw ;
wire  EKW ;
wire  ekx ;
wire  EKX ;
wire  ela ;
wire  ELA ;
wire  elb ;
wire  ELB ;
wire  elc ;
wire  ELC ;
wire  eld ;
wire  ELD ;
wire  ele ;
wire  ELE ;
wire  elf ;
wire  ELF ;
wire  elg ;
wire  ELG ;
wire  elh ;
wire  ELH ;
wire  eli ;
wire  ELI ;
wire  elj ;
wire  ELJ ;
wire  elk ;
wire  ELK ;
wire  ell ;
wire  ELL ;
wire  elm ;
wire  ELM ;
wire  eln ;
wire  ELN ;
wire  elo ;
wire  ELO ;
wire  elp ;
wire  ELP ;
wire  elq ;
wire  ELQ ;
wire  elr ;
wire  ELR ;
wire  els ;
wire  ELS ;
wire  elt ;
wire  ELT ;
wire  elu ;
wire  ELU ;
wire  elv ;
wire  ELV ;
wire  elw ;
wire  ELW ;
wire  elx ;
wire  ELX ;
wire  emr ;
wire  EMR ;
wire  ems ;
wire  EMS ;
wire  emt ;
wire  EMT ;
wire  emu ;
wire  EMU ;
wire  emv ;
wire  EMV ;
wire  emw ;
wire  EMW ;
wire  emx ;
wire  EMX ;
wire  ena ;
wire  ENA ;
wire  enb ;
wire  ENB ;
wire  enc ;
wire  ENC ;
wire  endd ;
wire  ENDD  ;
wire  ene ;
wire  ENE ;
wire  enf ;
wire  ENF ;
wire  eng ;
wire  ENG ;
wire  enh ;
wire  ENH ;
wire  eni ;
wire  ENI ;
wire  enj ;
wire  ENJ ;
wire  enk ;
wire  ENK ;
wire  enl ;
wire  ENL ;
wire  enm ;
wire  ENM ;
wire  enn ;
wire  ENN ;
wire  eno ;
wire  ENO ;
wire  enp ;
wire  ENP ;
wire  enq ;
wire  ENQ ;
wire  enr ;
wire  ENR ;
wire  ens ;
wire  ENS ;
wire  ent ;
wire  ENT ;
wire  enu ;
wire  ENU ;
wire  env ;
wire  ENV ;
wire  enw ;
wire  ENW ;
wire  enx ;
wire  ENX ;
wire  eos ;
wire  EOS ;
wire  eot ;
wire  EOT ;
wire  eou ;
wire  EOU ;
wire  eov ;
wire  EOV ;
wire  eow ;
wire  EOW ;
wire  eox ;
wire  EOX ;
wire  epa ;
wire  EPA ;
wire  epb ;
wire  EPB ;
wire  epc ;
wire  EPC ;
wire  epd ;
wire  EPD ;
wire  epe ;
wire  EPE ;
wire  epf ;
wire  EPF ;
wire  epg ;
wire  EPG ;
wire  eph ;
wire  EPH ;
wire  epi ;
wire  EPI ;
wire  epj ;
wire  EPJ ;
wire  epk ;
wire  EPK ;
wire  epl ;
wire  EPL ;
wire  epm ;
wire  EPM ;
wire  epn ;
wire  EPN ;
wire  epo ;
wire  EPO ;
wire  epp ;
wire  EPP ;
wire  epq ;
wire  EPQ ;
wire  epr ;
wire  EPR ;
wire  eps ;
wire  EPS ;
wire  ept ;
wire  EPT ;
wire  epu ;
wire  EPU ;
wire  epv ;
wire  EPV ;
wire  epw ;
wire  EPW ;
wire  epx ;
wire  EPX ;
wire  eqt ;
wire  EQT ;
wire  equ ;
wire  EQU ;
wire  eqv ;
wire  EQV ;
wire  eqw ;
wire  EQW ;
wire  eqx ;
wire  EQX ;
wire  era ;
wire  ERA ;
wire  erb ;
wire  ERB ;
wire  erc ;
wire  ERC ;
wire  erd ;
wire  ERD ;
wire  ere ;
wire  ERE ;
wire  erf ;
wire  ERF ;
wire  erg ;
wire  ERG ;
wire  erh ;
wire  ERH ;
wire  eri ;
wire  ERI ;
wire  erj ;
wire  ERJ ;
wire  erk ;
wire  ERK ;
wire  erl ;
wire  ERL ;
wire  erm ;
wire  ERM ;
wire  ern ;
wire  ERN ;
wire  ero ;
wire  ERO ;
wire  erp ;
wire  ERP ;
wire  erq ;
wire  ERQ ;
wire  err ;
wire  ERR ;
wire  ers ;
wire  ERS ;
wire  ert ;
wire  ERT ;
wire  eru ;
wire  ERU ;
wire  erv ;
wire  ERV ;
wire  erw ;
wire  ERW ;
wire  erx ;
wire  ERX ;
wire  esu ;
wire  ESU ;
wire  esv ;
wire  ESV ;
wire  esw ;
wire  ESW ;
wire  esx ;
wire  ESX ;
wire  eta ;
wire  ETA ;
wire  etb ;
wire  ETB ;
wire  etc ;
wire  ETC ;
wire  etd ;
wire  ETD ;
wire  ete ;
wire  ETE ;
wire  etf ;
wire  ETF ;
wire  etg ;
wire  ETG ;
wire  eth ;
wire  ETH ;
wire  eti ;
wire  ETI ;
wire  etj ;
wire  ETJ ;
wire  etk ;
wire  ETK ;
wire  etl ;
wire  ETL ;
wire  etm ;
wire  ETM ;
wire  etn ;
wire  ETN ;
wire  eto ;
wire  ETO ;
wire  etp ;
wire  ETP ;
wire  etq ;
wire  ETQ ;
wire  etr ;
wire  ETR ;
wire  ets ;
wire  ETS ;
wire  ett ;
wire  ETT ;
wire  etu ;
wire  ETU ;
wire  etv ;
wire  ETV ;
wire  etw ;
wire  ETW ;
wire  etx ;
wire  ETX ;
wire  euv ;
wire  EUV ;
wire  euw ;
wire  EUW ;
wire  eux ;
wire  EUX ;
wire  eva ;
wire  EVA ;
wire  evb ;
wire  EVB ;
wire  evc ;
wire  EVC ;
wire  evd ;
wire  EVD ;
wire  eve ;
wire  EVE ;
wire  evf ;
wire  EVF ;
wire  evg ;
wire  EVG ;
wire  evh ;
wire  EVH ;
wire  evi ;
wire  EVI ;
wire  evj ;
wire  EVJ ;
wire  evk ;
wire  EVK ;
wire  evl ;
wire  EVL ;
wire  evm ;
wire  EVM ;
wire  evn ;
wire  EVN ;
wire  evo ;
wire  EVO ;
wire  evp ;
wire  EVP ;
wire  evq ;
wire  EVQ ;
wire  evr ;
wire  EVR ;
wire  evs ;
wire  EVS ;
wire  evt ;
wire  EVT ;
wire  evu ;
wire  EVU ;
wire  evv ;
wire  EVV ;
wire  evw ;
wire  EVW ;
wire  evx ;
wire  EVX ;
wire  faa ;
wire  fab ;
wire  fac ;
wire  fad ;
wire  fae ;
wire  faf ;
wire  fag ;
wire  fah ;
wire  fai ;
wire  faj ;
wire  fak ;
wire  fal ;
wire  fam ;
wire  fan ;
wire  FBA ;
wire  FBB ;
wire  FBC ;
wire  FBD ;
wire  FBE ;
wire  FBF ;
wire  FBG ;
wire  FBH ;
wire  FBI ;
wire  FBJ ;
wire  FBK ;
wire  FBL ;
wire  fca ;
wire  fcb ;
wire  fcc ;
wire  fcd ;
wire  fce ;
wire  fcf ;
wire  fcg ;
wire  fch ;
wire  fci ;
wire  fcj ;
wire  fck ;
wire  fcl ;
wire  fcm ;
wire  FDA ;
wire  FDB ;
wire  FDC ;
wire  FDD ;
wire  FDE ;
wire  FDF ;
wire  FDG ;
wire  FDH ;
wire  FDI ;
wire  FDJ ;
wire  FDK ;
wire  FDL ;
wire  fea ;
wire  feb ;
wire  fec ;
wire  fed ;
wire  fee ;
wire  fef ;
wire  feg ;
wire  feh ;
wire  fei ;
wire  fej ;
wire  fek ;
wire  fel ;
wire  FFA ;
wire  FFB ;
wire  FFC ;
wire  FFD ;
wire  FFE ;
wire  FFF ;
wire  FFG ;
wire  FFH ;
wire  FFI ;
wire  FFJ ;
wire  FFK ;
wire  FFL ;
wire  fga ;
wire  fgb ;
wire  fgc ;
wire  fgd ;
wire  fge ;
wire  fgf ;
wire  fgg ;
wire  fgh ;
wire  fgi ;
wire  fgj ;
wire  fgk ;
wire  fgl ;
wire  fgm ;
wire  FHA ;
wire  FHB ;
wire  FHC ;
wire  FHD ;
wire  FHE ;
wire  FHF ;
wire  FHG ;
wire  FHH ;
wire  FHI ;
wire  FHJ ;
wire  FHK ;
wire  fia ;
wire  fib ;
wire  fic ;
wire  fid ;
wire  fie ;
wire  fif ;
wire  fig ;
wire  fih ;
wire  fii ;
wire  fij ;
wire  fik ;
wire  fil ;
wire  FJA ;
wire  FJB ;
wire  FJC ;
wire  FJD ;
wire  FJE ;
wire  FJF ;
wire  FJG ;
wire  FJH ;
wire  FJI ;
wire  FJJ ;
wire  FJK ;
wire  fka ;
wire  fkb ;
wire  fkc ;
wire  fkd ;
wire  fke ;
wire  fkf ;
wire  fkg ;
wire  fkh ;
wire  fki ;
wire  fkj ;
wire  fkk ;
wire  FLA ;
wire  FLB ;
wire  FLC ;
wire  FLD ;
wire  FLE ;
wire  FLF ;
wire  FLG ;
wire  FLH ;
wire  FLI ;
wire  FLJ ;
wire  FLK ;
wire  fma ;
wire  fmb ;
wire  fmc ;
wire  fmd ;
wire  fme ;
wire  fmf ;
wire  fmg ;
wire  fmh ;
wire  fmi ;
wire  fmj ;
wire  fmk ;
wire  fml ;
wire  FNA ;
wire  FNB ;
wire  FNC ;
wire  FND ;
wire  FNE ;
wire  FNF ;
wire  FNG ;
wire  FNH ;
wire  FNI ;
wire  FNJ ;
wire  foa ;
wire  fob ;
wire  foc ;
wire  fod ;
wire  foe ;
wire  fof ;
wire  fog ;
wire  foh ;
wire  foi ;
wire  foj ;
wire  fok ;
wire  FPA ;
wire  FPB ;
wire  FPC ;
wire  FPD ;
wire  FPE ;
wire  FPF ;
wire  FPG ;
wire  FPH ;
wire  FPI ;
wire  FPJ ;
wire  fqa ;
wire  fqb ;
wire  fqc ;
wire  fqd ;
wire  fqe ;
wire  fqf ;
wire  fqg ;
wire  fqh ;
wire  fqi ;
wire  fqj ;
wire  FRA ;
wire  FRB ;
wire  FRC ;
wire  FRD ;
wire  FRE ;
wire  FRF ;
wire  FRG ;
wire  FRH ;
wire  FRI ;
wire  FRJ ;
wire  fsa ;
wire  fsb ;
wire  fsc ;
wire  fsd ;
wire  fse ;
wire  fsf ;
wire  fsg ;
wire  fsh ;
wire  fsi ;
wire  fsj ;
wire  fsk ;
wire  FTA ;
wire  FTB ;
wire  FTC ;
wire  FTD ;
wire  FTE ;
wire  FTF ;
wire  FTG ;
wire  FTH ;
wire  FTI ;
wire  fua ;
wire  fub ;
wire  fuc ;
wire  fud ;
wire  fue ;
wire  fuf ;
wire  fug ;
wire  fuh ;
wire  fui ;
wire  fuj ;
wire  gaa ;
wire  GAA ;
wire  gab ;
wire  GAB ;
wire  gac ;
wire  GAC ;
wire  gad ;
wire  GAD ;
wire  gba ;
wire  GBA ;
wire  gbb ;
wire  GBB ;
wire  gbc ;
wire  GBC ;
wire  gbd ;
wire  GBD ;
wire  gca ;
wire  GCA ;
wire  gcb ;
wire  GCB ;
wire  gcc ;
wire  GCC ;
wire  gcd ;
wire  GCD ;
wire  gce ;
wire  GCE ;
wire  gcf ;
wire  GCF ;
wire  gcg ;
wire  GCG ;
wire  gch ;
wire  GCH ;
wire  gda ;
wire  GDA ;
wire  gdb ;
wire  GDB ;
wire  gdc ;
wire  GDC ;
wire  gdd ;
wire  GDD ;
wire  gde ;
wire  GDE ;
wire  gdf ;
wire  GDF ;
wire  gdg ;
wire  GDG ;
wire  gdh ;
wire  GDH ;
wire  gea ;
wire  GEA ;
wire  geb ;
wire  GEB ;
wire  gec ;
wire  GEC ;
wire  ged ;
wire  GED ;
wire  gee ;
wire  GEE ;
wire  gef ;
wire  GEF ;
wire  geg ;
wire  GEG ;
wire  geh ;
wire  GEH ;
wire  gfa ;
wire  GFA ;
wire  gfb ;
wire  GFB ;
wire  gfc ;
wire  GFC ;
wire  gfd ;
wire  GFD ;
wire  gfe ;
wire  GFE ;
wire  gff ;
wire  GFF ;
wire  gfg ;
wire  GFG ;
wire  gfh ;
wire  GFH ;
wire  gga ;
wire  GGA ;
wire  ggb ;
wire  GGB ;
wire  ggc ;
wire  GGC ;
wire  ggd ;
wire  GGD ;
wire  gge ;
wire  GGE ;
wire  ggf ;
wire  GGF ;
wire  ggg ;
wire  GGG ;
wire  ggh ;
wire  GGH ;
wire  gha ;
wire  GHA ;
wire  ghb ;
wire  GHB ;
wire  ghc ;
wire  GHC ;
wire  ghd ;
wire  GHD ;
wire  ghe ;
wire  GHE ;
wire  ghf ;
wire  GHF ;
wire  ghg ;
wire  GHG ;
wire  ghh ;
wire  GHH ;
wire  gia ;
wire  GIA ;
wire  gib ;
wire  GIB ;
wire  gic ;
wire  GIC ;
wire  gid ;
wire  GID ;
wire  gie ;
wire  GIE ;
wire  gif ;
wire  GIF ;
wire  gig ;
wire  GIG ;
wire  gja ;
wire  GJA ;
wire  gjb ;
wire  GJB ;
wire  gjc ;
wire  GJC ;
wire  gjd ;
wire  GJD ;
wire  gje ;
wire  GJE ;
wire  gjf ;
wire  GJF ;
wire  gjg ;
wire  GJG ;
wire  gka ;
wire  GKA ;
wire  gkb ;
wire  GKB ;
wire  gkc ;
wire  GKC ;
wire  gkd ;
wire  GKD ;
wire  gke ;
wire  GKE ;
wire  gkf ;
wire  GKF ;
wire  gkg ;
wire  GKG ;
wire  gla ;
wire  GLA ;
wire  glb ;
wire  GLB ;
wire  glc ;
wire  GLC ;
wire  gld ;
wire  GLD ;
wire  gle ;
wire  GLE ;
wire  glf ;
wire  GLF ;
wire  glg ;
wire  GLG ;
wire  gma ;
wire  GMA ;
wire  gmb ;
wire  GMB ;
wire  gmc ;
wire  GMC ;
wire  gmd ;
wire  GMD ;
wire  gme ;
wire  GME ;
wire  gmf ;
wire  GMF ;
wire  gmg ;
wire  GMG ;
wire  gna ;
wire  GNA ;
wire  gnb ;
wire  GNB ;
wire  gnc ;
wire  GNC ;
wire  gnd ;
wire  GND ;
wire  gne ;
wire  GNE ;
wire  gnf ;
wire  GNF ;
wire  gng ;
wire  GNG ;
wire  goa ;
wire  GOA ;
wire  gob ;
wire  GOB ;
wire  goc ;
wire  GOC ;
wire  god ;
wire  GOD ;
wire  goe ;
wire  GOE ;
wire  gof ;
wire  GOF ;
wire  gog ;
wire  GOG ;
wire  gpa ;
wire  GPA ;
wire  gpb ;
wire  GPB ;
wire  gpc ;
wire  GPC ;
wire  gpd ;
wire  GPD ;
wire  gpe ;
wire  GPE ;
wire  gpf ;
wire  GPF ;
wire  gpg ;
wire  GPG ;
wire  gqa ;
wire  GQA ;
wire  gqb ;
wire  GQB ;
wire  gqc ;
wire  GQC ;
wire  gqd ;
wire  GQD ;
wire  gqe ;
wire  GQE ;
wire  gqf ;
wire  GQF ;
wire  gra ;
wire  GRA ;
wire  grb ;
wire  GRB ;
wire  grc ;
wire  GRC ;
wire  grd ;
wire  GRD ;
wire  gre ;
wire  GRE ;
wire  grf ;
wire  GRF ;
wire  gsa ;
wire  GSA ;
wire  gsb ;
wire  GSB ;
wire  gsc ;
wire  GSC ;
wire  gsd ;
wire  GSD ;
wire  gse ;
wire  GSE ;
wire  gsf ;
wire  GSF ;
wire  gsg ;
wire  GSG ;
wire  gta ;
wire  GTA ;
wire  gtb ;
wire  GTB ;
wire  gtc ;
wire  GTC ;
wire  gtd ;
wire  GTD ;
wire  gte ;
wire  GTE ;
wire  gtf ;
wire  GTF ;
wire  gtg ;
wire  GTG ;
wire  gua ;
wire  GUA ;
wire  gub ;
wire  GUB ;
wire  guc ;
wire  GUC ;
wire  gud ;
wire  GUD ;
wire  gue ;
wire  GUE ;
wire  guf ;
wire  GUF ;
wire  gva ;
wire  GVA ;
wire  gvb ;
wire  GVB ;
wire  gvc ;
wire  GVC ;
wire  gvd ;
wire  GVD ;
wire  gve ;
wire  GVE ;
wire  gvf ;
wire  GVF ;
wire  haa ;
wire  hab ;
wire  hac ;
wire  had ;
wire  hae ;
wire  haf ;
wire  hag ;
wire  HBA ;
wire  HBB ;
wire  HBC ;
wire  HBD ;
wire  HBE ;
wire  HBF ;
wire  hca ;
wire  hcb ;
wire  hcc ;
wire  hcd ;
wire  hce ;
wire  HDA ;
wire  HDB ;
wire  HDC ;
wire  HDD ;
wire  hea ;
wire  heb ;
wire  hec ;
wire  hed ;
wire  hee ;
wire  hef ;
wire  HFA ;
wire  HFB ;
wire  HFC ;
wire  HFD ;
wire  HFE ;
wire  hga ;
wire  hgb ;
wire  hgc ;
wire  hgd ;
wire  hge ;
wire  hgf ;
wire  hgg ;
wire  HHA ;
wire  HHB ;
wire  HHC ;
wire  HHD ;
wire  HHE ;
wire  hia ;
wire  hib ;
wire  hic ;
wire  hid ;
wire  hie ;
wire  hif ;
wire  hig ;
wire  HJA ;
wire  HJB ;
wire  HJC ;
wire  HJD ;
wire  HJE ;
wire  hka ;
wire  hkb ;
wire  hkc ;
wire  hkd ;
wire  hke ;
wire  HLA ;
wire  HLB ;
wire  HLC ;
wire  HLD ;
wire  HLE ;
wire  hma ;
wire  hmb ;
wire  hmc ;
wire  hmd ;
wire  hme ;
wire  hmf ;
wire  HNA ;
wire  HNB ;
wire  HNC ;
wire  HND ;
wire  HNE ;
wire  hoa ;
wire  hob ;
wire  hoc ;
wire  hod ;
wire  hoe ;
wire  hof ;
wire  HPA ;
wire  HPB ;
wire  HPC ;
wire  HPD ;
wire  hqa ;
wire  hqb ;
wire  hqc ;
wire  hqd ;
wire  hqe ;
wire  HRA ;
wire  HRB ;
wire  HRC ;
wire  HRD ;
wire  HRE ;
wire  hsa ;
wire  hsb ;
wire  hsc ;
wire  hsd ;
wire  hse ;
wire  HTA ;
wire  HTB ;
wire  HTC ;
wire  HTD ;
wire  hua ;
wire  hub ;
wire  huc ;
wire  hud ;
wire  hue ;
wire  huf ;
wire  ial ;
wire  iam ;
wire  ian ;
wire  iao ;
wire  iap ;
wire  iba ;
wire  ibb ;
wire  ibc ;
wire  ibd ;
wire  ibe ;
wire  ibf ;
wire  ibg ;
wire  ibh ;
wire  ibi ;
wire  ibj ;
wire  ibk ;
wire  ibl ;
wire  ibm ;
wire  ibn ;
wire  ibo ;
wire  ibp ;
wire  ica ;
wire  icb ;
wire  icc ;
wire  icd ;
wire  ice ;
wire  icf ;
wire  icg ;
wire  ich ;
wire  ici ;
wire  icj ;
wire  ick ;
wire  icl ;
wire  icm ;
wire  icn ;
wire  ico ;
wire  icp ;
wire  idl ;
wire  idm ;
wire  idn ;
wire  ido ;
wire  idp ;
wire  iea ;
wire  ieb ;
wire  iec ;
wire  ied ;
wire  iee ;
wire  ief ;
wire  ieg ;
wire  ieh ;
wire  iei ;
wire  iej ;
wire  iek ;
wire  iel ;
wire  iem ;
wire  ien ;
wire  ieo ;
wire  iep ;
wire  ifa ;
wire  ifb ;
wire  ifc ;
wire  ifd ;
wire  ife ;
wire  ifff  ;
wire  ifg ;
wire  ifh ;
wire  ifi ;
wire  ifj ;
wire  ifk ;
wire  ifl ;
wire  ifm ;
wire  ifn ;
wire  ifo ;
wire  ifp ;
wire  iga ;
wire  igb ;
wire  igc ;
wire  igd ;
wire  ige ;
wire  igf ;
wire  igg ;
wire  igh ;
wire  igi ;
wire  igj ;
wire  ila ;
wire  ilb ;
wire  ilc ;
wire  ild ;
wire  ile ;
wire  ilf ;
wire  ilg ;
wire  ilh ;
wire  ili ;
wire  ilj ;
wire  ilk ;
wire  ill ;
wire  ilm ;
wire  ima ;
wire  imb ;
wire  imc ;
wire  imd ;
wire  ime ;
wire  imf ;
wire  img ;
wire  imh ;
wire  imi ;
wire  imj ;
wire  imk ;
wire  iml ;
wire  ina ;
wire  inb ;
wire  inc ;
wire  ind ;
wire  ine ;
wire  inf ;
wire  ioa ;
wire  iob ;
wire  iqc ;
wire  iqd ;
wire  iqe ;
wire  iqf ;
wire  iqg ;
wire  iqh ;
wire  ira ;
wire  irb ;
wire  irc ;
wire  jaa ;
wire  JAA ;
wire  jab ;
wire  JAB ;
wire  jba ;
wire  JBA ;
wire  jbb ;
wire  JBB ;
wire  jca ;
wire  JCA ;
wire  jcb ;
wire  JCB ;
wire  jcc ;
wire  JCC ;
wire  jda ;
wire  JDA ;
wire  jdb ;
wire  JDB ;
wire  jdc ;
wire  JDC ;
wire  jea ;
wire  JEA ;
wire  jeb ;
wire  JEB ;
wire  jec ;
wire  JEC ;
wire  jfa ;
wire  JFA ;
wire  jfb ;
wire  JFB ;
wire  jfc ;
wire  JFC ;
wire  jga ;
wire  JGA ;
wire  jgb ;
wire  JGB ;
wire  jgc ;
wire  JGC ;
wire  jgd ;
wire  JGD ;
wire  jha ;
wire  JHA ;
wire  jhb ;
wire  JHB ;
wire  jhc ;
wire  JHC ;
wire  jhd ;
wire  JHD ;
wire  jia ;
wire  JIA ;
wire  jib ;
wire  JIB ;
wire  jic ;
wire  JIC ;
wire  jid ;
wire  JID ;
wire  jja ;
wire  JJA ;
wire  jjb ;
wire  JJB ;
wire  jjc ;
wire  JJC ;
wire  jjd ;
wire  JJD ;
wire  jka ;
wire  JKA ;
wire  jkb ;
wire  JKB ;
wire  jkc ;
wire  JKC ;
wire  jla ;
wire  JLA ;
wire  jlb ;
wire  JLB ;
wire  jlc ;
wire  JLC ;
wire  jma ;
wire  JMA ;
wire  jmb ;
wire  JMB ;
wire  jmc ;
wire  JMC ;
wire  jna ;
wire  JNA ;
wire  jnb ;
wire  JNB ;
wire  jnc ;
wire  JNC ;
wire  joa ;
wire  JOA ;
wire  job ;
wire  JOB ;
wire  joc ;
wire  JOC ;
wire  jpa ;
wire  JPA ;
wire  jpb ;
wire  JPB ;
wire  jpc ;
wire  JPC ;
wire  jqa ;
wire  JQA ;
wire  jqb ;
wire  JQB ;
wire  jqc ;
wire  JQC ;
wire  jra ;
wire  JRA ;
wire  jrb ;
wire  JRB ;
wire  jrc ;
wire  JRC ;
wire  jsa ;
wire  JSA ;
wire  jsb ;
wire  JSB ;
wire  jsc ;
wire  JSC ;
wire  jta ;
wire  JTA ;
wire  jtb ;
wire  JTB ;
wire  jtc ;
wire  JTC ;
wire  jua ;
wire  JUA ;
wire  jub ;
wire  JUB ;
wire  juc ;
wire  JUC ;
wire  jva ;
wire  JVA ;
wire  jvb ;
wire  JVB ;
wire  jvc ;
wire  JVC ;
wire  kaa ;
wire  kab ;
wire  kac ;
wire  kad ;
wire  kae ;
wire  KBA ;
wire  KBB ;
wire  KBC ;
wire  KBD ;
wire  kca ;
wire  kcb ;
wire  kcc ;
wire  KDA ;
wire  KDB ;
wire  KDC ;
wire  kea ;
wire  keb ;
wire  kec ;
wire  KFA ;
wire  KFB ;
wire  kga ;
wire  kgb ;
wire  kgc ;
wire  KHA ;
wire  KHB ;
wire  kia ;
wire  kib ;
wire  kic ;
wire  kid ;
wire  KJA ;
wire  KJB ;
wire  kka ;
wire  kkb ;
wire  kkc ;
wire  kkd ;
wire  KLA ;
wire  KLB ;
wire  kma ;
wire  kmb ;
wire  kmc ;
wire  kmd ;
wire  KNA ;
wire  KNB ;
wire  koa ;
wire  kob ;
wire  koc ;
wire  kod ;
wire  KPA ;
wire  KPB ;
wire  kqa ;
wire  kqb ;
wire  KRA ;
wire  KRB ;
wire  ksa ;
wire  ksb ;
wire  ksc ;
wire  KTA ;
wire  KTB ;
wire  kua ;
wire  kub ;
wire  kuc ;
wire  laa ;
wire  LAA ;
wire  lba ;
wire  LBA ;
wire  lca ;
wire  LCA ;
wire  lcb ;
wire  LCB ;
wire  lda ;
wire  LDA ;
wire  ldb ;
wire  LDB ;
wire  lea ;
wire  LEA ;
wire  leb ;
wire  LEB ;
wire  lfa ;
wire  LFA ;
wire  lfb ;
wire  LFB ;
wire  lga ;
wire  LGA ;
wire  lha ;
wire  LHA ;
wire  lia ;
wire  LIA ;
wire  lib ;
wire  LIB ;
wire  lja ;
wire  LJA ;
wire  ljb ;
wire  LJB ;
wire  lka ;
wire  LKA ;
wire  lkb ;
wire  LKB ;
wire  lla ;
wire  LLA ;
wire  llb ;
wire  LLB ;
wire  lma ;
wire  LMA ;
wire  lmb ;
wire  LMB ;
wire  lna ;
wire  LNA ;
wire  lnb ;
wire  LNB ;
wire  loa ;
wire  LOA ;
wire  lob ;
wire  LOB ;
wire  lpa ;
wire  LPA ;
wire  lpb ;
wire  LPB ;
wire  lqa ;
wire  LQA ;
wire  lra ;
wire  LRA ;
wire  lsa ;
wire  LSA ;
wire  lta ;
wire  LTA ;
wire  lua ;
wire  LUA ;
wire  lva ;
wire  LVA ;
wire  maa ;
wire  mab ;
wire  mac ;
wire  mad ;
wire  MBA ;
wire  MBB ;
wire  mca ;
wire  mcb ;
wire  mcc ;
wire  MDA ;
wire  mea ;
wire  meb ;
wire  MFA ;
wire  mga ;
wire  mgb ;
wire  mgc ;
wire  MHA ;
wire  mia ;
wire  MJA ;
wire  mka ;
wire  mkb ;
wire  MLA ;
wire  mma ;
wire  mmb ;
wire  MNA ;
wire  moa ;
wire  mob ;
wire  MPA ;
wire  mqa ;
wire  mqb ;
wire  MRA ;
wire  msa ;
wire  msb ;
wire  MTA ;
wire  mua ;
wire  mub ;
wire  naa ;
wire  NAA ;
wire  nba ;
wire  NBA ;
wire  nca ;
wire  NCA ;
wire  nda ;
wire  NDA ;
wire  nea ;
wire  NEA ;
wire  nfa ;
wire  NFA ;
wire  nga ;
wire  NGA ;
wire  nha ;
wire  NHA ;
wire  OGA ;
wire  OGB ;
wire  OGC ;
wire  OGD ;
wire  OGE ;
wire  OGF ;
wire  OGG ;
wire  OGH ;
wire  OGI ;
wire  OHA ;
wire  OHB ;
wire  OHC ;
wire  OHD ;
wire  ohe ;
wire  ohf ;
wire  OIE ;
wire  OIF ;
wire  OKA ;
wire  OKB ;
wire  okc ;
wire  OLC ;
wire  OMA ;
wire  omb ;
wire  opa ;
wire  opb ;
wire  opc ;
wire  opd ;
wire  ope ;
wire  opf ;
wire  opg ;
wire  opi ;
wire  opk ;
wire  opm ;
wire  opo ;
wire  opq ;
wire  ops ;
wire  opu ;
wire  OQA ;
wire  OQC ;
wire  OQG ;
wire  OQI ;
wire  OQK ;
wire  OQM ;
wire  OQO ;
wire  OQQ ;
wire  OQS ;
wire  OQU ;
wire  qic ;
wire  qid ;
wire  qie ;
wire  qif ;
wire  qig ;
wire  qih ;
wire  qja ;
wire  qjb ;
wire  qjc ;
wire  taa ;
wire  tab ;
wire  ZZI ;
wire  ZZO ;
assign ZZI = 1'b1;
assign ZZO = 1'b0;
assign LAA =  KAA & kae & kab  |  kaa & KAE & kab  |  kaa & kae & KAB  |  KAA & KAE & KAB  ; 
assign laa = ~LAA; //complement 
assign lba =  KAA & kae & kab  |  kaa & KAE & kab  |  kaa & kae & KAB  |  kaa & kae & kab  ; 
assign LBA = ~lba;  //complement 
assign JAA =  HAC & haa & hab  |  hac & HAA & hab  |  hac & haa & HAB  |  HAC & HAA & HAB  ; 
assign jaa = ~JAA; //complement 
assign jba =  HAC & haa & hab  |  hac & HAA & hab  |  hac & haa & HAB  |  hac & haa & hab  ; 
assign JBA = ~jba;  //complement 
assign haa = ~HAA;  //complement 
assign HBA = ~hba;  //complement 
assign GAA =  FAA & fad & fag  |  faa & FAD & fag  |  faa & fad & FAG  |  FAA & FAD & FAG  ; 
assign gaa = ~GAA; //complement 
assign gba =  FAA & fad & fag  |  faa & FAD & fag  |  faa & fad & FAG  |  faa & fad & fag  ; 
assign GBA = ~gba;  //complement 
assign LKA =  KKA & kkc & kja  |  kka & KKC & kja  |  kka & kkc & KJA  |  KKA & KKC & KJA  ; 
assign lka = ~LKA; //complement 
assign lla =  KKA & kkc & kja  |  kka & KKC & kja  |  kka & kkc & KJA  |  kka & kkc & kja  ; 
assign LLA = ~lla;  //complement 
assign JGA =  HGA & hfa & hfb  |  hga & HFA & hfb  |  hga & hfa & HFB  |  HGA & HFA & HFB  ; 
assign jga = ~JGA; //complement 
assign jha =  HGA & hfa & hfb  |  hga & HFA & hfb  |  hga & hfa & HFB  |  hga & hfa & hfb  ; 
assign JHA = ~jha;  //complement 
assign hcc = ~HCC;  //complement 
assign HDC = ~hdc;  //complement 
assign GCE =  FBK & fbe & fch  |  fbk & FBE & fch  |  fbk & fbe & FCH  |  FBK & FBE & FCH  ; 
assign gce = ~GCE; //complement 
assign gde =  FBK & fbe & fch  |  fbk & FBE & fch  |  fbk & fbe & FCH  |  fbk & fbe & fch  ; 
assign GDE = ~gde;  //complement 
assign LUA =  KUA & kuc & kta  |  kua & KUC & kta  |  kua & kuc & KTA  |  KUA & KUC & KTA  ; 
assign lua = ~LUA; //complement 
assign lva =  KUA & kuc & kta  |  kua & KUC & kta  |  kua & kuc & KTA  |  kua & kuc & kta  ; 
assign LVA = ~lva;  //complement 
assign JKA =  HJA & hkb & hjb  |  hja & HKB & hjb  |  hja & hkb & HJB  |  HJA & HKB & HJB  ; 
assign jka = ~JKA; //complement 
assign jla =  HJA & hkb & hjb  |  hja & HKB & hjb  |  hja & hkb & HJB  |  hja & hkb & hjb  ; 
assign JLA = ~jla;  //complement 
assign hgb = ~HGB;  //complement 
assign HHB = ~hhb;  //complement 
assign GEE =  FEC & fda & fei  |  fec & FDA & fei  |  fec & fda & FEI  |  FEC & FDA & FEI  ; 
assign gee = ~GEE; //complement 
assign gfe =  FEC & fda & fei  |  fec & FDA & fei  |  fec & fda & FEI  |  fec & fda & fei  ; 
assign GFE = ~gfe;  //complement 
assign mma = ~MMA;  //complement 
assign MNA = ~mna;  //complement 
assign mmb = ~MMB;  //complement 
assign JOC =  HOD & hne & hoe  |  hod & HNE & hoe  |  hod & hne & HOE  |  HOD & HNE & HOE  ; 
assign joc = ~JOC; //complement 
assign jpc =  HOD & hne & hoe  |  hod & HNE & hoe  |  hod & hne & HOE  |  hod & hne & hoe  ; 
assign JPC = ~jpc;  //complement 
assign hie = ~HIE;  //complement 
assign HJE = ~hje;  //complement 
assign hig = ~HIG;  //complement 
assign GGE =  FGH & fgb & ffi  |  fgh & FGB & ffi  |  fgh & fgb & FFI  |  FGH & FGB & FFI  ; 
assign gge = ~GGE; //complement 
assign ghe =  FGH & fgb & ffi  |  fgh & FGB & ffi  |  fgh & fgb & FFI  |  fgh & fgb & ffi  ; 
assign GHE = ~ghe;  //complement 
assign NCA =  MCA & mcb & mba  |  mca & MCB & mba  |  mca & mcb & MBA  |  MCA & MCB & MBA  ; 
assign nca = ~NCA; //complement 
assign nda =  MCA & mcb & mba  |  mca & MCB & mba  |  mca & mcb & MBA  |  mca & mcb & mba  ; 
assign NDA = ~nda;  //complement 
assign JUB =  HUC & huf & hub  |  huc & HUF & hub  |  huc & huf & HUB  |  HUC & HUF & HUB  ; 
assign jub = ~JUB; //complement 
assign jvb =  HUC & huf & hub  |  huc & HUF & hub  |  huc & huf & HUB  |  huc & huf & hub  ; 
assign JVB = ~jvb;  //complement 
assign hmc = ~HMC;  //complement 
assign HNC = ~hnc;  //complement 
assign GIE =  FIE & fij & fhi  |  fie & FIJ & fhi  |  fie & fij & FHI  |  FIE & FIJ & FHI  ; 
assign gie = ~GIE; //complement 
assign gje =  FIE & fij & fhi  |  fie & FIJ & fhi  |  fie & fij & FHI  |  fie & fij & fhi  ; 
assign GJE = ~gje;  //complement 
assign opa = ~OPA;  //complement 
assign OQA = ~oqa;  //complement 
assign opb = ~OPB;  //complement 
assign kcc = ~KCC;  //complement 
assign KDC = ~kdc;  //complement 
assign hqb = ~HQB;  //complement 
assign HRB = ~hrb;  //complement 
assign GKF =  FKC & fjc & fki  |  fkc & FJC & fki  |  fkc & fjc & FKI  |  FKC & FJC & FKI  ; 
assign gkf = ~GKF; //complement 
assign glf =  FKC & fjc & fki  |  fkc & FJC & fki  |  fkc & fjc & FKI  |  fkc & fjc & fki  ; 
assign GLF = ~glf;  //complement 
assign ops = ~OPS;  //complement 
assign OQS = ~oqs;  //complement 
assign kkb = ~KKB;  //complement 
assign KLB = ~klb;  //complement 
assign kkd = ~KKD;  //complement 
assign hua = ~HUA;  //complement 
assign OHA = ~oha;  //complement 
assign GMG =  FMF & flf & fmj  |  fmf & FLF & fmj  |  fmf & flf & FMJ  |  FMF & FLF & FMJ  ; 
assign gmg = ~GMG; //complement 
assign gng =  FMF & flf & fmj  |  fmf & FLF & fmj  |  fmf & flf & FMJ  |  fmf & flf & fmj  ; 
assign GNG = ~gng;  //complement 
assign ksb = ~KSB;  //complement 
assign KTB = ~ktb;  //complement 
assign ksc = ~KSC;  //complement 
assign GSC =  FSH & frh & fsd  |  fsh & FRH & fsd  |  fsh & frh & FSD  |  FSH & FRH & FSD  ; 
assign gsc = ~GSC; //complement 
assign gtc =  FSH & frh & fsd  |  fsh & FRH & fsd  |  fsh & frh & FSD  |  fsh & frh & fsd  ; 
assign GTC = ~gtc;  //complement 
assign fqa = ~FQA;  //complement 
assign FRA = ~fra;  //complement 
assign faa = ~FAA;  //complement 
assign FBA = ~fba;  //complement 
assign faf = ~FAF;  //complement 
assign FBF = ~fbf;  //complement 
assign fqf = ~FQF;  //complement 
assign FRF = ~frf;  //complement 
assign fca = ~FCA;  //complement 
assign FDA = ~fda;  //complement 
assign fce = ~FCE;  //complement 
assign FDE = ~fde;  //complement 
assign fsa = ~FSA;  //complement 
assign FTA = ~fta;  //complement 
assign fea = ~FEA;  //complement 
assign FFA = ~ffa;  //complement 
assign fef = ~FEF;  //complement 
assign FFF = ~fff;  //complement 
assign fsh = ~FSH;  //complement 
assign FTH = ~fth;  //complement 
assign fsj = ~FSJ;  //complement 
assign fga = ~FGA;  //complement 
assign FHA = ~fha;  //complement 
assign fgf = ~FGF;  //complement 
assign FHF = ~fhf;  //complement 
assign fud = ~FUD;  //complement 
assign OGD = ~ogd;  //complement 
assign fia = ~FIA;  //complement 
assign FJA = ~fja;  //complement 
assign fif = ~FIF;  //complement 
assign FJF = ~fjf;  //complement 
assign fka = ~FKA;  //complement 
assign FLA = ~fla;  //complement 
assign fkf = ~FKF;  //complement 
assign FLF = ~flf;  //complement 
assign fma = ~FMA;  //complement 
assign FNA = ~fna;  //complement 
assign fmf = ~FMF;  //complement 
assign FNF = ~fnf;  //complement 
assign foa = ~FOA;  //complement 
assign FPA = ~fpa;  //complement 
assign fof = ~FOF;  //complement 
assign FPF = ~fpf;  //complement 
assign cal = ~CAL;  //complement 
assign cam = ~CAM;  //complement 
assign can = ~CAN;  //complement 
assign CGN = ~cgn;  //complement 
assign cao = ~CAO;  //complement 
assign CGO = ~cgo;  //complement 
assign cap = ~CAP;  //complement 
assign cdp = ~CDP;  //complement 
assign CGP = ~cgp;  //complement 
assign cba = ~CBA;  //complement 
assign cea = ~CEA;  //complement 
assign CHA = ~cha;  //complement 
assign cbb = ~CBB;  //complement 
assign ceb = ~CEB;  //complement 
assign CHB = ~chb;  //complement 
assign cbc = ~CBC;  //complement 
assign cec = ~CEC;  //complement 
assign CHC = ~chc;  //complement 
assign EAL =  CCP & DAL  ; 
assign eal = ~EAL;  //complement 
assign EAM =  CCO & DAM  ; 
assign eam = ~EAM;  //complement 
assign cbd = ~CBD;  //complement 
assign ced = ~CED;  //complement 
assign CHD = ~chd;  //complement 
assign LCA =  KBB & kca & kba  |  kbb & KCA & kba  |  kbb & kca & KBA  |  KBB & KCA & KBA  ; 
assign lca = ~LCA; //complement 
assign lda =  KBB & kca & kba  |  kbb & KCA & kba  |  kbb & kca & KBA  |  kbb & kca & kba  ; 
assign LDA = ~lda;  //complement 
assign JAB =  HAF & hag & had  |  haf & HAG & had  |  haf & hag & HAD  |  HAF & HAG & HAD  ; 
assign jab = ~JAB; //complement 
assign jbb =  HAF & hag & had  |  haf & HAG & had  |  haf & hag & HAD  |  haf & hag & had  ; 
assign JBB = ~jbb;  //complement 
assign hab = ~HAB;  //complement 
assign HBB = ~hbb;  //complement 
assign GAB =  FAJ & fah & fab  |  faj & FAH & fab  |  faj & fah & FAB  |  FAJ & FAH & FAB  ; 
assign gab = ~GAB; //complement 
assign gbb =  FAJ & fah & fab  |  faj & FAH & fab  |  faj & fah & FAB  |  faj & fah & fab  ; 
assign GBB = ~gbb;  //complement 
assign LKB =  KKB & kkd & kjb  |  kkb & KKD & kjb  |  kkb & kkd & KJB  |  KKB & KKD & KJB  ; 
assign lkb = ~LKB; //complement 
assign llb =  KKB & kkd & kjb  |  kkb & KKD & kjb  |  kkb & kkd & KJB  |  kkb & kkd & kjb  ; 
assign LLB = ~llb;  //complement 
assign JGB =  HGB & hgg & hfc  |  hgb & HGG & hfc  |  hgb & hgg & HFC  |  HGB & HGG & HFC  ; 
assign jgb = ~JGB; //complement 
assign jhb =  HGB & hgg & hfc  |  hgb & HGG & hfc  |  hgb & hgg & HFC  |  hgb & hgg & hfc  ; 
assign JHB = ~jhb;  //complement 
assign hcd = ~HCD;  //complement 
assign HDD = ~hdd;  //complement 
assign hce = ~HCE;  //complement 
assign GCF =  FCA & fcf & fcl  |  fca & FCF & fcl  |  fca & fcf & FCL  |  FCA & FCF & FCL  ; 
assign gcf = ~GCF; //complement 
assign gdf =  FCA & fcf & fcl  |  fca & FCF & fcl  |  fca & fcf & FCL  |  fca & fcf & fcl  ; 
assign GDF = ~gdf;  //complement 
assign maa = ~MAA;  //complement 
assign MBA = ~mba;  //complement 
assign mac = ~MAC;  //complement 
assign JKB =  HKA & hjc & hkc  |  hka & HJC & hkc  |  hka & hjc & HKC  |  HKA & HJC & HKC  ; 
assign jkb = ~JKB; //complement 
assign jlb =  HKA & hjc & hkc  |  hka & HJC & hkc  |  hka & hjc & HKC  |  hka & hjc & hkc  ; 
assign JLB = ~jlb;  //complement 
assign hgc = ~HGC;  //complement 
assign HHC = ~hhc;  //complement 
assign GEF =  FEE & fek & fdi  |  fee & FEK & fdi  |  fee & fek & FDI  |  FEE & FEK & FDI  ; 
assign gef = ~GEF; //complement 
assign gff =  FEE & fek & fdi  |  fee & FEK & fdi  |  fee & fek & FDI  |  fee & fek & fdi  ; 
assign GFF = ~gff;  //complement 
assign moa = ~MOA;  //complement 
assign MPA = ~mpa;  //complement 
assign mob = ~MOB;  //complement 
assign JQA =  HQB & hpa & hqa  |  hqb & HPA & hqa  |  hqb & hpa & HQA  |  HQB & HPA & HQA  ; 
assign jqa = ~JQA; //complement 
assign jra =  HQB & hpa & hqa  |  hqb & HPA & hqa  |  hqb & hpa & HQA  |  hqb & hpa & hqa  ; 
assign JRA = ~jra;  //complement 
assign hka = ~HKA;  //complement 
assign HLA = ~hla;  //complement 
assign GGF =  FFE & ffc & ffk  |  ffe & FFC & ffk  |  ffe & ffc & FFK  |  FFE & FFC & FFK  ; 
assign ggf = ~GGF; //complement 
assign ghf =  FFE & ffc & ffk  |  ffe & FFC & ffk  |  ffe & ffc & FFK  |  ffe & ffc & ffk  ; 
assign GHF = ~ghf;  //complement 
assign NEA =  MDA & mea & meb  |  mda & MEA & meb  |  mda & mea & MEB  |  MDA & MEA & MEB  ; 
assign nea = ~NEA; //complement 
assign nfa =  MDA & mea & meb  |  mda & MEA & meb  |  mda & mea & MEB  |  mda & mea & meb  ; 
assign NFA = ~nfa;  //complement 
assign JUC =  HUD & htc & htd  |  hud & HTC & htd  |  hud & htc & HTD  |  HUD & HTC & HTD  ; 
assign juc = ~JUC; //complement 
assign jvc =  HUD & htc & htd  |  hud & HTC & htd  |  hud & htc & HTD  |  hud & htc & htd  ; 
assign JVC = ~jvc;  //complement 
assign hmd = ~HMD;  //complement 
assign HND = ~hnd;  //complement 
assign GIF =  FIC & fhc & fii  |  fic & FHC & fii  |  fic & fhc & FII  |  FIC & FHC & FII  ; 
assign gif = ~GIF; //complement 
assign gjf =  FIC & fhc & fii  |  fic & FHC & fii  |  fic & fhc & FII  |  fic & fhc & fii  ; 
assign GJF = ~gjf;  //complement 
assign opc = ~OPC;  //complement 
assign OQC = ~oqc;  //complement 
assign opd = ~OPD;  //complement 
assign kea = ~KEA;  //complement 
assign KFA = ~kfa;  //complement 
assign hqc = ~HQC;  //complement 
assign HRC = ~hrc;  //complement 
assign GKG =  FJK & fji & fjf  |  fjk & FJI & fjf  |  fjk & fji & FJF  |  FJK & FJI & FJF  ; 
assign gkg = ~GKG; //complement 
assign glg =  FJK & fji & fjf  |  fjk & FJI & fjf  |  fjk & fji & FJF  |  fjk & fji & fjf  ; 
assign GLG = ~glg;  //complement 
assign opu = ~OPU;  //complement 
assign OQU = ~oqu;  //complement 
assign kma = ~KMA;  //complement 
assign KNA = ~kna;  //complement 
assign kmc = ~KMC;  //complement 
assign hub = ~HUB;  //complement 
assign OHB = ~ohb;  //complement 
assign GOA =  FOA & fna & fog  |  foa & FNA & fog  |  foa & fna & FOG  |  FOA & FNA & FOG  ; 
assign goa = ~GOA; //complement 
assign gpa =  FOA & fna & fog  |  foa & FNA & fog  |  foa & fna & FOG  |  foa & fna & fog  ; 
assign GPA = ~gpa;  //complement 
assign kua = ~KUA;  //complement 
assign OKA = ~oka;  //complement 
assign GSE =  FSE & fre & fsi  |  fse & FRE & fsi  |  fse & fre & FSI  |  FSE & FRE & FSI  ; 
assign gse = ~GSE; //complement 
assign gte =  FSE & fre & fsi  |  fse & FRE & fsi  |  fse & fre & FSI  |  fse & fre & fsi  ; 
assign GTE = ~gte;  //complement 
assign GQB =  FPG & fqd & fpd  |  fpg & FQD & fpd  |  fpg & fqd & FPD  |  FPG & FQD & FPD  ; 
assign gqb = ~GQB; //complement 
assign grb =  FPG & fqd & fpd  |  fpg & FQD & fpd  |  fpg & fqd & FPD  |  fpg & fqd & fpd  ; 
assign GRB = ~grb;  //complement 
assign fqb = ~FQB;  //complement 
assign FRB = ~frb;  //complement 
assign fab = ~FAB;  //complement 
assign FBB = ~fbb;  //complement 
assign fag = ~FAG;  //complement 
assign FBG = ~fbg;  //complement 
assign fqg = ~FQG;  //complement 
assign FRG = ~frg;  //complement 
assign ECM =  CCP & DAM  ; 
assign ecm = ~ECM;  //complement 
assign fcb = ~FCB;  //complement 
assign FDB = ~fdb;  //complement 
assign fcf = ~FCF;  //complement 
assign FDF = ~fdf;  //complement 
assign fsb = ~FSB;  //complement 
assign FTB = ~ftb;  //complement 
assign feb = ~FEB;  //complement 
assign FFB = ~ffb;  //complement 
assign feg = ~FEG;  //complement 
assign FFG = ~ffg;  //complement 
assign fsi = ~FSI;  //complement 
assign FTI = ~fti;  //complement 
assign fsk = ~FSK;  //complement 
assign fgb = ~FGB;  //complement 
assign FHB = ~fhb;  //complement 
assign fgg = ~FGG;  //complement 
assign FHG = ~fhg;  //complement 
assign fue = ~FUE;  //complement 
assign OGE = ~oge;  //complement 
assign fib = ~FIB;  //complement 
assign FJB = ~fjb;  //complement 
assign fig = ~FIG;  //complement 
assign FJG = ~fjg;  //complement 
assign fkb = ~FKB;  //complement 
assign FLB = ~flb;  //complement 
assign fkg = ~FKG;  //complement 
assign FLG = ~flg;  //complement 
assign fmb = ~FMB;  //complement 
assign FNB = ~fnb;  //complement 
assign fmg = ~FMG;  //complement 
assign FNG = ~fng;  //complement 
assign GSD =  FSB & fsj & fsg  |  fsb & FSJ & fsg  |  fsb & fsj & FSG  |  FSB & FSJ & FSG  ; 
assign gsd = ~GSD; //complement 
assign gtd =  FSB & fsj & fsg  |  fsb & FSJ & fsg  |  fsb & fsj & FSG  |  fsb & fsj & fsg  ; 
assign GTD = ~gtd;  //complement 
assign fob = ~FOB;  //complement 
assign FPB = ~fpb;  //complement 
assign fog = ~FOG;  //complement 
assign FPG = ~fpg;  //complement 
assign cbe = ~CBE;  //complement 
assign cee = ~CEE;  //complement 
assign CHE = ~che;  //complement 
assign CHL = ~chl;  //complement 
assign cbf = ~CBF;  //complement 
assign cef = ~CEF;  //complement 
assign CHF = ~chf;  //complement 
assign CKL = ~ckl;  //complement 
assign cbg = ~CBG;  //complement 
assign ceg = ~CEG;  //complement 
assign CHG = ~chg;  //complement 
assign CHH = ~chh;  //complement 
assign cbh = ~CBH;  //complement 
assign ceh = ~CEH;  //complement 
assign taa = ~TAA;  //complement 
assign tab = ~TAB;  //complement 
assign cbi = ~CBI;  //complement 
assign cei = ~CEI;  //complement 
assign qic = ~QIC;  //complement 
assign qid = ~QID;  //complement 
assign qie = ~QIE;  //complement 
assign qif = ~QIF;  //complement 
assign qig = ~QIG;  //complement 
assign qih = ~QIH;  //complement 
assign CHI = ~chi;  //complement 
assign CKI = ~cki;  //complement 
assign CHJ = ~chj;  //complement 
assign CKJ = ~ckj;  //complement 
assign cbj = ~CBJ;  //complement 
assign cej = ~CEJ;  //complement 
assign cbk = ~CBK;  //complement 
assign cek = ~CEK;  //complement 
assign CHK = ~chk;  //complement 
assign CKK = ~ckk;  //complement 
assign GSB =  FSA & frb & fsf  |  fsa & FRB & fsf  |  fsa & frb & FSF  |  FSA & FRB & FSF  ; 
assign gsb = ~GSB; //complement 
assign gtb =  FSA & frb & fsf  |  fsa & FRB & fsf  |  fsa & frb & FSF  |  fsa & frb & fsf  ; 
assign GTB = ~gtb;  //complement 
assign cbl = ~CBL;  //complement 
assign cel = ~CEL;  //complement 
assign LCB =  KBC & kbd & kcb  |  kbc & KBD & kcb  |  kbc & kbd & KCB  |  KBC & KBD & KCB  ; 
assign lcb = ~LCB; //complement 
assign ldb =  KBC & kbd & kcb  |  kbc & KBD & kcb  |  kbc & kbd & KCB  |  kbc & kbd & kcb  ; 
assign LDB = ~ldb;  //complement 
assign JCA =  HBA & hca & hbb  |  hba & HCA & hbb  |  hba & hca & HBB  |  HBA & HCA & HBB  ; 
assign jca = ~JCA; //complement 
assign jda =  HBA & hca & hbb  |  hba & HCA & hbb  |  hba & hca & HBB  |  hba & hca & hbb  ; 
assign JDA = ~jda;  //complement 
assign hac = ~HAC;  //complement 
assign HBC = ~hbc;  //complement 
assign GAC =  FAK & fae & fac  |  fak & FAE & fac  |  fak & fae & FAC  |  FAK & FAE & FAC  ; 
assign gac = ~GAC; //complement 
assign gbc =  FAK & fae & fac  |  fak & FAE & fac  |  fak & fae & FAC  |  fak & fae & fac  ; 
assign GBC = ~gbc;  //complement 
assign LMA =  KMB & kma & kla  |  kmb & KMA & kla  |  kmb & kma & KLA  |  KMB & KMA & KLA  ; 
assign lma = ~LMA; //complement 
assign lna =  KMB & kma & kla  |  kmb & KMA & kla  |  kmb & kma & KLA  |  kmb & kma & kla  ; 
assign LNA = ~lna;  //complement 
assign JGC =  HGC & hgf & hfd  |  hgc & HGF & hfd  |  hgc & hgf & HFD  |  HGC & HGF & HFD  ; 
assign jgc = ~JGC; //complement 
assign jhc =  HGC & hgf & hfd  |  hgc & HGF & hfd  |  hgc & hgf & HFD  |  hgc & hgf & hfd  ; 
assign JHC = ~jhc;  //complement 
assign hea = ~HEA;  //complement 
assign HFA = ~hfa;  //complement 
assign GCG =  FBF & fbl & fbc  |  fbf & FBL & fbc  |  fbf & fbl & FBC  |  FBF & FBL & FBC  ; 
assign gcg = ~GCG; //complement 
assign gdg =  FBF & fbl & fbc  |  fbf & FBL & fbc  |  fbf & fbl & FBC  |  fbf & fbl & fbc  ; 
assign GDG = ~gdg;  //complement 
assign mab = ~MAB;  //complement 
assign MBB = ~mbb;  //complement 
assign mad = ~MAD;  //complement 
assign JKC =  HKE & hje & hkd  |  hke & HJE & hkd  |  hke & hje & HKD  |  HKE & HJE & HKD  ; 
assign jkc = ~JKC; //complement 
assign jlc =  HKE & hje & hkd  |  hke & HJE & hkd  |  hke & hje & HKD  |  hke & hje & hkd  ; 
assign JLC = ~jlc;  //complement 
assign hgd = ~HGD;  //complement 
assign HHD = ~hhd;  //complement 
assign hgf = ~HGF;  //complement 
assign GEG =  FDL & fdh & fdf  |  fdl & FDH & fdf  |  fdl & fdh & FDF  |  FDL & FDH & FDF  ; 
assign geg = ~GEG; //complement 
assign gfg =  FDL & fdh & fdf  |  fdl & FDH & fdf  |  fdl & fdh & FDF  |  fdl & fdh & fdf  ; 
assign GFG = ~gfg;  //complement 
assign JQB =  HQC & hpc & hpb  |  hqc & HPC & hpb  |  hqc & hpc & HPB  |  HQC & HPC & HPB  ; 
assign jqb = ~JQB; //complement 
assign jrb =  HQC & hpc & hpb  |  hqc & HPC & hpb  |  hqc & hpc & HPB  |  hqc & hpc & hpb  ; 
assign JRB = ~jrb;  //complement 
assign hkb = ~HKB;  //complement 
assign HLB = ~hlb;  //complement 
assign GGG =  FGC & fff & fgi  |  fgc & FFF & fgi  |  fgc & fff & FGI  |  FGC & FFF & FGI  ; 
assign ggg = ~GGG; //complement 
assign ghg =  FGC & fff & fgi  |  fgc & FFF & fgi  |  fgc & fff & FGI  |  fgc & fff & fgi  ; 
assign GHG = ~ghg;  //complement 
assign NGA =  MFA & mga & mgc  |  mfa & MGA & mgc  |  mfa & mga & MGC  |  MFA & MGA & MGC  ; 
assign nga = ~NGA; //complement 
assign nha =  MFA & mga & mgc  |  mfa & MGA & mgc  |  mfa & mga & MGC  |  mfa & mga & mgc  ; 
assign NHA = ~nha;  //complement 
assign kaa = ~KAA;  //complement 
assign KBA = ~kba;  //complement 
assign hme = ~HME;  //complement 
assign HNE = ~hne;  //complement 
assign hmf = ~HMF;  //complement 
assign GIG =  FIK & fhk & fif  |  fik & FHK & fif  |  fik & fhk & FIF  |  FIK & FHK & FIF  ; 
assign gig = ~GIG; //complement 
assign gjg =  FIK & fhk & fif  |  fik & FHK & fif  |  fik & fhk & FIF  |  fik & fhk & fif  ; 
assign GJG = ~gjg;  //complement 
assign opg = ~OPG;  //complement 
assign OQG = ~oqg;  //complement 
assign keb = ~KEB;  //complement 
assign KFB = ~kfb;  //complement 
assign kec = ~KEC;  //complement 
assign hqd = ~HQD;  //complement 
assign HRD = ~hrd;  //complement 
assign GMA =  FMA & fld & fmg  |  fma & FLD & fmg  |  fma & fld & FMG  |  FMA & FLD & FMG  ; 
assign gma = ~GMA; //complement 
assign gna =  FMA & fld & fmg  |  fma & FLD & fmg  |  fma & fld & FMG  |  fma & fld & fmg  ; 
assign GNA = ~gna;  //complement 
assign kmb = ~KMB;  //complement 
assign KNB = ~knb;  //complement 
assign kmd = ~KMD;  //complement 
assign huc = ~HUC;  //complement 
assign OHC = ~ohc;  //complement 
assign hue = ~HUE;  //complement 
assign GOB =  FOD & fng & fok  |  fod & FNG & fok  |  fod & fng & FOK  |  FOD & FNG & FOK  ; 
assign gob = ~GOB; //complement 
assign gpb =  FOD & fng & fok  |  fod & FNG & fok  |  fod & fng & FOK  |  fod & fng & fok  ; 
assign GPB = ~gpb;  //complement 
assign kub = ~KUB;  //complement 
assign OKB = ~okb;  //complement 
assign kuc = ~KUC;  //complement 
assign GSF =  FSC & frc & fsk  |  fsc & FRC & fsk  |  fsc & frc & FSK  |  FSC & FRC & FSK  ; 
assign gsf = ~GSF; //complement 
assign gtf =  FSC & frc & fsk  |  fsc & FRC & fsk  |  fsc & frc & FSK  |  fsc & frc & fsk  ; 
assign GTF = ~gtf;  //complement 
assign GQC =  FQH & fqb & fpi  |  fqh & FQB & fpi  |  fqh & fqb & FPI  |  FQH & FQB & FPI  ; 
assign gqc = ~GQC; //complement 
assign grc =  FQH & fqb & fpi  |  fqh & FQB & fpi  |  fqh & fqb & FPI  |  fqh & fqb & fpi  ; 
assign GRC = ~grc;  //complement 
assign fac = ~FAC;  //complement 
assign FBC = ~fbc;  //complement 
assign fah = ~FAH;  //complement 
assign FBH = ~fbh;  //complement 
assign fcg = ~FCG;  //complement 
assign FDG = ~fdg;  //complement 
assign cbm = ~CBM;  //complement 
assign cem = ~CEM;  //complement 
assign CHM = ~chm;  //complement 
assign CKM = ~ckm;  //complement 
assign cbn = ~CBN;  //complement 
assign cen = ~CEN;  //complement 
assign CHN = ~chn;  //complement 
assign CKN = ~ckn;  //complement 
assign cbo = ~CBO;  //complement 
assign ceo = ~CEO;  //complement 
assign CHO = ~cho;  //complement 
assign CKO = ~cko;  //complement 
assign cbp = ~CBP;  //complement 
assign cep = ~CEP;  //complement 
assign CHP = ~chp;  //complement 
assign CKP = ~ckp;  //complement 
assign cca = ~CCA;  //complement 
assign cfa = ~CFA;  //complement 
assign CIA = ~cia;  //complement 
assign CLA = ~cla;  //complement 
assign ccb = ~CCB;  //complement 
assign cfb = ~CFB;  //complement 
assign CIB = ~cib;  //complement 
assign CLB = ~clb;  //complement 
assign ccc = ~CCC;  //complement 
assign cfc = ~CFC;  //complement 
assign CIC = ~cic;  //complement 
assign CLC = ~clc;  //complement 
assign qja = ~QJA;  //complement 
assign qjb = ~QJB;  //complement 
assign qjc = ~QJC;  //complement 
assign ccd = ~CCD;  //complement 
assign cfd = ~CFD;  //complement 
assign CID = ~cid;  //complement 
assign CLD = ~cld;  //complement 
assign LEA =  KEA & kdb & kda  |  kea & KDB & kda  |  kea & kdb & KDA  |  KEA & KDB & KDA  ; 
assign lea = ~LEA; //complement 
assign lfa =  KEA & kdb & kda  |  kea & KDB & kda  |  kea & kdb & KDA  |  kea & kdb & kda  ; 
assign LFA = ~lfa;  //complement 
assign JCB =  HBD & hcb & hbc  |  hbd & HCB & hbc  |  hbd & hcb & HBC  |  HBD & HCB & HBC  ; 
assign jcb = ~JCB; //complement 
assign jdb =  HBD & hcb & hbc  |  hbd & HCB & hbc  |  hbd & hcb & HBC  |  hbd & hcb & hbc  ; 
assign JDB = ~jdb;  //complement 
assign had = ~HAD;  //complement 
assign HBD = ~hbd;  //complement 
assign GAD =  FAL & fai & faf  |  fal & FAI & faf  |  fal & fai & FAF  |  FAL & FAI & FAF  ; 
assign gad = ~GAD; //complement 
assign gbd =  FAL & fai & faf  |  fal & FAI & faf  |  fal & fai & FAF  |  fal & fai & faf  ; 
assign GBD = ~gbd;  //complement 
assign LMB =  KLB & kmc & kmd  |  klb & KMC & kmd  |  klb & kmc & KMD  |  KLB & KMC & KMD  ; 
assign lmb = ~LMB; //complement 
assign lnb =  KLB & kmc & kmd  |  klb & KMC & kmd  |  klb & kmc & KMD  |  klb & kmc & kmd  ; 
assign LNB = ~lnb;  //complement 
assign JGD =  HFE & hgd & hge  |  hfe & HGD & hge  |  hfe & hgd & HGE  |  HFE & HGD & HGE  ; 
assign jgd = ~JGD; //complement 
assign jhd =  HFE & hgd & hge  |  hfe & HGD & hge  |  hfe & hgd & HGE  |  hfe & hgd & hge  ; 
assign JHD = ~jhd;  //complement 
assign heb = ~HEB;  //complement 
assign HFB = ~hfb;  //complement 
assign GCH =  FCG & fci & fbi  |  fcg & FCI & fbi  |  fcg & fci & FBI  |  FCG & FCI & FBI  ; 
assign gch = ~GCH; //complement 
assign gdh =  FCG & fci & fbi  |  fcg & FCI & fbi  |  fcg & fci & FBI  |  fcg & fci & fbi  ; 
assign GDH = ~gdh;  //complement 
assign mca = ~MCA;  //complement 
assign MDA = ~mda;  //complement 
assign mcb = ~MCB;  //complement 
assign JMA =  HMA & hla & hlb  |  hma & HLA & hlb  |  hma & hla & HLB  |  HMA & HLA & HLB  ; 
assign jma = ~JMA; //complement 
assign jna =  HMA & hla & hlb  |  hma & HLA & hlb  |  hma & hla & HLB  |  hma & hla & hlb  ; 
assign JNA = ~jna;  //complement 
assign hge = ~HGE;  //complement 
assign HHE = ~hhe;  //complement 
assign hgg = ~HGG;  //complement 
assign GEH =  FEF & fel & fdc  |  fef & FEL & fdc  |  fef & fel & FDC  |  FEF & FEL & FDC  ; 
assign geh = ~GEH; //complement 
assign gfh =  FEF & fel & fdc  |  fef & FEL & fdc  |  fef & fel & FDC  |  fef & fel & fdc  ; 
assign GFH = ~gfh;  //complement 
assign mqa = ~MQA;  //complement 
assign MRA = ~mra;  //complement 
assign mqb = ~MQB;  //complement 
assign JQC =  HQE & hpd & hqd  |  hqe & HPD & hqd  |  hqe & hpd & HQD  |  HQE & HPD & HQD  ; 
assign jqc = ~JQC; //complement 
assign jrc =  HQE & hpd & hqd  |  hqe & HPD & hqd  |  hqe & hpd & HQD  |  hqe & hpd & hqd  ; 
assign JRC = ~jrc;  //complement 
assign hkc = ~HKC;  //complement 
assign HLC = ~hlc;  //complement 
assign GGH =  FGK & ffl & fgf  |  fgk & FFL & fgf  |  fgk & ffl & FGF  |  FGK & FFL & FGF  ; 
assign ggh = ~GGH; //complement 
assign ghh =  FGK & ffl & fgf  |  fgk & FFL & fgf  |  fgk & ffl & FGF  |  fgk & ffl & fgf  ; 
assign GHH = ~ghh;  //complement 
assign mgc = ~MGC;  //complement 
assign mcc = ~MCC;  //complement 
assign ope = ~OPE;  //complement 
assign opf = ~OPF;  //complement 
assign kab = ~KAB;  //complement 
assign KBB = ~kbb;  //complement 
assign hoa = ~HOA;  //complement 
assign HPA = ~hpa;  //complement 
assign GKA =  FJA & fjg & fkd  |  fja & FJG & fkd  |  fja & fjg & FKD  |  FJA & FJG & FKD  ; 
assign gka = ~GKA; //complement 
assign gla =  FJA & fjg & fkd  |  fja & FJG & fkd  |  fja & fjg & FKD  |  fja & fjg & fkd  ; 
assign GLA = ~gla;  //complement 
assign opi = ~OPI;  //complement 
assign OQI = ~oqi;  //complement 
assign kga = ~KGA;  //complement 
assign KHA = ~kha;  //complement 
assign hqe = ~HQE;  //complement 
assign HRE = ~hre;  //complement 
assign GMB =  FLA & flg & fle  |  fla & FLG & fle  |  fla & flg & FLE  |  FLA & FLG & FLE  ; 
assign gmb = ~GMB; //complement 
assign gnb =  FLA & flg & fle  |  fla & FLG & fle  |  fla & flg & FLE  |  fla & flg & fle  ; 
assign GNB = ~gnb;  //complement 
assign koa = ~KOA;  //complement 
assign KPA = ~kpa;  //complement 
assign koc = ~KOC;  //complement 
assign hud = ~HUD;  //complement 
assign OHD = ~ohd;  //complement 
assign huf = ~HUF;  //complement 
assign GOC =  FNE & fnd & fni  |  fne & FND & fni  |  fne & fnd & FNI  |  FNE & FND & FNI  ; 
assign goc = ~GOC; //complement 
assign gpc =  FNE & fnd & fni  |  fne & FND & fni  |  fne & fnd & FNI  |  fne & fnd & fni  ; 
assign GPC = ~gpc;  //complement 
assign GSG =  FRJ & fri & frf  |  frj & FRI & frf  |  frj & fri & FRF  |  FRJ & FRI & FRF  ; 
assign gsg = ~GSG; //complement 
assign gtg =  FRJ & fri & frf  |  frj & FRI & frf  |  frj & fri & FRF  |  frj & fri & frf  ; 
assign GTG = ~gtg;  //complement 
assign GQD =  FQI & fph & fqe  |  fqi & FPH & fqe  |  fqi & fph & FQE  |  FQI & FPH & FQE  ; 
assign gqd = ~GQD; //complement 
assign grd =  FQI & fph & fqe  |  fqi & FPH & fqe  |  fqi & fph & FQE  |  fqi & fph & fqe  ; 
assign GRD = ~grd;  //complement 
assign fqc = ~FQC;  //complement 
assign FRC = ~frc;  //complement 
assign fad = ~FAD;  //complement 
assign FBD = ~fbd;  //complement 
assign fai = ~FAI;  //complement 
assign FBI = ~fbi;  //complement 
assign fqh = ~FQH;  //complement 
assign FRH = ~frh;  //complement 
assign fcc = ~FCC;  //complement 
assign FDC = ~fdc;  //complement 
assign fch = ~FCH;  //complement 
assign FDH = ~fdh;  //complement 
assign fsc = ~FSC;  //complement 
assign FTC = ~ftc;  //complement 
assign fec = ~FEC;  //complement 
assign FFC = ~ffc;  //complement 
assign feh = ~FEH;  //complement 
assign FFH = ~ffh;  //complement 
assign fua = ~FUA;  //complement 
assign OGA = ~oga;  //complement 
assign fgc = ~FGC;  //complement 
assign FHC = ~fhc;  //complement 
assign fgh = ~FGH;  //complement 
assign FHH = ~fhh;  //complement 
assign fuf = ~FUF;  //complement 
assign OGF = ~ogf;  //complement 
assign fic = ~FIC;  //complement 
assign FJC = ~fjc;  //complement 
assign fih = ~FIH;  //complement 
assign FJH = ~fjh;  //complement 
assign fkc = ~FKC;  //complement 
assign FLC = ~flc;  //complement 
assign fkh = ~FKH;  //complement 
assign FLH = ~flh;  //complement 
assign fmc = ~FMC;  //complement 
assign FNC = ~fnc;  //complement 
assign fmh = ~FMH;  //complement 
assign FNH = ~fnh;  //complement 
assign foc = ~FOC;  //complement 
assign FPC = ~fpc;  //complement 
assign foh = ~FOH;  //complement 
assign FPH = ~fph;  //complement 
assign cce = ~CCE;  //complement 
assign cfe = ~CFE;  //complement 
assign CIE = ~cie;  //complement 
assign ccf = ~CCF;  //complement 
assign cff = ~CFF;  //complement 
assign CIF = ~cif;  //complement 
assign ccg = ~CCG;  //complement 
assign cfg = ~CFG;  //complement 
assign CIG = ~cig;  //complement 
assign cch = ~CCH;  //complement 
assign cfh = ~CFH;  //complement 
assign CIH = ~cih;  //complement 
assign cci = ~CCI;  //complement 
assign cfi = ~CFI;  //complement 
assign CII = ~cii;  //complement 
assign ccj = ~CCJ;  //complement 
assign cfj = ~CFJ;  //complement 
assign CIJ = ~cij;  //complement 
assign ERW = DIO & CHE ; 
assign erw = ~ERW ; //complement 
assign ETW = DIO & CHF ; 
assign etw = ~ETW ;  //complement 
assign EVW = DIO & CHG ; 
assign evw = ~EVW ;  //complement 
assign cck = ~CCK;  //complement 
assign cfk = ~CFK;  //complement 
assign CIK = ~cik;  //complement 
assign ERX = DIP & CHD ; 
assign erx = ~ERX ; //complement 
assign ETX = DIP & CHE ; 
assign etx = ~ETX ;  //complement 
assign EVX = DIP & CHF ; 
assign evx = ~EVX ;  //complement 
assign ccl = ~CCL;  //complement 
assign cfl = ~CFL;  //complement 
assign CIL = ~cil;  //complement 
assign LEB =  KEB & kec & kdc  |  keb & KEC & kdc  |  keb & kec & KDC  |  KEB & KEC & KDC  ; 
assign leb = ~LEB; //complement 
assign lfb =  KEB & kec & kdc  |  keb & KEC & kdc  |  keb & kec & KDC  |  keb & kec & kdc  ; 
assign LFB = ~lfb;  //complement 
assign JCC =  HCD & hce & hbf  |  hcd & HCE & hbf  |  hcd & hce & HBF  |  HCD & HCE & HBF  ; 
assign jcc = ~JCC; //complement 
assign jdc =  HCD & hce & hbf  |  hcd & HCE & hbf  |  hcd & hce & HBF  |  hcd & hce & hbf  ; 
assign JDC = ~jdc;  //complement 
assign hae = ~HAE;  //complement 
assign HBE = ~hbe;  //complement 
assign GCA =  FBG & fba & fbj  |  fbg & FBA & fbj  |  fbg & fba & FBJ  |  FBG & FBA & FBJ  ; 
assign gca = ~GCA; //complement 
assign gda =  FBG & fba & fbj  |  fbg & FBA & fbj  |  fbg & fba & FBJ  |  fbg & fba & fbj  ; 
assign GDA = ~gda;  //complement 
assign LOA =  KNA & kod & knb  |  kna & KOD & knb  |  kna & kod & KNB  |  KNA & KOD & KNB  ; 
assign loa = ~LOA; //complement 
assign lpa =  KNA & kod & knb  |  kna & KOD & knb  |  kna & kod & KNB  |  kna & kod & knb  ; 
assign LPA = ~lpa;  //complement 
assign JIA =  HIA & hha & hib  |  hia & HHA & hib  |  hia & hha & HIB  |  HIA & HHA & HIB  ; 
assign jia = ~JIA; //complement 
assign jja =  HIA & hha & hib  |  hia & HHA & hib  |  hia & hha & HIB  |  hia & hha & hib  ; 
assign JJA = ~jja;  //complement 
assign hec = ~HEC;  //complement 
assign HFC = ~hfc;  //complement 
assign GEA =  FEA & feg & fdj  |  fea & FEG & fdj  |  fea & feg & FDJ  |  FEA & FEG & FDJ  ; 
assign gea = ~GEA; //complement 
assign gfa =  FEA & feg & fdj  |  fea & FEG & fdj  |  fea & feg & FDJ  |  fea & feg & fdj  ; 
assign GFA = ~gfa;  //complement 
assign mea = ~MEA;  //complement 
assign MFA = ~mfa;  //complement 
assign meb = ~MEB;  //complement 
assign JMB =  HMB & hmf & hmd  |  hmb & HMF & hmd  |  hmb & hmf & HMD  |  HMB & HMF & HMD  ; 
assign jmb = ~JMB; //complement 
assign jnb =  HMB & hmf & hmd  |  hmb & HMF & hmd  |  hmb & hmf & HMD  |  hmb & hmf & hmd  ; 
assign JNB = ~jnb;  //complement 
assign hia = ~HIA;  //complement 
assign HJA = ~hja;  //complement 
assign GGA =  FGA & ffa & fgg  |  fga & FFA & fgg  |  fga & ffa & FGG  |  FGA & FFA & FGG  ; 
assign gga = ~GGA; //complement 
assign gha =  FGA & ffa & fgg  |  fga & FFA & fgg  |  fga & ffa & FGG  |  fga & ffa & fgg  ; 
assign GHA = ~gha;  //complement 
assign msa = ~MSA;  //complement 
assign MTA = ~mta;  //complement 
assign msb = ~MSB;  //complement 
assign JSA =  HSA & hra & hrb  |  hsa & HRA & hrb  |  hsa & hra & HRB  |  HSA & HRA & HRB  ; 
assign jsa = ~JSA; //complement 
assign jta =  HSA & hra & hrb  |  hsa & HRA & hrb  |  hsa & hra & HRB  |  hsa & hra & hrb  ; 
assign JTA = ~jta;  //complement 
assign hkd = ~HKD;  //complement 
assign HLD = ~hld;  //complement 
assign GIA =  FIA & fig & fhg  |  fia & FIG & fhg  |  fia & fig & FHG  |  FIA & FIG & FHG  ; 
assign gia = ~GIA; //complement 
assign gja =  FIA & fig & fhg  |  fia & FIG & fhg  |  fia & fig & FHG  |  fia & fig & fhg  ; 
assign GJA = ~gja;  //complement 
assign omb = ~OMB;  //complement 
assign kac = ~KAC;  //complement 
assign KBC = ~kbc;  //complement 
assign hob = ~HOB;  //complement 
assign HPB = ~hpb;  //complement 
assign GKB =  FKA & fjb & fkg  |  fka & FJB & fkg  |  fka & fjb & FKG  |  FKA & FJB & FKG  ; 
assign gkb = ~GKB; //complement 
assign glb =  FKA & fjb & fkg  |  fka & FJB & fkg  |  fka & fjb & FKG  |  fka & fjb & fkg  ; 
assign GLB = ~glb;  //complement 
assign opk = ~OPK;  //complement 
assign OQK = ~oqk;  //complement 
assign kgb = ~KGB;  //complement 
assign KHB = ~khb;  //complement 
assign kgc = ~KGC;  //complement 
assign hsa = ~HSA;  //complement 
assign HTA = ~hta;  //complement 
assign GMC =  FME & fmi & fmd  |  fme & FMI & fmd  |  fme & fmi & FMD  |  FME & FMI & FMD  ; 
assign gmc = ~GMC; //complement 
assign gnc =  FME & fmi & fmd  |  fme & FMI & fmd  |  fme & fmi & FMD  |  fme & fmi & fmd  ; 
assign GNC = ~gnc;  //complement 
assign kob = ~KOB;  //complement 
assign KPB = ~kpb;  //complement 
assign kod = ~KOD;  //complement 
assign GOD =  FOE & foi & fnh  |  foe & FOI & fnh  |  foe & foi & FNH  |  FOE & FOI & FNH  ; 
assign god = ~GOD; //complement 
assign gpd =  FOE & foi & fnh  |  foe & FOI & fnh  |  foe & foi & FNH  |  foe & foi & fnh  ; 
assign GPD = ~gpd;  //complement 
assign GUA =  FUF & fuj & fua  |  fuf & FUJ & fua  |  fuf & fuj & FUA  |  FUF & FUJ & FUA  ; 
assign gua = ~GUA; //complement 
assign gva =  FUF & fuj & fua  |  fuf & FUJ & fua  |  fuf & fuj & FUA  |  fuf & fuj & fua  ; 
assign GVA = ~gva;  //complement 
assign GQE =  FQC & fpc & fpj  |  fqc & FPC & fpj  |  fqc & fpc & FPJ  |  FQC & FPC & FPJ  ; 
assign gqe = ~GQE; //complement 
assign gre =  FQC & fpc & fpj  |  fqc & FPC & fpj  |  fqc & fpc & FPJ  |  fqc & fpc & fpj  ; 
assign GRE = ~gre;  //complement 
assign fqd = ~FQD;  //complement 
assign FRD = ~frd;  //complement 
assign fae = ~FAE;  //complement 
assign FBE = ~fbe;  //complement 
assign faj = ~FAJ;  //complement 
assign FBJ = ~fbj;  //complement 
assign fam = ~FAM;  //complement 
assign fqi = ~FQI;  //complement 
assign FRI = ~fri;  //complement 
assign fcd = ~FCD;  //complement 
assign FDD = ~fdd;  //complement 
assign fci = ~FCI;  //complement 
assign FDI = ~fdi;  //complement 
assign fsd = ~FSD;  //complement 
assign FTD = ~ftd;  //complement 
assign fed = ~FED;  //complement 
assign FFD = ~ffd;  //complement 
assign fei = ~FEI;  //complement 
assign FFI = ~ffi;  //complement 
assign fub = ~FUB;  //complement 
assign OGB = ~ogb;  //complement 
assign fgd = ~FGD;  //complement 
assign FHD = ~fhd;  //complement 
assign fgi = ~FGI;  //complement 
assign FHI = ~fhi;  //complement 
assign fug = ~FUG;  //complement 
assign OGG = ~ogg;  //complement 
assign fid = ~FID;  //complement 
assign FJD = ~fjd;  //complement 
assign fii = ~FII;  //complement 
assign FJI = ~fji;  //complement 
assign fkd = ~FKD;  //complement 
assign FLD = ~fld;  //complement 
assign fki = ~FKI;  //complement 
assign FLI = ~fli;  //complement 
assign fmd = ~FMD;  //complement 
assign FND = ~fnd;  //complement 
assign fmi = ~FMI;  //complement 
assign FNI = ~fni;  //complement 
assign fmk = ~FMK;  //complement 
assign fod = ~FOD;  //complement 
assign FPD = ~fpd;  //complement 
assign foi = ~FOI;  //complement 
assign FPI = ~fpi;  //complement 
assign ccm = ~CCM;  //complement 
assign cfm = ~CFM;  //complement 
assign CIM = ~cim;  //complement 
assign EBD = DBL & CBP ; 
assign ebd = ~EBD ; //complement 
assign EDD = DBL & CCA ; 
assign edd = ~EDD ;  //complement 
assign EFD = DBL & CCB ; 
assign efd = ~EFD ;  //complement 
assign EHD = DBL & CCC; 
assign ehd = ~EHD; 
assign ccn = ~CCN;  //complement 
assign cfn = ~CFN;  //complement 
assign CIN = ~cin;  //complement 
assign cco = ~CCO;  //complement 
assign cfo = ~CFO;  //complement 
assign CIO = ~cio;  //complement 
assign ccp = ~CCP;  //complement 
assign cfp = ~CFP;  //complement 
assign CIP = ~cip;  //complement 
assign EAO = DAO & CCM ; 
assign eao = ~EAO ; //complement 
assign ECO = DAO & CCN ; 
assign eco = ~ECO ;  //complement 
assign EEO = DAO & CCO ; 
assign eeo = ~EEO ;  //complement 
assign EGO = DAO & CCP; 
assign ego = ~EGO; 
assign EEN = DAN & CCP ; 
assign een = ~EEN ; //complement 
assign EAN = DAN & CCN ; 
assign ean = ~EAN ;  //complement 
assign ECN = DAN & CCO ; 
assign ecn = ~ECN ;  //complement 
assign dal = ~DAL;  //complement 
assign dam = ~DAM;  //complement 
assign dan = ~DAN;  //complement 
assign dao = ~DAO;  //complement 
assign ddo = ~DDO;  //complement 
assign ddp = ~DDP;  //complement 
assign EAP = DAP & CCL ; 
assign eap = ~EAP ; //complement 
assign ECP = DAP & CCM ; 
assign ecp = ~ECP ;  //complement 
assign EEP = DAP & CCN ; 
assign eep = ~EEP ;  //complement 
assign EGP = DAP & CCO; 
assign egp = ~EGP; 
assign dap = ~DAP;  //complement 
assign EAQ = DBA & CCK ; 
assign eaq = ~EAQ ; //complement 
assign ECQ = DBA & CCL ; 
assign ecq = ~ECQ ;  //complement 
assign EEQ = DBA & CCM ; 
assign eeq = ~EEQ ;  //complement 
assign EGQ = DBA & CCN; 
assign egq = ~EGQ; 
assign dba = ~DBA;  //complement 
assign dea = ~DEA;  //complement 
assign DHA = ~dha;  //complement 
assign EAR = DBB & CCJ ; 
assign ear = ~EAR ; //complement 
assign ECR = DBB & CCK ; 
assign ecr = ~ECR ;  //complement 
assign EER = DBB & CCL ; 
assign eer = ~EER ;  //complement 
assign EGR = DBB & CCM; 
assign egr = ~EGR; 
assign EIR = DEB & CFN ; 
assign eir = ~EIR ; //complement 
assign EKR = DEB & CFO ; 
assign ekr = ~EKR ;  //complement 
assign EMR = DEB & CFP ; 
assign emr = ~EMR ;  //complement 
assign dbb = ~DBB;  //complement 
assign deb = ~DEB;  //complement 
assign DHB = ~dhb;  //complement 
assign LGA =  KFA & kga & kgc  |  kfa & KGA & kgc  |  kfa & kga & KGC  |  KFA & KGA & KGC  ; 
assign lga = ~LGA; //complement 
assign lha =  KFA & kga & kgc  |  kfa & KGA & kgc  |  kfa & kga & KGC  |  kfa & kga & kgc  ; 
assign LHA = ~lha;  //complement 
assign JEA =  HEB & hef & hda  |  heb & HEF & hda  |  heb & hef & HDA  |  HEB & HEF & HDA  ; 
assign jea = ~JEA; //complement 
assign jfa =  HEB & hef & hda  |  heb & HEF & hda  |  heb & hef & HDA  |  heb & hef & hda  ; 
assign JFA = ~jfa;  //complement 
assign haf = ~HAF;  //complement 
assign HBF = ~hbf;  //complement 
assign hag = ~HAG;  //complement 
assign GCB =  FBD & fcd & fcj  |  fbd & FCD & fcj  |  fbd & fcd & FCJ  |  FBD & FCD & FCJ  ; 
assign gcb = ~GCB; //complement 
assign gdb =  FBD & fcd & fcj  |  fbd & FCD & fcj  |  fbd & fcd & FCJ  |  fbd & fcd & fcj  ; 
assign GDB = ~gdb;  //complement 
assign LOB =  KOA & koc & kob  |  koa & KOC & kob  |  koa & koc & KOB  |  KOA & KOC & KOB  ; 
assign lob = ~LOB; //complement 
assign lpb =  KOA & koc & kob  |  koa & KOC & kob  |  koa & koc & KOB  |  koa & koc & kob  ; 
assign LPB = ~lpb;  //complement 
assign JIB =  HIC & hhc & hhb  |  hic & HHC & hhb  |  hic & hhc & HHB  |  HIC & HHC & HHB  ; 
assign jib = ~JIB; //complement 
assign jjb =  HIC & hhc & hhb  |  hic & HHC & hhb  |  hic & hhc & HHB  |  hic & hhc & hhb  ; 
assign JJB = ~jjb;  //complement 
assign hed = ~HED;  //complement 
assign HFD = ~hfd;  //complement 
assign GEB =  FEB & feh & fdd  |  feb & FEH & fdd  |  feb & feh & FDD  |  FEB & FEH & FDD  ; 
assign geb = ~GEB; //complement 
assign gfb =  FEB & feh & fdd  |  feb & FEH & fdd  |  feb & feh & FDD  |  feb & feh & fdd  ; 
assign GFB = ~gfb;  //complement 
assign mga = ~MGA;  //complement 
assign MHA = ~mha;  //complement 
assign mgb = ~MGB;  //complement 
assign JMC =  HLE & hme & hld  |  hle & HME & hld  |  hle & hme & HLD  |  HLE & HME & HLD  ; 
assign jmc = ~JMC; //complement 
assign jnc =  HLE & hme & hld  |  hle & HME & hld  |  hle & hme & HLD  |  hle & hme & hld  ; 
assign JNC = ~jnc;  //complement 
assign hib = ~HIB;  //complement 
assign HJB = ~hjb;  //complement 
assign GGB =  FGD & ffg & fgl  |  fgd & FFG & fgl  |  fgd & ffg & FGL  |  FGD & FFG & FGL  ; 
assign ggb = ~GGB; //complement 
assign ghb =  FGD & ffg & fgl  |  fgd & FFG & fgl  |  fgd & ffg & FGL  |  fgd & ffg & fgl  ; 
assign GHB = ~ghb;  //complement 
assign JSB =  HSC & hrd & hrc  |  hsc & HRD & hrc  |  hsc & hrd & HRC  |  HSC & HRD & HRC  ; 
assign jsb = ~JSB; //complement 
assign jtb =  HSC & hrd & hrc  |  hsc & HRD & hrc  |  hsc & hrd & HRC  |  hsc & hrd & hrc  ; 
assign JTB = ~jtb;  //complement 
assign hke = ~HKE;  //complement 
assign HLE = ~hle;  //complement 
assign GIB =  FHA & fid & fhd  |  fha & FID & fhd  |  fha & fid & FHD  |  FHA & FID & FHD  ; 
assign gib = ~GIB; //complement 
assign gjb =  FHA & fid & fhd  |  fha & FID & fhd  |  fha & fid & FHD  |  fha & fid & fhd  ; 
assign GJB = ~gjb;  //complement 
assign ohe = ~OHE;  //complement 
assign OIE = ~oie;  //complement 
assign kad = ~KAD;  //complement 
assign KBD = ~kbd;  //complement 
assign kae = ~KAE;  //complement 
assign hoc = ~HOC;  //complement 
assign HPC = ~hpc;  //complement 
assign hoe = ~HOE;  //complement 
assign GKC =  FKJ & fjh & fke  |  fkj & FJH & fke  |  fkj & fjh & FKE  |  FKJ & FJH & FKE  ; 
assign gkc = ~GKC; //complement 
assign glc =  FKJ & fjh & fke  |  fkj & FJH & fke  |  fkj & fjh & FKE  |  fkj & fjh & fke  ; 
assign GLC = ~glc;  //complement 
assign opm = ~OPM;  //complement 
assign OQM = ~oqm;  //complement 
assign kia = ~KIA;  //complement 
assign KJA = ~kja;  //complement 
assign kic = ~KIC;  //complement 
assign hsb = ~HSB;  //complement 
assign HTB = ~htb;  //complement 
assign GMD =  FMC & fmh & fmb  |  fmc & FMH & fmb  |  fmc & fmh & FMB  |  FMC & FMH & FMB  ; 
assign gmd = ~GMD; //complement 
assign gnd =  FMC & fmh & fmb  |  fmc & FMH & fmb  |  fmc & fmh & FMB  |  fmc & fmh & fmb  ; 
assign GND = ~gnd;  //complement 
assign kqa = ~KQA;  //complement 
assign KRA = ~kra;  //complement 
assign GOE =  FOB & fnc & foh  |  fob & FNC & foh  |  fob & fnc & FOH  |  FOB & FNC & FOH  ; 
assign goe = ~GOE; //complement 
assign gpe =  FOB & fnc & foh  |  fob & FNC & foh  |  fob & fnc & FOH  |  fob & fnc & foh  ; 
assign GPE = ~gpe;  //complement 
assign GQA =  FQA & fpa & fqg  |  fqa & FPA & fqg  |  fqa & fpa & FQG  |  FQA & FPA & FQG  ; 
assign gqa = ~GQA; //complement 
assign gra =  FQA & fpa & fqg  |  fqa & FPA & fqg  |  fqa & fpa & FQG  |  fqa & fpa & fqg  ; 
assign GRA = ~gra;  //complement 
assign GUB =  FUB & fta & fug  |  fub & FTA & fug  |  fub & fta & FUG  |  FUB & FTA & FUG  ; 
assign gub = ~GUB; //complement 
assign gvb =  FUB & fta & fug  |  fub & FTA & fug  |  fub & fta & FUG  |  fub & fta & fug  ; 
assign GVB = ~gvb;  //complement 
assign GQF =  FQF & fpf & fqj  |  fqf & FPF & fqj  |  fqf & fpf & FQJ  |  FQF & FPF & FQJ  ; 
assign gqf = ~GQF; //complement 
assign grf =  FQF & fpf & fqj  |  fqf & FPF & fqj  |  fqf & fpf & FQJ  |  fqf & fpf & fqj  ; 
assign GRF = ~grf;  //complement 
assign fqe = ~FQE;  //complement 
assign FRE = ~fre;  //complement 
assign fee = ~FEE;  //complement 
assign FFE = ~ffe;  //complement 
assign fsg = ~FSG;  //complement 
assign FTG = ~ftg;  //complement 
assign fak = ~FAK;  //complement 
assign FBK = ~fbk;  //complement 
assign fan = ~FAN;  //complement 
assign fal = ~FAL;  //complement 
assign FBL = ~fbl;  //complement 
assign fqj = ~FQJ;  //complement 
assign FRJ = ~frj;  //complement 
assign fcj = ~FCJ;  //complement 
assign FDJ = ~fdj;  //complement 
assign fck = ~FCK;  //complement 
assign FDK = ~fdk;  //complement 
assign fse = ~FSE;  //complement 
assign FTE = ~fte;  //complement 
assign EQU = DHE & CIO ; 
assign equ = ~EQU ; //complement 
assign ESU = DHE & CIP ; 
assign esu = ~ESU ;  //complement 
assign EQT = DHD & CIP ; 
assign eqt = ~EQT ;  //complement 
assign fsf = ~FSF;  //complement 
assign FTF = ~ftf;  //complement 
assign fej = ~FEJ;  //complement 
assign FFJ = ~ffj;  //complement 
assign fuc = ~FUC;  //complement 
assign OGC = ~ogc;  //complement 
assign fel = ~FEL;  //complement 
assign FFL = ~ffl;  //complement 
assign fge = ~FGE;  //complement 
assign FHE = ~fhe;  //complement 
assign fgj = ~FGJ;  //complement 
assign FHJ = ~fhj;  //complement 
assign fgl = ~FGL;  //complement 
assign fuh = ~FUH;  //complement 
assign OGH = ~ogh;  //complement 
assign fui = ~FUI;  //complement 
assign OGI = ~ogi;  //complement 
assign fuj = ~FUJ;  //complement 
assign fie = ~FIE;  //complement 
assign FJE = ~fje;  //complement 
assign EQW = DHG & CIM ; 
assign eqw = ~EQW ; //complement 
assign ESW = DHG & CIN ; 
assign esw = ~ESW ;  //complement 
assign EUW = DHG & CIO ; 
assign euw = ~EUW ;  //complement 
assign fik = ~FIK;  //complement 
assign FJK = ~fjk;  //complement 
assign fil = ~FIL;  //complement 
assign fek = ~FEK;  //complement 
assign FFK = ~ffk;  //complement 
assign fke = ~FKE;  //complement 
assign FLE = ~fle;  //complement 
assign EQX = DHH & CIL ; 
assign eqx = ~EQX ; //complement 
assign ESX = DHH & CIM ; 
assign esx = ~ESX ;  //complement 
assign EUX = DHH & CIN ; 
assign eux = ~EUX ;  //complement 
assign fkk = ~FKK;  //complement 
assign FLK = ~flk;  //complement 
assign EQV = DHF & CIN ; 
assign eqv = ~EQV ; //complement 
assign ESV = DHF & CIO ; 
assign esv = ~ESV ;  //complement 
assign EUV = DHF & CIP ; 
assign euv = ~EUV ;  //complement 
assign fme = ~FME;  //complement 
assign FNE = ~fne;  //complement 
assign ERA = DHI & CIK ; 
assign era = ~ERA ; //complement 
assign ETA = DHI & CIL ; 
assign eta = ~ETA ;  //complement 
assign EVA = DHI & CIM ; 
assign eva = ~EVA ;  //complement 
assign fmj = ~FMJ;  //complement 
assign FNJ = ~fnj;  //complement 
assign fml = ~FML;  //complement 
assign foe = ~FOE;  //complement 
assign FPE = ~fpe;  //complement 
assign ERB = DHJ & CIJ ; 
assign erb = ~ERB ; //complement 
assign ETB = DHJ & CIK ; 
assign etb = ~ETB ;  //complement 
assign EVB = DHJ & CIL ; 
assign evb = ~EVB ;  //complement 
assign foj = ~FOJ;  //complement 
assign FPJ = ~fpj;  //complement 
assign fok = ~FOK;  //complement 
assign EIS = DEC & CFM ; 
assign eis = ~EIS ; //complement 
assign EKS = DEC & CFN ; 
assign eks = ~EKS ;  //complement 
assign EMS = DEC & CFO ; 
assign ems = ~EMS ;  //complement 
assign EOS = DEC & CFP; 
assign eos = ~EOS; 
assign ERN = DIF & CHN ; 
assign ern = ~ERN ; //complement 
assign ETN = DIF & CHO ; 
assign etn = ~ETN ;  //complement 
assign EVN = DIF & CHP ; 
assign evn = ~EVN ;  //complement 
assign EAS = DBC & CCI ; 
assign eas = ~EAS ; //complement 
assign ECS = DBC & CCJ ; 
assign ecs = ~ECS ;  //complement 
assign EES = DBC & CCK ; 
assign ees = ~EES ;  //complement 
assign EGS = DBC & CCL; 
assign egs = ~EGS; 
assign dbc = ~DBC;  //complement 
assign dec = ~DEC;  //complement 
assign DHC = ~dhc;  //complement 
assign EIT = DED & CFL ; 
assign eit = ~EIT ; //complement 
assign EKT = DED & CFM ; 
assign ekt = ~EKT ;  //complement 
assign EMT = DED & CFN ; 
assign emt = ~EMT ;  //complement 
assign EOT = DED & CFO; 
assign eot = ~EOT; 
assign ERM = DIE & CHO ; 
assign erm = ~ERM ; //complement 
assign ETM = DIE & CHP ; 
assign etm = ~ETM ;  //complement 
assign EVM = DIE & CIA ; 
assign evm = ~EVM ;  //complement 
assign EAT = DBD & CCH ; 
assign eat = ~EAT ; //complement 
assign ECT = DBD & CCI ; 
assign ect = ~ECT ;  //complement 
assign EET = DBD & CCJ ; 
assign eet = ~EET ;  //complement 
assign EGT = DBD & CCK; 
assign egt = ~EGT; 
assign dbd = ~DBD;  //complement 
assign ded = ~DED;  //complement 
assign DHD = ~dhd;  //complement 
assign EIU = DEE & CFK ; 
assign eiu = ~EIU ; //complement 
assign EKU = DEE & CFL ; 
assign eku = ~EKU ;  //complement 
assign EMU = DEE & CFM ; 
assign emu = ~EMU ;  //complement 
assign EOU = DEE & CFN; 
assign eou = ~EOU; 
assign dca = ~DCA;  //complement 
assign dfa = ~DFA;  //complement 
assign DIA = ~dia;  //complement 
assign EAU = DBE & CCG ; 
assign eau = ~EAU ; //complement 
assign ECU = DBE & CCH ; 
assign ecu = ~ECU ;  //complement 
assign EEU = DBE & CCI ; 
assign eeu = ~EEU ;  //complement 
assign EGU = DBE & CCJ; 
assign egu = ~EGU; 
assign dbe = ~DBE;  //complement 
assign dee = ~DEE;  //complement 
assign DHE = ~dhe;  //complement 
assign EIV = DEF & CFJ ; 
assign eiv = ~EIV ; //complement 
assign EKV = DEF & CFK ; 
assign ekv = ~EKV ;  //complement 
assign EMV = DEF & CFL ; 
assign emv = ~EMV ;  //complement 
assign EOV = DEF & CFM; 
assign eov = ~EOV; 
assign EBJ = DCB & CBJ ; 
assign ebj = ~EBJ ; //complement 
assign EDJ = DCB & CBK ; 
assign edj = ~EDJ ;  //complement 
assign EFJ = DCB & CBL ; 
assign efj = ~EFJ ;  //complement 
assign EHJ = DCB & CBM; 
assign ehj = ~EHJ; 
assign EAV = DBF & CCF ; 
assign eav = ~EAV ; //complement 
assign ECV = DBF & CCG ; 
assign ecv = ~ECV ;  //complement 
assign EEV = DBF & CCH ; 
assign eev = ~EEV ;  //complement 
assign EGV = DBF & CCI; 
assign egv = ~EGV; 
assign dbf = ~DBF;  //complement 
assign def = ~DEF;  //complement 
assign DHF = ~dhf;  //complement 
assign EIW = DEG & CFI ; 
assign eiw = ~EIW ; //complement 
assign EKW = DEG & CFJ ; 
assign ekw = ~EKW ;  //complement 
assign EMW = DEG & CFK ; 
assign emw = ~EMW ;  //complement 
assign EOW = DEG & CFL; 
assign eow = ~EOW; 
assign EBC = DBK & CCA ; 
assign ebc = ~EBC ; //complement 
assign EDC = DBK & CCB ; 
assign edc = ~EDC ;  //complement 
assign EFC = DBK & CCC ; 
assign efc = ~EFC ;  //complement 
assign EHC = DBK & CCD; 
assign ehc = ~EHC; 
assign EAW = DBG & CCE ; 
assign eaw = ~EAW ; //complement 
assign ECW = DBG & CCF ; 
assign ecw = ~ECW ;  //complement 
assign EEW = DBG & CCG ; 
assign eew = ~EEW ;  //complement 
assign EGW = DBG & CCH; 
assign egw = ~EGW; 
assign dbg = ~DBG;  //complement 
assign deg = ~DEG;  //complement 
assign DHG = ~dhg;  //complement 
assign EIX = DEH & CFH ; 
assign eix = ~EIX ; //complement 
assign EKX = DEH & CFI ; 
assign ekx = ~EKX ;  //complement 
assign EMX = DEH & CFJ ; 
assign emx = ~EMX ;  //complement 
assign EOX = DEH & CFK; 
assign eox = ~EOX; 
assign ERJ = DIB & CIB ; 
assign erj = ~ERJ ; //complement 
assign ETJ = DIB & CIC ; 
assign etj = ~ETJ ;  //complement 
assign EVJ = DIB & CID ; 
assign evj = ~EVJ ;  //complement 
assign dbk = ~DBK;  //complement 
assign dek = ~DEK;  //complement 
assign DHK = ~dhk;  //complement 
assign dbh = ~DBH;  //complement 
assign deh = ~DEH;  //complement 
assign DHH = ~dhh;  //complement 
assign EJA = DEI & CFG ; 
assign eja = ~EJA ; //complement 
assign ELA = DEI & CFH ; 
assign ela = ~ELA ;  //complement 
assign ENA = DEI & CFI ; 
assign ena = ~ENA ;  //complement 
assign EPA = DEI & CFJ; 
assign epa = ~EPA; 
assign fkj = ~FKJ;  //complement 
assign FLJ = ~flj;  //complement 
assign EAX = DBH & CCD ; 
assign eax = ~EAX ; //complement 
assign ECX = DBH & CCE ; 
assign ecx = ~ECX ;  //complement 
assign EEX = DBH & CCF ; 
assign eex = ~EEX ;  //complement 
assign EGX = DBH & CCG; 
assign egx = ~EGX; 
assign dbi = ~DBI;  //complement 
assign dei = ~DEI;  //complement 
assign DHI = ~dhi;  //complement 
assign EJB = DEJ & CFF ; 
assign ejb = ~EJB ; //complement 
assign ELB = DEJ & CFG ; 
assign elb = ~ELB ;  //complement 
assign ENB = DEJ & CFH ; 
assign enb = ~ENB ;  //complement 
assign EPB = DEJ & CFI; 
assign epb = ~EPB; 
assign EBB = DBJ & CCB ; 
assign ebb = ~EBB ; //complement 
assign EDB = DBJ & CCC ; 
assign edb = ~EDB ;  //complement 
assign EFB = DBJ & CCD ; 
assign efb = ~EFB ;  //complement 
assign EHB = DBJ & CCE; 
assign ehb = ~EHB; 
assign EBA = DBI & CCC ; 
assign eba = ~EBA ; //complement 
assign EDA = DBI & CCD ; 
assign eda = ~EDA ;  //complement 
assign EFA = DBI & CCE ; 
assign efa = ~EFA ;  //complement 
assign EHA = DBI & CCF; 
assign eha = ~EHA; 
assign dbj = ~DBJ;  //complement 
assign dej = ~DEJ;  //complement 
assign DHJ = ~dhj;  //complement 
assign LIA =  KIA & kic & kha  |  kia & KIC & kha  |  kia & kic & KHA  |  KIA & KIC & KHA  ; 
assign lia = ~LIA; //complement 
assign lja =  KIA & kic & kha  |  kia & KIC & kha  |  kia & kic & KHA  |  kia & kic & kha  ; 
assign LJA = ~lja;  //complement 
assign JEB =  HEC & hed & hdb  |  hec & HED & hdb  |  hec & hed & HDB  |  HEC & HED & HDB  ; 
assign jeb = ~JEB; //complement 
assign jfb =  HEC & hed & hdb  |  hec & HED & hdb  |  hec & hed & HDB  |  hec & hed & hdb  ; 
assign JFB = ~jfb;  //complement 
assign hca = ~HCA;  //complement 
assign HDA = ~hda;  //complement 
assign GCC =  FBB & fbh & fce  |  fbb & FBH & fce  |  fbb & fbh & FCE  |  FBB & FBH & FCE  ; 
assign gcc = ~GCC; //complement 
assign gdc =  FBB & fbh & fce  |  fbb & FBH & fce  |  fbb & fbh & FCE  |  fbb & fbh & fce  ; 
assign GDC = ~gdc;  //complement 
assign LQA =  KPA & kpb & kqb  |  kpa & KPB & kqb  |  kpa & kpb & KQB  |  KPA & KPB & KQB  ; 
assign lqa = ~LQA; //complement 
assign lra =  KPA & kpb & kqb  |  kpa & KPB & kqb  |  kpa & kpb & KQB  |  kpa & kpb & kqb  ; 
assign LRA = ~lra;  //complement 
assign JIC =  HID & hig & hhe  |  hid & HIG & hhe  |  hid & hig & HHE  |  HID & HIG & HHE  ; 
assign jic = ~JIC; //complement 
assign jjc =  HID & hig & hhe  |  hid & HIG & hhe  |  hid & hig & HHE  |  hid & hig & hhe  ; 
assign JJC = ~jjc;  //complement 
assign hee = ~HEE;  //complement 
assign HFE = ~hfe;  //complement 
assign hef = ~HEF;  //complement 
assign GEC =  FDB & fdg & fde  |  fdb & FDG & fde  |  fdb & fdg & FDE  |  FDB & FDG & FDE  ; 
assign gec = ~GEC; //complement 
assign gfc =  FDB & fdg & fde  |  fdb & FDG & fde  |  fdb & fdg & FDE  |  fdb & fdg & fde  ; 
assign GFC = ~gfc;  //complement 
assign mia = ~MIA;  //complement 
assign MJA = ~mja;  //complement 
assign JOA =  HOA & hof & hna  |  hoa & HOF & hna  |  hoa & hof & HNA  |  HOA & HOF & HNA  ; 
assign joa = ~JOA; //complement 
assign jpa =  HOA & hof & hna  |  hoa & HOF & hna  |  hoa & hof & HNA  |  hoa & hof & hna  ; 
assign JPA = ~jpa;  //complement 
assign hic = ~HIC;  //complement 
assign HJC = ~hjc;  //complement 
assign GGC =  FFB & ffh & ffj  |  ffb & FFH & ffj  |  ffb & ffh & FFJ  |  FFB & FFH & FFJ  ; 
assign ggc = ~GGC; //complement 
assign ghc =  FFB & ffh & ffj  |  ffb & FFH & ffj  |  ffb & ffh & FFJ  |  ffb & ffh & ffj  ; 
assign GHC = ~ghc;  //complement 
assign mua = ~MUA;  //complement 
assign OMA = ~oma;  //complement 
assign mub = ~MUB;  //complement 
assign JSC =  HSD & hse & hre  |  hsd & HSE & hre  |  hsd & hse & HRE  |  HSD & HSE & HRE  ; 
assign jsc = ~JSC; //complement 
assign jtc =  HSD & hse & hre  |  hsd & HSE & hre  |  hsd & hse & HRE  |  hsd & hse & hre  ; 
assign JTC = ~jtc;  //complement 
assign hma = ~HMA;  //complement 
assign HNA = ~hna;  //complement 
assign GIC =  FIH & fib & fhj  |  fih & FIB & fhj  |  fih & fib & FHJ  |  FIH & FIB & FHJ  ; 
assign gic = ~GIC; //complement 
assign gjc =  FIH & fib & fhj  |  fih & FIB & fhj  |  fih & fib & FHJ  |  fih & fib & fhj  ; 
assign GJC = ~gjc;  //complement 
assign ohf = ~OHF;  //complement 
assign OIF = ~oif;  //complement 
assign kca = ~KCA;  //complement 
assign KDA = ~kda;  //complement 
assign hod = ~HOD;  //complement 
assign HPD = ~hpd;  //complement 
assign hof = ~HOF;  //complement 
assign GKD =  FKB & fkh & fje  |  fkb & FKH & fje  |  fkb & fkh & FJE  |  FKB & FKH & FJE  ; 
assign gkd = ~GKD; //complement 
assign gld =  FKB & fkh & fje  |  fkb & FKH & fje  |  fkb & fkh & FJE  |  fkb & fkh & fje  ; 
assign GLD = ~gld;  //complement 
assign opo = ~OPO;  //complement 
assign OQO = ~oqo;  //complement 
assign kib = ~KIB;  //complement 
assign KJB = ~kjb;  //complement 
assign kid = ~KID;  //complement 
assign hsc = ~HSC;  //complement 
assign HTC = ~htc;  //complement 
assign GME =  FMK & flh & fml  |  fmk & FLH & fml  |  fmk & flh & FML  |  FMK & FLH & FML  ; 
assign gme = ~GME; //complement 
assign gne =  FMK & flh & fml  |  fmk & FLH & fml  |  fmk & flh & FML  |  fmk & flh & fml  ; 
assign GNE = ~gne;  //complement 
assign kqb = ~KQB;  //complement 
assign KRB = ~krb;  //complement 
assign GOF =  FNB & foc & fnf  |  fnb & FOC & fnf  |  fnb & foc & FNF  |  FNB & FOC & FNF  ; 
assign gof = ~GOF; //complement 
assign gpf =  FNB & foc & fnf  |  fnb & FOC & fnf  |  fnb & foc & FNF  |  fnb & foc & fnf  ; 
assign GPF = ~gpf;  //complement 
assign GUC =  FTD & ftf & fth  |  ftd & FTF & fth  |  ftd & ftf & FTH  |  FTD & FTF & FTH  ; 
assign guc = ~GUC; //complement 
assign gvc =  FTD & ftf & fth  |  ftd & FTF & fth  |  ftd & ftf & FTH  |  ftd & ftf & fth  ; 
assign GVC = ~gvc;  //complement 
assign GSA =  FRD & fra & frg  |  frd & FRA & frg  |  frd & fra & FRG  |  FRD & FRA & FRG  ; 
assign gsa = ~GSA; //complement 
assign gta =  FRD & fra & frg  |  frd & FRA & frg  |  frd & fra & FRG  |  frd & fra & frg  ; 
assign GTA = ~gta;  //complement 
assign EJC = DEK & CFE ; 
assign ejc = ~EJC ; //complement 
assign ELC = DEK & CFF ; 
assign elc = ~ELC ;  //complement 
assign ENC = DEK & CFG ; 
assign enc = ~ENC ;  //complement 
assign EPC = DEK & CFH; 
assign epc = ~EPC; 
assign ERS = DIK & CHI ; 
assign ers = ~ERS ; //complement 
assign ETS = DIK & CHJ ; 
assign ets = ~ETS ;  //complement 
assign EVS = DIK & CHK ; 
assign evs = ~EVS ;  //complement 
assign ERK = DIC & CIA ; 
assign erk = ~ERK ; //complement 
assign ETK = DIC & CIB ; 
assign etk = ~ETK ;  //complement 
assign EVK = DIC & CIC ; 
assign evk = ~EVK ;  //complement 
assign ERC = DHK & CII ; 
assign erc = ~ERC ; //complement 
assign ETC = DHK & CIJ ; 
assign etc = ~ETC ;  //complement 
assign EVC = DHK & CIK ; 
assign evc = ~EVC ;  //complement 
assign EJD = DEL & CFD ; 
assign ejd = ~EJD ; //complement 
assign ELD = DEL & CFE ; 
assign eld = ~ELD ;  //complement 
assign ENDD  = DEL & CFF ; 
assign endd = ~ENDD  ;  //complement 
assign EPD = DEL & CFG; 
assign epd = ~EPD; 
assign ERQ = DII & CHK ; 
assign erq = ~ERQ ; //complement 
assign ETQ = DII & CHL ; 
assign etq = ~ETQ ;  //complement 
assign EVQ = DII & CHM ; 
assign evq = ~EVQ ;  //complement 
assign ERL = DID & CHP ; 
assign erl = ~ERL ; //complement 
assign ETL = DID & CIA ; 
assign etl = ~ETL ;  //complement 
assign EVL = DID & CIB ; 
assign evl = ~EVL ;  //complement 
assign ERD = DHL & CIH ; 
assign erd = ~ERD ; //complement 
assign ETD = DHL & CII ; 
assign etd = ~ETD ;  //complement 
assign EVD = DHL & CIJ ; 
assign evd = ~EVD ;  //complement 
assign EJE = DEM & CFC ; 
assign eje = ~EJE ; //complement 
assign ELE = DEM & CFD ; 
assign ele = ~ELE ;  //complement 
assign ENE = DEM & CFE ; 
assign ene = ~ENE ;  //complement 
assign EPE = DEM & CFF; 
assign epe = ~EPE; 
assign dbl = ~DBL;  //complement 
assign del = ~DEL;  //complement 
assign DHL = ~dhl;  //complement 
assign EBE = DBM & CBO ; 
assign ebe = ~EBE ; //complement 
assign EDE = DBM & CBP ; 
assign ede = ~EDE ;  //complement 
assign EFE = DBM & CCA ; 
assign efe = ~EFE ;  //complement 
assign EHE = DBM & CCB; 
assign ehe = ~EHE; 
assign ERE = DHM & CIG ; 
assign ere = ~ERE ; //complement 
assign ETE = DHM & CIH ; 
assign ete = ~ETE ;  //complement 
assign EVE = DHM & CII ; 
assign eve = ~EVE ;  //complement 
assign EJF = DEN & CFB ; 
assign ejf = ~EJF ; //complement 
assign ELF = DEN & CFC ; 
assign elf = ~ELF ;  //complement 
assign ENF = DEN & CFD ; 
assign enf = ~ENF ;  //complement 
assign EPF = DEN & CFE; 
assign epf = ~EPF; 
assign dbm = ~DBM;  //complement 
assign dem = ~DEM;  //complement 
assign DHM = ~dhm;  //complement 
assign EBF = DBN & CBN ; 
assign ebf = ~EBF ; //complement 
assign EDF = DBN & CBO ; 
assign edf = ~EDF ;  //complement 
assign EFF = DBN & CBP ; 
assign eff = ~EFF ;  //complement 
assign EHF = DBN & CCA; 
assign ehf = ~EHF; 
assign ERF = DHN & CIF ; 
assign erf = ~ERF ; //complement 
assign ETF = DHN & CIG ; 
assign etf = ~ETF ;  //complement 
assign EVF = DHN & CIH ; 
assign evf = ~EVF ;  //complement 
assign EJG = DEO & CFA ; 
assign ejg = ~EJG ; //complement 
assign ELG = DEO & CFB ; 
assign elg = ~ELG ;  //complement 
assign ENG = DEO & CFC ; 
assign eng = ~ENG ;  //complement 
assign EPG = DEO & CFD; 
assign epg = ~EPG; 
assign ERV = DIN & CHF ; 
assign erv = ~ERV ; //complement 
assign ETV = DIN & CHG ; 
assign etv = ~ETV ;  //complement 
assign EVV = DIN & CHH ; 
assign evv = ~EVV ;  //complement 
assign EBG = DBO & CBM ; 
assign ebg = ~EBG ; //complement 
assign EDG = DBO & CBN ; 
assign edg = ~EDG ;  //complement 
assign EFG = DBO & CBO ; 
assign efg = ~EFG ;  //complement 
assign EHG = DBO & CBP; 
assign ehg = ~EHG; 
assign ERO = DIG & CHM ; 
assign ero = ~ERO ; //complement 
assign ETO = DIG & CHN ; 
assign eto = ~ETO ;  //complement 
assign EVO = DIG & CHO ; 
assign evo = ~EVO ;  //complement 
assign EJH = DEP & CEP ; 
assign ejh = ~EJH ; //complement 
assign ELH = DEP & CFA ; 
assign elh = ~ELH ;  //complement 
assign ENH = DEP & CFB ; 
assign enh = ~ENH ;  //complement 
assign EPH = DEP & CFC; 
assign eph = ~EPH; 
assign dbn = ~DBN;  //complement 
assign den = ~DEN;  //complement 
assign DHN = ~dhn;  //complement 
assign EBH = DBP & CBL ; 
assign ebh = ~EBH ; //complement 
assign EDH = DBP & CBM ; 
assign edh = ~EDH ;  //complement 
assign EFH = DBP & CBN ; 
assign efh = ~EFH ;  //complement 
assign EHH = DBP & CBO; 
assign ehh = ~EHH; 
assign dbp = ~DBP;  //complement 
assign dep = ~DEP;  //complement 
assign DHP = ~dhp;  //complement 
assign EJI = DFA & CEO ; 
assign eji = ~EJI ; //complement 
assign ELI = DFA & CEP ; 
assign eli = ~ELI ;  //complement 
assign ENI = DFA & CFA ; 
assign eni = ~ENI ;  //complement 
assign EPI = DFA & CFB; 
assign epi = ~EPI; 
assign ERT = DIL & CHH ; 
assign ert = ~ERT ; //complement 
assign ETT = DIL & CHI ; 
assign ett = ~ETT ;  //complement 
assign EVT = DIL & CHJ ; 
assign evt = ~EVT ;  //complement 
assign EBI = DCA & CBK ; 
assign ebi = ~EBI ; //complement 
assign EDI = DCA & CBL ; 
assign edi = ~EDI ;  //complement 
assign EFI = DCA & CBM ; 
assign efi = ~EFI ;  //complement 
assign EHI = DCA & CBN; 
assign ehi = ~EHI; 
assign ERI = DIA & CIC ; 
assign eri = ~ERI ; //complement 
assign ETI = DIA & CID ; 
assign eti = ~ETI ;  //complement 
assign EVI = DIA & CIE ; 
assign evi = ~EVI ;  //complement 
assign EJJ = DFB & CEN ; 
assign ejj = ~EJJ ; //complement 
assign ELJ = DFB & CEO ; 
assign elj = ~ELJ ;  //complement 
assign ENJ = DFB & CEP ; 
assign enj = ~ENJ ;  //complement 
assign EPJ = DFB & CFA; 
assign epj = ~EPJ; 
assign ERU = DIM & CHG ; 
assign eru = ~ERU ; //complement 
assign ETU = DIM & CHH ; 
assign etu = ~ETU ;  //complement 
assign EVU = DIM & CHI ; 
assign evu = ~EVU ;  //complement 
assign ERR = DIJ & CHJ ; 
assign err = ~ERR ; //complement 
assign ETR = DIJ & CHK ; 
assign etr = ~ETR ;  //complement 
assign EVR = DIJ & CHL ; 
assign evr = ~EVR ;  //complement 
assign dcb = ~DCB;  //complement 
assign dfb = ~DFB;  //complement 
assign DIB = ~dib;  //complement 
assign LIB =  KIB & kid & khb  |  kib & KID & khb  |  kib & kid & KHB  |  KIB & KID & KHB  ; 
assign lib = ~LIB; //complement 
assign ljb =  KIB & kid & khb  |  kib & KID & khb  |  kib & kid & KHB  |  kib & kid & khb  ; 
assign LJB = ~ljb;  //complement 
assign JEC =  HDD & hee & hdc  |  hdd & HEE & hdc  |  hdd & hee & HDC  |  HDD & HEE & HDC  ; 
assign jec = ~JEC; //complement 
assign jfc =  HDD & hee & hdc  |  hdd & HEE & hdc  |  hdd & hee & HDC  |  hdd & hee & hdc  ; 
assign JFC = ~jfc;  //complement 
assign hcb = ~HCB;  //complement 
assign HDB = ~hdb;  //complement 
assign GCD =  FCC & fck & fcb  |  fcc & FCK & fcb  |  fcc & fck & FCB  |  FCC & FCK & FCB  ; 
assign gcd = ~GCD; //complement 
assign gdd =  FCC & fck & fcb  |  fcc & FCK & fcb  |  fcc & fck & FCB  |  fcc & fck & fcb  ; 
assign GDD = ~gdd;  //complement 
assign LSA =  KSB & ksc & krb  |  ksb & KSC & krb  |  ksb & ksc & KRB  |  KSB & KSC & KRB  ; 
assign lsa = ~LSA; //complement 
assign lta =  KSB & ksc & krb  |  ksb & KSC & krb  |  ksb & ksc & KRB  |  ksb & ksc & krb  ; 
assign LTA = ~lta;  //complement 
assign JID =  HIE & hif & hhd  |  hie & HIF & hhd  |  hie & hif & HHD  |  HIE & HIF & HHD  ; 
assign jid = ~JID; //complement 
assign jjd =  HIE & hif & hhd  |  hie & HIF & hhd  |  hie & hif & HHD  |  hie & hif & hhd  ; 
assign JJD = ~jjd;  //complement 
assign hga = ~HGA;  //complement 
assign HHA = ~hha;  //complement 
assign GED =  FED & fej & fdk  |  fed & FEJ & fdk  |  fed & fej & FDK  |  FED & FEJ & FDK  ; 
assign ged = ~GED; //complement 
assign gfd =  FED & fej & fdk  |  fed & FEJ & fdk  |  fed & fej & FDK  |  fed & fej & fdk  ; 
assign GFD = ~gfd;  //complement 
assign mka = ~MKA;  //complement 
assign MLA = ~mla;  //complement 
assign mkb = ~MKB;  //complement 
assign JOB =  HOB & hnd & hnb  |  hob & HND & hnb  |  hob & hnd & HNB  |  HOB & HND & HNB  ; 
assign job = ~JOB; //complement 
assign jpb =  HOB & hnd & hnb  |  hob & HND & hnb  |  hob & hnd & HNB  |  hob & hnd & hnb  ; 
assign JPB = ~jpb;  //complement 
assign hid = ~HID;  //complement 
assign HJD = ~hjd;  //complement 
assign hif = ~HIF;  //complement 
assign GGD =  FGJ & fge & ffd  |  fgj & FGE & ffd  |  fgj & fge & FFD  |  FGJ & FGE & FFD  ; 
assign ggd = ~GGD; //complement 
assign ghd =  FGJ & fge & ffd  |  fgj & FGE & ffd  |  fgj & fge & FFD  |  fgj & fge & ffd  ; 
assign GHD = ~ghd;  //complement 
assign NAA =  MAB & mac & mad  |  mab & MAC & mad  |  mab & mac & MAD  |  MAB & MAC & MAD  ; 
assign naa = ~NAA; //complement 
assign nba =  MAB & mac & mad  |  mab & MAC & mad  |  mab & mac & MAD  |  mab & mac & mad  ; 
assign NBA = ~nba;  //complement 
assign JUA =  HUA & hue & htb  |  hua & HUE & htb  |  hua & hue & HTB  |  HUA & HUE & HTB  ; 
assign jua = ~JUA; //complement 
assign jva =  HUA & hue & htb  |  hua & HUE & htb  |  hua & hue & HTB  |  hua & hue & htb  ; 
assign JVA = ~jva;  //complement 
assign hmb = ~HMB;  //complement 
assign HNB = ~hnb;  //complement 
assign GID =  FHB & fhh & fhe  |  fhb & FHH & fhe  |  fhb & fhh & FHE  |  FHB & FHH & FHE  ; 
assign gid = ~GID; //complement 
assign gjd =  FHB & fhh & fhe  |  fhb & FHH & fhe  |  fhb & fhh & FHE  |  fhb & fhh & fhe  ; 
assign GJD = ~gjd;  //complement 
assign okc = ~OKC;  //complement 
assign OLC = ~olc;  //complement 
assign kcb = ~KCB;  //complement 
assign KDB = ~kdb;  //complement 
assign hqa = ~HQA;  //complement 
assign HRA = ~hra;  //complement 
assign GKE =  FKF & fkk & fjj  |  fkf & FKK & fjj  |  fkf & fkk & FJJ  |  FKF & FKK & FJJ  ; 
assign gke = ~GKE; //complement 
assign gle =  FKF & fkk & fjj  |  fkf & FKK & fjj  |  fkf & fkk & FJJ  |  fkf & fkk & fjj  ; 
assign GLE = ~gle;  //complement 
assign opq = ~OPQ;  //complement 
assign OQQ = ~oqq;  //complement 
assign kka = ~KKA;  //complement 
assign KLA = ~kla;  //complement 
assign kkc = ~KKC;  //complement 
assign hsd = ~HSD;  //complement 
assign HTD = ~htd;  //complement 
assign hse = ~HSE;  //complement 
assign GMF =  FLC & fli & flk  |  flc & FLI & flk  |  flc & fli & FLK  |  FLC & FLI & FLK  ; 
assign gmf = ~GMF; //complement 
assign gnf =  FLC & fli & flk  |  flc & FLI & flk  |  flc & fli & FLK  |  flc & fli & flk  ; 
assign GNF = ~gnf;  //complement 
assign ERP = DIH & CHL ; 
assign erp = ~ERP ; //complement 
assign ETP = DIH & CHM ; 
assign etp = ~ETP ;  //complement 
assign EVP = DIH & CHN ; 
assign evp = ~EVP ;  //complement 
assign ksa = ~KSA;  //complement 
assign KTA = ~kta;  //complement 
assign ERG = DHO & CIE ; 
assign erg = ~ERG ; //complement 
assign ETG = DHO & CIF ; 
assign etg = ~ETG ;  //complement 
assign EVG = DHO & CIG ; 
assign evg = ~EVG ;  //complement 
assign GOG =  FOF & foj & fnj  |  fof & FOJ & fnj  |  fof & foj & FNJ  |  FOF & FOJ & FNJ  ; 
assign gog = ~GOG; //complement 
assign gpg =  FOF & foj & fnj  |  fof & FOJ & fnj  |  fof & foj & FNJ  |  fof & foj & fnj  ; 
assign GPG = ~gpg;  //complement 
assign GUF =  FUI & fue & ftc  |  fui & FUE & ftc  |  fui & fue & FTC  |  FUI & FUE & FTC  ; 
assign guf = ~GUF; //complement 
assign gvf =  FUI & fue & ftc  |  fui & FUE & ftc  |  fui & fue & FTC  |  fui & fue & ftc  ; 
assign GVF = ~gvf;  //complement 
assign GUE =  FUD & fuh & fti  |  fud & FUH & fti  |  fud & fuh & FTI  |  FUD & FUH & FTI  ; 
assign gue = ~GUE; //complement 
assign gve =  FUD & fuh & fti  |  fud & FUH & fti  |  fud & fuh & FTI  |  fud & fuh & fti  ; 
assign GVE = ~gve;  //complement 
assign GUD =  FUC & ftb & ftg  |  fuc & FTB & ftg  |  fuc & ftb & FTG  |  FUC & FTB & FTG  ; 
assign gud = ~GUD; //complement 
assign gvd =  FUC & ftb & ftg  |  fuc & FTB & ftg  |  fuc & ftb & FTG  |  fuc & ftb & ftg  ; 
assign GVD = ~gvd;  //complement 
assign dbo = ~DBO;  //complement 
assign deo = ~DEO;  //complement 
assign DHO = ~dho;  //complement 
assign EJS = DFK & CEE ; 
assign ejs = ~EJS ; //complement 
assign ELS = DFK & CEF ; 
assign els = ~ELS ;  //complement 
assign ENS = DFK & CEG ; 
assign ens = ~ENS ;  //complement 
assign EPS = DFK & CEH; 
assign eps = ~EPS; 
assign EBS = DCK & CBA ; 
assign ebs = ~EBS ; //complement 
assign EDS = DCK & CBB ; 
assign eds = ~EDS ;  //complement 
assign EFS = DCK & CBC ; 
assign efs = ~EFS ;  //complement 
assign EHS = DCK & CBD; 
assign ehs = ~EHS; 
assign EJT = DFL & CED ; 
assign ejt = ~EJT ; //complement 
assign ELT = DFL & CEE ; 
assign elt = ~ELT ;  //complement 
assign ENT = DFL & CEF ; 
assign ent = ~ENT ;  //complement 
assign EPT = DFL & CEG; 
assign ept = ~EPT; 
assign EBT = DCL & CAP ; 
assign ebt = ~EBT ; //complement 
assign EDT = DCL & CBA ; 
assign edt = ~EDT ;  //complement 
assign EFT = DCL & CBB ; 
assign eft = ~EFT ;  //complement 
assign EHT = DCL & CBC; 
assign eht = ~EHT; 
assign EJU = DFM & CEC ; 
assign eju = ~EJU ; //complement 
assign ELU = DFM & CED ; 
assign elu = ~ELU ;  //complement 
assign ENU = DFM & CEE ; 
assign enu = ~ENU ;  //complement 
assign EPU = DFM & CEF; 
assign epu = ~EPU; 
assign EBU = DCM & CAO ; 
assign ebu = ~EBU ; //complement 
assign EDU = DCM & CAP ; 
assign edu = ~EDU ;  //complement 
assign EFU = DCM & CBA ; 
assign efu = ~EFU ;  //complement 
assign EHU = DCM & CBB; 
assign ehu = ~EHU; 
assign EJV = DFN & CEB ; 
assign ejv = ~EJV ; //complement 
assign ELV = DFN & CEC ; 
assign elv = ~ELV ;  //complement 
assign ENV = DFN & CED ; 
assign env = ~ENV ;  //complement 
assign EPV = DFN & CEE; 
assign epv = ~EPV; 
assign EJW = DFO & CEA ; 
assign ejw = ~EJW ; //complement 
assign ELW = DFO & CEB ; 
assign elw = ~ELW ;  //complement 
assign ENW = DFO & CEC ; 
assign enw = ~ENW ;  //complement 
assign EPW = DFO & CED; 
assign epw = ~EPW; 
assign EBV = DCN & CAN ; 
assign ebv = ~EBV ; //complement 
assign EDV = DCN & CAO ; 
assign edv = ~EDV ;  //complement 
assign EFV = DCN & CAP ; 
assign efv = ~EFV ;  //complement 
assign EHV = DCN & CBA; 
assign ehv = ~EHV; 
assign EJX = DFP & CDP ; 
assign ejx = ~EJX ; //complement 
assign ELX = DFP & CEA ; 
assign elx = ~ELX ;  //complement 
assign ENX = DFP & CEB ; 
assign enx = ~ENX ;  //complement 
assign EPX = DFP & CEC; 
assign epx = ~EPX; 
assign EBW = DCO & CAM ; 
assign ebw = ~EBW ; //complement 
assign EDW = DCO & CAN ; 
assign edw = ~EDW ;  //complement 
assign EFW = DCO & CAO ; 
assign efw = ~EFW ;  //complement 
assign EHW = DCO & CAP; 
assign ehw = ~EHW; 
assign fgk = ~FGK;  //complement 
assign FHK = ~fhk;  //complement 
assign fgm = ~FGM;  //complement 
assign fij = ~FIJ;  //complement 
assign FJJ = ~fjj;  //complement 
assign EBX = DCP & CAL ; 
assign ebx = ~EBX ; //complement 
assign EDX = DCP & CAM ; 
assign edx = ~EDX ;  //complement 
assign EFX = DCP & CAN ; 
assign efx = ~EFX ;  //complement 
assign EHX = DCP & CAO; 
assign ehx = ~EHX; 
assign EIQ = DEA & CFO ; 
assign eiq = ~EIQ ; //complement 
assign EKQ = DEA & CFP ; 
assign ekq = ~EKQ ;  //complement 
assign EIP = DDP & CFP ; 
assign eip = ~EIP ;  //complement 
assign EBK = DCC & CBI ; 
assign ebk = ~EBK ; //complement 
assign EDK = DCC & CBJ ; 
assign edk = ~EDK ;  //complement 
assign EFK = DCC & CBK ; 
assign efk = ~EFK ;  //complement 
assign EHK = DCC & CBL; 
assign ehk = ~EHK; 
assign EJK = DFC & CEM ; 
assign ejk = ~EJK ; //complement 
assign ELK = DFC & CEN ; 
assign elk = ~ELK ;  //complement 
assign ENK = DFC & CEO ; 
assign enk = ~ENK ;  //complement 
assign EPK = DFC & CEP; 
assign epk = ~EPK; 
assign dck = ~DCK;  //complement 
assign dfk = ~DFK;  //complement 
assign DIK = ~dik;  //complement 
assign dcc = ~DCC;  //complement 
assign dfc = ~DFC;  //complement 
assign DIC = ~dic;  //complement 
assign EBL = DCD & CBH ; 
assign ebl = ~EBL ; //complement 
assign EDL = DCD & CBI ; 
assign edl = ~EDL ;  //complement 
assign EFL = DCD & CBJ ; 
assign efl = ~EFL ;  //complement 
assign EHL = DCD & CBK; 
assign ehl = ~EHL; 
assign EJL = DFD & CEL ; 
assign ejl = ~EJL ; //complement 
assign ELL = DFD & CEM ; 
assign ell = ~ELL ;  //complement 
assign ENL = DFD & CEN ; 
assign enl = ~ENL ;  //complement 
assign EPL = DFD & CEO; 
assign epl = ~EPL; 
assign dcl = ~DCL;  //complement 
assign dfl = ~DFL;  //complement 
assign DIL = ~dil;  //complement 
assign dcd = ~DCD;  //complement 
assign dfd = ~DFD;  //complement 
assign DID = ~did;  //complement 
assign EBM = DCE & CBG ; 
assign ebm = ~EBM ; //complement 
assign EDM = DCE & CBH ; 
assign edm = ~EDM ;  //complement 
assign EFM = DCE & CBI ; 
assign efm = ~EFM ;  //complement 
assign EHM = DCE & CBJ; 
assign ehm = ~EHM; 
assign EJM = DFE & CEK ; 
assign ejm = ~EJM ; //complement 
assign ELM = DFE & CEL ; 
assign elm = ~ELM ;  //complement 
assign ENM = DFE & CEM ; 
assign enm = ~ENM ;  //complement 
assign EPM = DFE & CEN; 
assign epm = ~EPM; 
assign dcm = ~DCM;  //complement 
assign dfm = ~DFM;  //complement 
assign DIM = ~dim;  //complement 
assign dce = ~DCE;  //complement 
assign dfe = ~DFE;  //complement 
assign DIE = ~die;  //complement 
assign EBN = DCF & CBF ; 
assign ebn = ~EBN ; //complement 
assign EDN = DCF & CBG ; 
assign edn = ~EDN ;  //complement 
assign EFN = DCF & CBH ; 
assign efn = ~EFN ;  //complement 
assign EHN = DCF & CBI; 
assign ehn = ~EHN; 
assign EJN = DFF & CEJ ; 
assign ejn = ~EJN ; //complement 
assign ELN = DFF & CEK ; 
assign eln = ~ELN ;  //complement 
assign ENN = DFF & CEL ; 
assign enn = ~ENN ;  //complement 
assign EPN = DFF & CEM; 
assign epn = ~EPN; 
assign dcn = ~DCN;  //complement 
assign dfn = ~DFN;  //complement 
assign DIN = ~din;  //complement 
assign dcf = ~DCF;  //complement 
assign dff = ~DFF;  //complement 
assign DIF = ~dif;  //complement 
assign EBO = DCG & CBE ; 
assign ebo = ~EBO ; //complement 
assign EDO = DCG & CBF ; 
assign edo = ~EDO ;  //complement 
assign EFO = DCG & CBG ; 
assign efo = ~EFO ;  //complement 
assign EHO = DCG & CBH; 
assign eho = ~EHO; 
assign EJO = DFG & CEI ; 
assign ejo = ~EJO ; //complement 
assign ELO = DFG & CEJ ; 
assign elo = ~ELO ;  //complement 
assign ENO = DFG & CEK ; 
assign eno = ~ENO ;  //complement 
assign EPO = DFG & CEL; 
assign epo = ~EPO; 
assign dco = ~DCO;  //complement 
assign dfo = ~DFO;  //complement 
assign DIO = ~dio;  //complement 
assign dcg = ~DCG;  //complement 
assign dfg = ~DFG;  //complement 
assign DIG = ~dig;  //complement 
assign EBP = DCH & CBD ; 
assign ebp = ~EBP ; //complement 
assign EDP = DCH & CBE ; 
assign edp = ~EDP ;  //complement 
assign EFP = DCH & CBF ; 
assign efp = ~EFP ;  //complement 
assign EHP = DCH & CBG; 
assign ehp = ~EHP; 
assign EJP = DFH & CEH ; 
assign ejp = ~EJP ; //complement 
assign ELP = DFH & CEI ; 
assign elp = ~ELP ;  //complement 
assign ENP = DFH & CEJ ; 
assign enp = ~ENP ;  //complement 
assign EPP = DFH & CEK; 
assign epp = ~EPP; 
assign dcp = ~DCP;  //complement 
assign dfp = ~DFP;  //complement 
assign DIP = ~dip;  //complement 
assign dch = ~DCH;  //complement 
assign dfh = ~DFH;  //complement 
assign DIH = ~dih;  //complement 
assign EBQ = DCI & CBC ; 
assign ebq = ~EBQ ; //complement 
assign EDQ = DCI & CBD ; 
assign edq = ~EDQ ;  //complement 
assign EFQ = DCI & CBE ; 
assign efq = ~EFQ ;  //complement 
assign EHQ = DCI & CBF; 
assign ehq = ~EHQ; 
assign EJQ = DFI & CEG ; 
assign ejq = ~EJQ ; //complement 
assign ELQ = DFI & CEH ; 
assign elq = ~ELQ ;  //complement 
assign ENQ = DFI & CEI ; 
assign enq = ~ENQ ;  //complement 
assign EPQ = DFI & CEJ; 
assign epq = ~EPQ; 
assign ERH = DHP & CID ; 
assign erh = ~ERH ; //complement 
assign ETH = DHP & CIE ; 
assign eth = ~ETH ;  //complement 
assign EVH = DHP & CIF ; 
assign evh = ~EVH ;  //complement 
assign dci = ~DCI;  //complement 
assign dfi = ~DFI;  //complement 
assign DII = ~dii;  //complement 
assign EBR = DCJ & CBB ; 
assign ebr = ~EBR ; //complement 
assign EDR = DCJ & CBC ; 
assign edr = ~EDR ;  //complement 
assign EFR = DCJ & CBD ; 
assign efr = ~EFR ;  //complement 
assign EHR = DCJ & CBE; 
assign ehr = ~EHR; 
assign EJR = DFJ & CEF ; 
assign ejr = ~EJR ; //complement 
assign ELR = DFJ & CEG ; 
assign elr = ~ELR ;  //complement 
assign ENR = DFJ & CEH ; 
assign enr = ~ENR ;  //complement 
assign EPR = DFJ & CEI; 
assign epr = ~EPR; 
assign fcl = ~FCL;  //complement 
assign FDL = ~fdl;  //complement 
assign fcm = ~FCM;  //complement 
assign dcj = ~DCJ;  //complement 
assign dfj = ~DFJ;  //complement 
assign DIJ = ~dij;  //complement 
assign ial = ~IAL; //complement 
assign iam = ~IAM; //complement 
assign ian = ~IAN; //complement 
assign iao = ~IAO; //complement 
assign iap = ~IAP; //complement 
assign iba = ~IBA; //complement 
assign ibb = ~IBB; //complement 
assign ibc = ~IBC; //complement 
assign ibd = ~IBD; //complement 
assign ibe = ~IBE; //complement 
assign ibf = ~IBF; //complement 
assign ibg = ~IBG; //complement 
assign ibh = ~IBH; //complement 
assign ibi = ~IBI; //complement 
assign ibj = ~IBJ; //complement 
assign ibk = ~IBK; //complement 
assign ibl = ~IBL; //complement 
assign ibm = ~IBM; //complement 
assign ibn = ~IBN; //complement 
assign ibo = ~IBO; //complement 
assign ibp = ~IBP; //complement 
assign ica = ~ICA; //complement 
assign icb = ~ICB; //complement 
assign icc = ~ICC; //complement 
assign icd = ~ICD; //complement 
assign ice = ~ICE; //complement 
assign icf = ~ICF; //complement 
assign icg = ~ICG; //complement 
assign ich = ~ICH; //complement 
assign ici = ~ICI; //complement 
assign icj = ~ICJ; //complement 
assign ick = ~ICK; //complement 
assign icl = ~ICL; //complement 
assign icm = ~ICM; //complement 
assign icn = ~ICN; //complement 
assign ico = ~ICO; //complement 
assign icp = ~ICP; //complement 
assign idl = ~IDL; //complement 
assign idm = ~IDM; //complement 
assign idn = ~IDN; //complement 
assign ido = ~IDO; //complement 
assign idp = ~IDP; //complement 
assign iea = ~IEA; //complement 
assign ieb = ~IEB; //complement 
assign iec = ~IEC; //complement 
assign ied = ~IED; //complement 
assign iee = ~IEE; //complement 
assign ief = ~IEF; //complement 
assign ieg = ~IEG; //complement 
assign ieh = ~IEH; //complement 
assign iei = ~IEI; //complement 
assign iej = ~IEJ; //complement 
assign iek = ~IEK; //complement 
assign iel = ~IEL; //complement 
assign iem = ~IEM; //complement 
assign ien = ~IEN; //complement 
assign ieo = ~IEO; //complement 
assign iep = ~IEP; //complement 
assign ifa = ~IFA; //complement 
assign ifb = ~IFB; //complement 
assign ifc = ~IFC; //complement 
assign ifd = ~IFD; //complement 
assign ife = ~IFE; //complement 
assign ifff  = ~IFFF ; //complement 
assign ifg = ~IFG; //complement 
assign ifh = ~IFH; //complement 
assign ifi = ~IFI; //complement 
assign ifj = ~IFJ; //complement 
assign ifk = ~IFK; //complement 
assign ifl = ~IFL; //complement 
assign ifm = ~IFM; //complement 
assign ifn = ~IFN; //complement 
assign ifo = ~IFO; //complement 
assign ifp = ~IFP; //complement 
assign iga = ~IGA; //complement 
assign igb = ~IGB; //complement 
assign igc = ~IGC; //complement 
assign igd = ~IGD; //complement 
assign ige = ~IGE; //complement 
assign igf = ~IGF; //complement 
assign igg = ~IGG; //complement 
assign igh = ~IGH; //complement 
assign igi = ~IGI; //complement 
assign igj = ~IGJ; //complement 
assign ila = ~ILA; //complement 
assign ilb = ~ILB; //complement 
assign ilc = ~ILC; //complement 
assign ild = ~ILD; //complement 
assign ile = ~ILE; //complement 
assign ilf = ~ILF; //complement 
assign ilg = ~ILG; //complement 
assign ilh = ~ILH; //complement 
assign ili = ~ILI; //complement 
assign ilj = ~ILJ; //complement 
assign ilk = ~ILK; //complement 
assign ill = ~ILL; //complement 
assign ilm = ~ILM; //complement 
assign ima = ~IMA; //complement 
assign imb = ~IMB; //complement 
assign imc = ~IMC; //complement 
assign imd = ~IMD; //complement 
assign ime = ~IME; //complement 
assign imf = ~IMF; //complement 
assign img = ~IMG; //complement 
assign imh = ~IMH; //complement 
assign imi = ~IMI; //complement 
assign imj = ~IMJ; //complement 
assign imk = ~IMK; //complement 
assign iml = ~IML; //complement 
assign ina = ~INA; //complement 
assign inb = ~INB; //complement 
assign inc = ~INC; //complement 
assign ind = ~IND; //complement 
assign ine = ~INE; //complement 
assign inf = ~INF; //complement 
assign ioa = ~IOA; //complement 
assign iob = ~IOB; //complement 
assign iqc = ~IQC; //complement 
assign iqd = ~IQD; //complement 
assign iqe = ~IQE; //complement 
assign iqf = ~IQF; //complement 
assign iqg = ~IQG; //complement 
assign iqh = ~IQH; //complement 
assign ira = ~IRA; //complement 
assign irb = ~IRB; //complement 
assign irc = ~IRC; //complement 
always@(posedge IZZ )
   begin 
 HAA <=  ILA & ilc & ilk  |  ila & ILC & ilk  |  ila & ilc & ILK  |  ILA & ILC & ILK  ;
 hba <=  ILA & ilc & ilk  |  ila & ILC & ilk  |  ila & ilc & ILK  |  ila & ilc & ilk  ;
 HCC <=  GBC & gcf & gcg  |  gbc & GCF & gcg  |  gbc & gcf & GCG  |  GBC & GCF & GCG  ;
 hdc <=  GBC & gcf & gcg  |  gbc & GCF & gcg  |  gbc & gcf & GCG  |  gbc & gcf & gcg  ;
 HGB <=  GGC & gfd & gge  |  ggc & GFD & gge  |  ggc & gfd & GGE  |  GGC & GFD & GGE  ;
 hhb <=  GGC & gfd & gge  |  ggc & GFD & gge  |  ggc & gfd & GGE  |  ggc & gfd & gge  ;
 MMA <=  LLB & lma & lmb  |  llb & LMA & lmb  |  llb & lma & LMB  |  LLB & LMA & LMB  ;
 mna <=  LLB & lma & lmb  |  llb & LMA & lmb  |  llb & lma & LMB  |  llb & lma & lmb  ;
 MMB <= LLA ; 
 HIE <=  GIE & gig & ghh  |  gie & GIG & ghh  |  gie & gig & GHH  |  GIE & GIG & GHH  ;
 hje <=  GIE & gig & ghh  |  gie & GIG & ghh  |  gie & gig & GHH  |  gie & gig & ghh  ;
 HIG <= FIL ; 
 HMC <=  GLE & gmf & flb  |  gle & GMF & flb  |  gle & gmf & FLB  |  GLE & GMF & FLB  ;
 hnc <=  GLE & gmf & flb  |  gle & GMF & flb  |  gle & gmf & FLB  |  gle & gmf & flb  ;
 OPA <=  MAA & naa & iob  |  maa & NAA & iob  |  maa & naa & IOB  |  MAA & NAA & IOB  ;
 oqa <=  MAA & naa & iob  |  maa & NAA & iob  |  maa & naa & IOB  |  maa & naa & iob  ;
 OPB <= IOA ; 
 KCC <=  JCC & jbb & hcc  |  jcc & JBB & hcc  |  jcc & jbb & HCC  |  JCC & JBB & HCC  ;
 kdc <=  JCC & jbb & hcc  |  jcc & JBB & hcc  |  jcc & jbb & HCC  |  jcc & jbb & hcc  ;
 HQB <=  GQC & gpb & gqb  |  gqc & GPB & gqb  |  gqc & gpb & GQB  |  GQC & GPB & GQB  ;
 hrb <=  GQC & gpb & gqb  |  gqc & GPB & gqb  |  gqc & gpb & GQB  |  gqc & gpb & gqb  ;
 OPS <=  MSA & msb & mra  |  msa & MSB & mra  |  msa & msb & MRA  |  MSA & MSB & MRA  ;
 oqs <=  MSA & msb & mra  |  msa & MSB & mra  |  msa & msb & MRA  |  msa & msb & mra  ;
 KKB <=  JJD & jkc & jjc  |  jjd & JKC & jjc  |  jjd & jkc & JJC  |  JJD & JKC & JJC  ;
 klb <=  JJD & jkc & jjc  |  jjd & JKC & jjc  |  jjd & jkc & JJC  |  jjd & jkc & jjc  ;
 KKD <= HJD ; 
 HUA <=  GTB & gub & gta  |  gtb & GUB & gta  |  gtb & gub & GTA  |  GTB & GUB & GTA  ;
 oha <=  GTB & gub & gta  |  gtb & GUB & gta  |  gtb & gub & GTA  |  gtb & gub & gta  ;
 KSB <=  JRC & jsb & jrb  |  jrc & JSB & jrb  |  jrc & jsb & JRB  |  JRC & JSB & JRB  ;
 ktb <=  JRC & jsb & jrb  |  jrc & JSB & jrb  |  jrc & jsb & JRB  |  jrc & jsb & jrb  ;
 KSC <= JSC ; 
 FQA <=  EQT & equ & eqv  |  eqt & EQU & eqv  |  eqt & equ & EQV  |  EQT & EQU & EQV  ;
 fra <=  EQT & equ & eqv  |  eqt & EQU & eqv  |  eqt & equ & EQV  |  eqt & equ & eqv  ;
 FAA <=  EAL & eam & ean  |  eal & EAM & ean  |  eal & eam & EAN  |  EAL & EAM & EAN  ;
 fba <=  EAL & eam & ean  |  eal & EAM & ean  |  eal & eam & EAN  |  eal & eam & ean  ;
 FAF <=  EAO & eap & eaq  |  eao & EAP & eaq  |  eao & eap & EAQ  |  EAO & EAP & EAQ  ;
 fbf <=  EAO & eap & eaq  |  eao & EAP & eaq  |  eao & eap & EAQ  |  eao & eap & eaq  ;
 FQF <=  EQW & eqx & era  |  eqw & EQX & era  |  eqw & eqx & ERA  |  EQW & EQX & ERA  ;
 frf <=  EQW & eqx & era  |  eqw & EQX & era  |  eqw & eqx & ERA  |  eqw & eqx & era  ;
 FCA <=  EDA & edb & edc  |  eda & EDB & edc  |  eda & edb & EDC  |  EDA & EDB & EDC  ;
 fda <=  EDA & edb & edc  |  eda & EDB & edc  |  eda & edb & EDC  |  eda & edb & edc  ;
 FCE <=  EDD & ede & edf  |  edd & EDE & edf  |  edd & ede & EDF  |  EDD & EDE & EDF  ;
 fde <=  EDD & ede & edf  |  edd & EDE & edf  |  edd & ede & EDF  |  edd & ede & edf  ;
 FSA <=  ESU & esv & esw  |  esu & ESV & esw  |  esu & esv & ESW  |  ESU & ESV & ESW  ;
 fta <=  ESU & esv & esw  |  esu & ESV & esw  |  esu & esv & ESW  |  esu & esv & esw  ;
 FEA <=  EEN & eeo & eep  |  een & EEO & eep  |  een & eeo & EEP  |  EEN & EEO & EEP  ;
 ffa <=  EEN & eeo & eep  |  een & EEO & eep  |  een & eeo & EEP  |  een & eeo & eep  ;
 FEF <=  EEQ & eer & ees  |  eeq & EER & ees  |  eeq & eer & EES  |  EEQ & EER & EES  ;
 fff <=  EEQ & eer & ees  |  eeq & EER & ees  |  eeq & eer & EES  |  eeq & eer & ees  ;
 FSH <=  ETR & ets & ett  |  etr & ETS & ett  |  etr & ets & ETT  |  ETR & ETS & ETT  ;
 fth <=  ETR & ets & ett  |  etr & ETS & ett  |  etr & ets & ETT  |  etr & ets & ett  ;
 FSJ <= ETX ; 
 FGA <=  EGO & egp & egq  |  ego & EGP & egq  |  ego & egp & EGQ  |  EGO & EGP & EGQ  ;
 fha <=  EGO & egp & egq  |  ego & EGP & egq  |  ego & egp & EGQ  |  ego & egp & egq  ;
 FGF <=  EGR & egs & egt  |  egr & EGS & egt  |  egr & egs & EGT  |  EGR & EGS & EGT  ;
 fhf <=  EGR & egs & egt  |  egr & EGS & egt  |  egr & egs & EGT  |  egr & egs & egt  ;
 FUD <=  EVM & evn & evo  |  evm & EVN & evo  |  evm & evn & EVO  |  EVM & EVN & EVO  ;
 ogd <=  EVM & evn & evo  |  evm & EVN & evo  |  evm & evn & EVO  |  evm & evn & evo  ;
 FIA <=  EIP & eiq & eir  |  eip & EIQ & eir  |  eip & eiq & EIR  |  EIP & EIQ & EIR  ;
 fja <=  EIP & eiq & eir  |  eip & EIQ & eir  |  eip & eiq & EIR  |  eip & eiq & eir  ;
 FIF <=  EIS & eit & eiu  |  eis & EIT & eiu  |  eis & eit & EIU  |  EIS & EIT & EIU  ;
 fjf <=  EIS & eit & eiu  |  eis & EIT & eiu  |  eis & eit & EIU  |  eis & eit & eiu  ;
 FKA <=  EKQ & ekr & eks  |  ekq & EKR & eks  |  ekq & ekr & EKS  |  EKQ & EKR & EKS  ;
 fla <=  EKQ & ekr & eks  |  ekq & EKR & eks  |  ekq & ekr & EKS  |  ekq & ekr & eks  ;
 FKF <=  EKT & eku & ekv  |  ekt & EKU & ekv  |  ekt & eku & EKV  |  EKT & EKU & EKV  ;
 flf <=  EKT & eku & ekv  |  ekt & EKU & ekv  |  ekt & eku & EKV  |  ekt & eku & ekv  ;
 FMA <=  EMR & ems & emt  |  emr & EMS & emt  |  emr & ems & EMT  |  EMR & EMS & EMT  ;
 fna <=  EMR & ems & emt  |  emr & EMS & emt  |  emr & ems & EMT  |  emr & ems & emt  ;
 FMF <=  EMU & emv & emw  |  emu & EMV & emw  |  emu & emv & EMW  |  EMU & EMV & EMW  ;
 fnf <=  EMU & emv & emw  |  emu & EMV & emw  |  emu & emv & EMW  |  emu & emv & emw  ;
 FOA <=  EOS & eot & eou  |  eos & EOT & eou  |  eos & eot & EOU  |  EOS & EOT & EOU  ;
 fpa <=  EOS & eot & eou  |  eos & EOT & eou  |  eos & eot & EOU  |  eos & eot & eou  ;
 FOF <=  EOV & eow & eox  |  eov & EOW & eox  |  eov & eow & EOX  |  EOV & EOW & EOX  ;
 fpf <=  EOV & eow & eox  |  eov & EOW & eox  |  eov & eow & EOX  |  eov & eow & eox  ;
 CAL <= IAL ; 
 CAM <= IAM ; 
 CAN <= IAN ; 
 cgn <= ian ; 
 CAO <= IAO ; 
 cgo <= iao ; 
 CAP <= IAP ; 
 CDP <= IAP ; 
 cgp <= iap ; 
 CBA <= IBA ; 
 CEA <= IBA ; 
 cha <= iba ; 
 CBB <= IBB ; 
 CEB <= IBB ; 
 chb <= ibb ; 
 CBC <= IBC ; 
 CEC <= IBC ; 
 chc <= ibc ; 
 CBD <= IBD ; 
 CED <= IBD ; 
 chd <= ibd ; 
 HAB <=  ILG & gaa & ilb  |  ilg & GAA & ilb  |  ilg & gaa & ILB  |  ILG & GAA & ILB  ;
 hbb <=  ILG & gaa & ilb  |  ilg & GAA & ilb  |  ilg & gaa & ILB  |  ilg & gaa & ilb  ;
 HCD <=  GCE & gch & gbd  |  gce & GCH & gbd  |  gce & gch & GBD  |  GCE & GCH & GBD  ;
 hdd <=  GCE & gch & gbd  |  gce & GCH & gbd  |  gce & gch & GBD  |  gce & gch & gbd  ;
 HCE <= FCM ; 
 MAA <=  INA & ind & laa  |  ina & IND & laa  |  ina & ind & LAA  |  INA & IND & LAA  ;
 mba <=  INA & ind & laa  |  ina & IND & laa  |  ina & ind & LAA  |  ina & ind & laa  ;
 MAC <= INB ; 
 HGC <=  GFE & ggd & gfb  |  gfe & GGD & gfb  |  gfe & ggd & GFB  |  GFE & GGD & GFB  ;
 hhc <=  GFE & ggd & gfb  |  gfe & GGD & gfb  |  gfe & ggd & GFB  |  gfe & ggd & gfb  ;
 MOA <=  LOA & lna & lob  |  loa & LNA & lob  |  loa & lna & LOB  |  LOA & LNA & LOB  ;
 mpa <=  LOA & lna & lob  |  loa & LNA & lob  |  loa & lna & LOB  |  loa & lna & lob  ;
 MOB <= LNB ; 
 HKA <=  GKA & gjb & gkb  |  gka & GJB & gkb  |  gka & gjb & GKB  |  GKA & GJB & GKB  ;
 hla <=  GKA & gjb & gkb  |  gka & GJB & gkb  |  gka & gjb & GKB  |  gka & gjb & gkb  ;
 HMD <=  GMC & gmd & gld  |  gmc & GMD & gld  |  gmc & gmd & GLD  |  GMC & GMD & GLD  ;
 hnd <=  GMC & gmd & gld  |  gmc & GMD & gld  |  gmc & gmd & GLD  |  gmc & gmd & gld  ;
 OPC <=  MCC & mbb & nba  |  mcc & MBB & nba  |  mcc & mbb & NBA  |  MCC & MBB & NBA  ;
 oqc <=  MCC & mbb & nba  |  mcc & MBB & nba  |  mcc & mbb & NBA  |  mcc & mbb & nba  ;
 OPD <= NCA ; 
 KEA <=  JEA & jda & hea  |  jea & JDA & hea  |  jea & jda & HEA  |  JEA & JDA & HEA  ;
 kfa <=  JEA & jda & hea  |  jea & JDA & hea  |  jea & jda & HEA  |  jea & jda & hea  ;
 HQC <=  GPD & gpe & fpe  |  gpd & GPE & fpe  |  gpd & gpe & FPE  |  GPD & GPE & FPE  ;
 hrc <=  GPD & gpe & fpe  |  gpd & GPE & fpe  |  gpd & gpe & FPE  |  gpd & gpe & fpe  ;
 OPU <=  MTA & mua & mub  |  mta & MUA & mub  |  mta & mua & MUB  |  MTA & MUA & MUB  ;
 oqu <=  MTA & mua & mub  |  mta & MUA & mub  |  mta & mua & MUB  |  mta & mua & mub  ;
 KMA <=  JLA & jma & jlb  |  jla & JMA & jlb  |  jla & jma & JLB  |  JLA & JMA & JLB  ;
 kna <=  JLA & jma & jlb  |  jla & JMA & jlb  |  jla & jma & JLB  |  jla & jma & jlb  ;
 KMC <= JLC ; 
 HUB <=  GTC & guc & gue  |  gtc & GUC & gue  |  gtc & guc & GUE  |  GTC & GUC & GUE  ;
 ohb <=  GTC & guc & gue  |  gtc & GUC & gue  |  gtc & guc & GUE  |  gtc & guc & gue  ;
 KUA <=  HTA & jta & jua  |  hta & JTA & jua  |  hta & jta & JUA  |  HTA & JTA & JUA  ;
 oka <=  HTA & jta & jua  |  hta & JTA & jua  |  hta & jta & JUA  |  hta & jta & jua  ;
 FQB <=  ERH & eri & erj  |  erh & ERI & erj  |  erh & eri & ERJ  |  ERH & ERI & ERJ  ;
 frb <=  ERH & eri & erj  |  erh & ERI & erj  |  erh & eri & ERJ  |  erh & eri & erj  ;
 FAB <=  EAX & eba & ebb  |  eax & EBA & ebb  |  eax & eba & EBB  |  EAX & EBA & EBB  ;
 fbb <=  EAX & eba & ebb  |  eax & EBA & ebb  |  eax & eba & EBB  |  eax & eba & ebb  ;
 FAG <=  EAR & eas & eat  |  ear & EAS & eat  |  ear & eas & EAT  |  EAR & EAS & EAT  ;
 fbg <=  EAR & eas & eat  |  ear & EAS & eat  |  ear & eas & EAT  |  ear & eas & eat  ;
 FQG <=  ERB & erc & erd  |  erb & ERC & erd  |  erb & erc & ERD  |  ERB & ERC & ERD  ;
 frg <=  ERB & erc & erd  |  erb & ERC & erd  |  erb & erc & ERD  |  erb & erc & erd  ;
 FCB <=  ECM & ecn & eco  |  ecm & ECN & eco  |  ecm & ecn & ECO  |  ECM & ECN & ECO  ;
 fdb <=  ECM & ecn & eco  |  ecm & ECN & eco  |  ecm & ecn & ECO  |  ecm & ecn & eco  ;
 FCF <=  ECP & ecq & ecr  |  ecp & ECQ & ecr  |  ecp & ecq & ECR  |  ECP & ECQ & ECR  ;
 fdf <=  ECP & ecq & ecr  |  ecp & ECQ & ecr  |  ecp & ecq & ECR  |  ecp & ecq & ecr  ;
 FSB <=  ETI & etj & etk  |  eti & ETJ & etk  |  eti & etj & ETK  |  ETI & ETJ & ETK  ;
 ftb <=  ETI & etj & etk  |  eti & ETJ & etk  |  eti & etj & ETK  |  eti & etj & etk  ;
 FEB <=  EFB & efc & efd  |  efb & EFC & efd  |  efb & efc & EFD  |  EFB & EFC & EFD  ;
 ffb <=  EFB & efc & efd  |  efb & EFC & efd  |  efb & efc & EFD  |  efb & efc & efd  ;
 FEG <=  EET & eeu & eev  |  eet & EEU & eev  |  eet & eeu & EEV  |  EET & EEU & EEV  ;
 ffg <=  EET & eeu & eev  |  eet & EEU & eev  |  eet & eeu & EEV  |  eet & eeu & eev  ;
 FSI <=  ETF & etg & eth  |  etf & ETG & eth  |  etf & etg & ETH  |  ETF & ETG & ETH  ;
 fti <=  ETF & etg & eth  |  etf & ETG & eth  |  etf & etg & ETH  |  etf & etg & eth  ;
 FSK <= QIC ; 
 FGB <=  EHC & ehd & ehe  |  ehc & EHD & ehe  |  ehc & ehd & EHE  |  EHC & EHD & EHE  ;
 fhb <=  EHC & ehd & ehe  |  ehc & EHD & ehe  |  ehc & ehd & EHE  |  ehc & ehd & ehe  ;
 FGG <=  EGU & egv & egw  |  egu & EGV & egw  |  egu & egv & EGW  |  EGU & EGV & EGW  ;
 fhg <=  EGU & egv & egw  |  egu & EGV & egw  |  egu & egv & EGW  |  egu & egv & egw  ;
 FUE <=  EVA & evb & evc  |  eva & EVB & evc  |  eva & evb & EVC  |  EVA & EVB & EVC  ;
 oge <=  EVA & evb & evc  |  eva & EVB & evc  |  eva & evb & EVC  |  eva & evb & evc  ;
 FIB <=  EJD & eje & ejf  |  ejd & EJE & ejf  |  ejd & eje & EJF  |  EJD & EJE & EJF  ;
 fjb <=  EJD & eje & ejf  |  ejd & EJE & ejf  |  ejd & eje & EJF  |  ejd & eje & ejf  ;
 FIG <=  EIV & eiw & eix  |  eiv & EIW & eix  |  eiv & eiw & EIX  |  EIV & EIW & EIX  ;
 fjg <=  EIV & eiw & eix  |  eiv & EIW & eix  |  eiv & eiw & EIX  |  eiv & eiw & eix  ;
 FKB <=  ELE & elf & elg  |  ele & ELF & elg  |  ele & elf & ELG  |  ELE & ELF & ELG  ;
 flb <=  ELE & elf & elg  |  ele & ELF & elg  |  ele & elf & ELG  |  ele & elf & elg  ;
 FKG <=  EKW & ekx & ela  |  ekw & EKX & ela  |  ekw & ekx & ELA  |  EKW & EKX & ELA  ;
 flg <=  EKW & ekx & ela  |  ekw & EKX & ela  |  ekw & ekx & ELA  |  ekw & ekx & ela  ;
 FMB <=  ENR & ens & ent  |  enr & ENS & ent  |  enr & ens & ENT  |  ENR & ENS & ENT  ;
 fnb <=  ENR & ens & ent  |  enr & ENS & ent  |  enr & ens & ENT  |  enr & ens & ent  ;
 FMG <=  EMX & ena & enb  |  emx & ENA & enb  |  emx & ena & ENB  |  EMX & ENA & ENB  ;
 fng <=  EMX & ena & enb  |  emx & ENA & enb  |  emx & ena & ENB  |  emx & ena & enb  ;
 FOB <=  EPG & eph & epi  |  epg & EPH & epi  |  epg & eph & EPI  |  EPG & EPH & EPI  ;
 fpb <=  EPG & eph & epi  |  epg & EPH & epi  |  epg & eph & EPI  |  epg & eph & epi  ;
 FOG <=  EPA & epb & epc  |  epa & EPB & epc  |  epa & epb & EPC  |  EPA & EPB & EPC  ;
 fpg <=  EPA & epb & epc  |  epa & EPB & epc  |  epa & epb & EPC  |  epa & epb & epc  ;
 CBE <= IBE ; 
 CEE <= IBE ; 
 che <= ibe ; 
 chl <= ibl ; 
 CBF <= IBF ; 
 CEF <= IBF ; 
 chf <= ibf ; 
 ckl <= ibl ; 
 CBG <= IGA & TAA |  IBG & taa ; 
 CEG <= IGA & TAA |  IBG & taa ; 
 chg <= ibg ; 
 chh <= ibh ; 
 CBH <= IGB & TAA |  IBH & taa ; 
 CEH <= IGB & TAA |  IBH & taa ; 
 TAA <= QJA ; 
 TAB <= QJA ; 
 CBI <= IGC & TAA |  IBI & taa ; 
 CEI <= IGC & TAA |  IBI & taa ; 
 QIC <= IQC ; 
 QID <= IQD ; 
 QIE <= IQE ; 
 QIF <= IQF ; 
 QIG <= IQG ; 
 QIH <= IQH ; 
 chi <= ibi ; 
 cki <= ibi ; 
 chj <= ibj ; 
 ckj <= ibj ; 
 CBJ <= IGD & TAA |  IBJ & taa ; 
 CEJ <= IGD & TAA |  IBJ & taa ; 
 CBK <= TAA & IGE ; 
 CEK <= TAA & IGE ; 
 chk <= TAA & ibk ; 
 ckk <= TAA & ibk ; 
 CBL <= IGF & TAB |  IBL & tab ; 
 CEL <= IGF & TAB |  IBL & tab ; 
 HAC <=  ILL & ild & ilh  |  ill & ILD & ilh  |  ill & ild & ILH  |  ILL & ILD & ILH  ;
 hbc <=  ILL & ild & ilh  |  ill & ILD & ilh  |  ill & ild & ILH  |  ill & ild & ilh  ;
 HEA <=  GEA & gda & gdb  |  gea & GDA & gdb  |  gea & gda & GDB  |  GEA & GDA & GDB  ;
 hfa <=  GEA & gda & gdb  |  gea & GDA & gdb  |  gea & gda & GDB  |  gea & gda & gdb  ;
 MAB <=  KAC & kad & inc  |  kac & KAD & inc  |  kac & kad & INC  |  KAC & KAD & INC  ;
 mbb <=  KAC & kad & inc  |  kac & KAD & inc  |  kac & kad & INC  |  kac & kad & inc  ;
 MAD <= INE ; 
 HGD <=  GGH & gfg & gff  |  ggh & GFG & gff  |  ggh & gfg & GFF  |  GGH & GFG & GFF  ;
 hhd <=  GGH & gfg & gff  |  ggh & GFG & gff  |  ggh & gfg & GFF  |  ggh & gfg & gff  ;
 HGF <= GFC ; 
 HKB <=  FJD & gja & gjc  |  fjd & GJA & gjc  |  fjd & gja & GJC  |  FJD & GJA & GJC  ;
 hlb <=  FJD & gja & gjc  |  fjd & GJA & gjc  |  fjd & gja & GJC  |  fjd & gja & gjc  ;
 KAA <=  IMA & jaa & img  |  ima & JAA & img  |  ima & jaa & IMG  |  IMA & JAA & IMG  ;
 kba <=  IMA & jaa & img  |  ima & JAA & img  |  ima & jaa & IMG  |  ima & jaa & img  ;
 HME <=  GLF & gmg & glg  |  glf & GMG & glg  |  glf & gmg & GLG  |  GLF & GMG & GLG  ;
 hne <=  GLF & gmg & glg  |  glf & GMG & glg  |  glf & gmg & GLG  |  glf & gmg & glg  ;
 HMF <= GME ; 
 OPG <=  NFA & mgb & nga  |  nfa & MGB & nga  |  nfa & mgb & NGA  |  NFA & MGB & NGA  ;
 oqg <=  NFA & mgb & nga  |  nfa & MGB & nga  |  nfa & mgb & NGA  |  nfa & mgb & nga  ;
 KEB <=  JDB & jdc & jec  |  jdb & JDC & jec  |  jdb & jdc & JEC  |  JDB & JDC & JEC  ;
 kfb <=  JDB & jdc & jec  |  jdb & JDC & jec  |  jdb & jdc & JEC  |  jdb & jdc & jec  ;
 KEC <= JEB ; 
 HQD <=  GQD & gqe & gpg  |  gqd & GQE & gpg  |  gqd & gqe & GPG  |  GQD & GQE & GPG  ;
 hrd <=  GQD & gqe & gpg  |  gqd & GQE & gpg  |  gqd & gqe & GPG  |  gqd & gqe & gpg  ;
 KMB <=  JMB & hlc & hmc  |  jmb & HLC & hmc  |  jmb & hlc & HMC  |  JMB & HLC & HMC  ;
 knb <=  JMB & hlc & hmc  |  jmb & HLC & hmc  |  jmb & hlc & HMC  |  jmb & hlc & hmc  ;
 KMD <= JMC ; 
 HUC <=  GTD & gud & gte  |  gtd & GUD & gte  |  gtd & gud & GTE  |  GTD & GUD & GTE  ;
 ohc <=  GTD & gud & gte  |  gtd & GUD & gte  |  gtd & gud & GTE  |  gtd & gud & gte  ;
 HUE <= GUA ; 
 KUB <=  JTB & juc & jtc  |  jtb & JUC & jtc  |  jtb & juc & JTC  |  JTB & JUC & JTC  ;
 okb <=  JTB & juc & jtc  |  jtb & JUC & jtc  |  jtb & juc & JTC  |  jtb & juc & jtc  ;
 KUC <= JUB ; 
 FAC <=  EBL & ebm & ebn  |  ebl & EBM & ebn  |  ebl & ebm & EBN  |  EBL & EBM & EBN  ;
 fbc <=  EBL & ebm & ebn  |  ebl & EBM & ebn  |  ebl & ebm & EBN  |  ebl & ebm & ebn  ;
 FAH <=  EBF & ebg & ebh  |  ebf & EBG & ebh  |  ebf & ebg & EBH  |  EBF & EBG & EBH  ;
 fbh <=  EBF & ebg & ebh  |  ebf & EBG & ebh  |  ebf & ebg & EBH  |  ebf & ebg & ebh  ;
 FCG <=  ECS & ect & ecu  |  ecs & ECT & ecu  |  ecs & ect & ECU  |  ECS & ECT & ECU  ;
 fdg <=  ECS & ect & ecu  |  ecs & ECT & ecu  |  ecs & ect & ECU  |  ecs & ect & ecu  ;
 CBM <= IGG & TAB |  IBM & tab ; 
 CEM <= IGG & TAB |  IBM & tab ; 
 chm <= ibm ; 
 ckm <= ibm ; 
 CBN <= IGH & TAB |  IBN & tab ; 
 CEN <= IGH & TAB |  IBN & tab ; 
 chn <= ibn ; 
 ckn <= ibn ; 
 CBO <= TAB & IGI ; 
 CEO <= TAB & IGI ; 
 cho <= TAB & ibo ; 
 cko <= TAB & ibo ; 
 CBP <= IGJ & TAB |  IBP & tab ; 
 CEP <= IGJ & TAB |  IBP & tab ; 
 chp <= ibp ; 
 ckp <= ibp ; 
 CCA <= ICA ; 
 CFA <= ICA ; 
 cia <= ica ; 
 cla <= ica ; 
 CCB <= ICB ; 
 CFB <= ICB ; 
 cib <= icb ; 
 clb <= icb ; 
 CCC <= ICC ; 
 CFC <= ICC ; 
 cic <= icc ; 
 clc <= icc ; 
 QJA <= IRA ; 
 QJB <= IRB ; 
 QJC <= IRC ; 
 CCD <= ICD ; 
 CFD <= ICD ; 
 cid <= icd ; 
 cld <= icd ; 
 HAD <=  GAC & ilm & ile  |  gac & ILM & ile  |  gac & ilm & ILE  |  GAC & ILM & ILE  ;
 hbd <=  GAC & ilm & ile  |  gac & ILM & ile  |  gac & ilm & ILE  |  gac & ilm & ile  ;
 HEB <=  GDC & gec & geb  |  gdc & GEC & geb  |  gdc & gec & GEB  |  GDC & GEC & GEB  ;
 hfb <=  GDC & gec & geb  |  gdc & GEC & geb  |  gdc & gec & GEB  |  gdc & gec & geb  ;
 MCA <=  LCA & lba & lcb  |  lca & LBA & lcb  |  lca & lba & LCB  |  LCA & LBA & LCB  ;
 mda <=  LCA & lba & lcb  |  lca & LBA & lcb  |  lca & lba & LCB  |  lca & lba & lcb  ;
 MCB <= INF ; 
 HGE <=  GFH & ggg & ggf  |  gfh & GGG & ggf  |  gfh & ggg & GGF  |  GFH & GGG & GGF  ;
 hhe <=  GFH & ggg & ggf  |  gfh & GGG & ggf  |  gfh & ggg & GGF  |  gfh & ggg & ggf  ;
 HGG <= FGM ; 
 MQA <=  KQA & lpa & lpb  |  kqa & LPA & lpb  |  kqa & lpa & LPB  |  KQA & LPA & LPB  ;
 mra <=  KQA & lpa & lpb  |  kqa & LPA & lpb  |  kqa & lpa & LPB  |  kqa & lpa & lpb  ;
 MQB <= LQA ; 
 HKC <=  GKC & gje & gjd  |  gkc & GJE & gjd  |  gkc & gje & GJD  |  GKC & GJE & GJD  ;
 hlc <=  GKC & gje & gjd  |  gkc & GJE & gjd  |  gkc & gje & GJD  |  gkc & gje & gjd  ;
 MGC <= LGA ; 
 MCC <= KCC ; 
 OPE <= NDA ; 
 OPF <= NEA ; 
 KAB <=  IMD & imc & imj  |  imd & IMC & imj  |  imd & imc & IMJ  |  IMD & IMC & IMJ  ;
 kbb <=  IMD & imc & imj  |  imd & IMC & imj  |  imd & imc & IMJ  |  imd & imc & imj  ;
 HOA <=  GOB & gna & goa  |  gob & GNA & goa  |  gob & gna & GOA  |  GOB & GNA & GOA  ;
 hpa <=  GOB & gna & goa  |  gob & GNA & goa  |  gob & gna & GOA  |  gob & gna & goa  ;
 OPI <=  MIA & nha & mha  |  mia & NHA & mha  |  mia & nha & MHA  |  MIA & NHA & MHA  ;
 oqi <=  MIA & nha & mha  |  mia & NHA & mha  |  mia & nha & MHA  |  mia & nha & mha  ;
 KGA <=  JGA & jfb & jgb  |  jga & JFB & jgb  |  jga & jfb & JGB  |  JGA & JFB & JGB  ;
 kha <=  JGA & jfb & jgb  |  jga & JFB & jgb  |  jga & jfb & JGB  |  jga & jfb & jgb  ;
 HQE <=  FPB & gpf & gqf  |  fpb & GPF & gqf  |  fpb & gpf & GQF  |  FPB & GPF & GQF  ;
 hre <=  FPB & gpf & gqf  |  fpb & GPF & gqf  |  fpb & gpf & GQF  |  fpb & gpf & gqf  ;
 KOA <=  JOA & jna & job  |  joa & JNA & job  |  joa & jna & JOB  |  JOA & JNA & JOB  ;
 kpa <=  JOA & jna & job  |  joa & JNA & job  |  joa & jna & JOB  |  joa & jna & job  ;
 KOC <= HNC ; 
 HUD <=  GTF & gtg & guf  |  gtf & GTG & guf  |  gtf & gtg & GUF  |  GTF & GTG & GUF  ;
 ohd <=  GTF & gtg & guf  |  gtf & GTG & guf  |  gtf & gtg & GUF  |  gtf & gtg & guf  ;
 HUF <= FTE ; 
 FQC <=  ERT & eru & erv  |  ert & ERU & erv  |  ert & eru & ERV  |  ERT & ERU & ERV  ;
 frc <=  ERT & eru & erv  |  ert & ERU & erv  |  ert & eru & ERV  |  ert & eru & erv  ;
 FAD <=  EBO & ebp & ebq  |  ebo & EBP & ebq  |  ebo & ebp & EBQ  |  EBO & EBP & EBQ  ;
 fbd <=  EBO & ebp & ebq  |  ebo & EBP & ebq  |  ebo & ebp & EBQ  |  ebo & ebp & ebq  ;
 FAI <=  EBR & ebs & ebt  |  ebr & EBS & ebt  |  ebr & ebs & EBT  |  EBR & EBS & EBT  ;
 fbi <=  EBR & ebs & ebt  |  ebr & EBS & ebt  |  ebr & ebs & EBT  |  ebr & ebs & ebt  ;
 FQH <=  ERN & ero & erp  |  ern & ERO & erp  |  ern & ero & ERP  |  ERN & ERO & ERP  ;
 frh <=  ERN & ero & erp  |  ern & ERO & erp  |  ern & ero & ERP  |  ern & ero & erp  ;
 FCC <=  EDM & edn & edo  |  edm & EDN & edo  |  edm & edn & EDO  |  EDM & EDN & EDO  ;
 fdc <=  EDM & edn & edo  |  edm & EDN & edo  |  edm & edn & EDO  |  edm & edn & edo  ;
 FCH <=  EDG & edh & edi  |  edg & EDH & edi  |  edg & edh & EDI  |  EDG & EDH & EDI  ;
 fdh <=  EDG & edh & edi  |  edg & EDH & edi  |  edg & edh & EDI  |  edg & edh & edi  ;
 FSC <=  ETU & etv & etw  |  etu & ETV & etw  |  etu & etv & ETW  |  ETU & ETV & ETW  ;
 ftc <=  ETU & etv & etw  |  etu & ETV & etw  |  etu & etv & ETW  |  etu & etv & etw  ;
 FEC <=  EFN & efo & efp  |  efn & EFO & efp  |  efn & efo & EFP  |  EFN & EFO & EFP  ;
 ffc <=  EFN & efo & efp  |  efn & EFO & efp  |  efn & efo & EFP  |  efn & efo & efp  ;
 FEH <=  EFH & efi & efj  |  efh & EFI & efj  |  efh & efi & EFJ  |  EFH & EFI & EFJ  ;
 ffh <=  EFH & efi & efj  |  efh & EFI & efj  |  efh & efi & EFJ  |  efh & efi & efj  ;
 FUA <=  EUV & euw & eux  |  euv & EUW & eux  |  euv & euw & EUX  |  EUV & EUW & EUX  ;
 oga <=  EUV & euw & eux  |  euv & EUW & eux  |  euv & euw & EUX  |  euv & euw & eux  ;
 FGC <=  EHO & ehp & ehq  |  eho & EHP & ehq  |  eho & ehp & EHQ  |  EHO & EHP & EHQ  ;
 fhc <=  EHO & ehp & ehq  |  eho & EHP & ehq  |  eho & ehp & EHQ  |  eho & ehp & ehq  ;
 FGH <=  EHI & ehj & ehk  |  ehi & EHJ & ehk  |  ehi & ehj & EHK  |  EHI & EHJ & EHK  ;
 fhh <=  EHI & ehj & ehk  |  ehi & EHJ & ehk  |  ehi & ehj & EHK  |  ehi & ehj & ehk  ;
 FUF <=  EVD & eve & evf  |  evd & EVE & evf  |  evd & eve & EVF  |  EVD & EVE & EVF  ;
 ogf <=  EVD & eve & evf  |  evd & EVE & evf  |  evd & eve & EVF  |  evd & eve & evf  ;
 FIC <=  EJP & ejq & ejr  |  ejp & EJQ & ejr  |  ejp & ejq & EJR  |  EJP & EJQ & EJR  ;
 fjc <=  EJP & ejq & ejr  |  ejp & EJQ & ejr  |  ejp & ejq & EJR  |  ejp & ejq & ejr  ;
 FIH <=  EJJ & ejk & ejl  |  ejj & EJK & ejl  |  ejj & ejk & EJL  |  EJJ & EJK & EJL  ;
 fjh <=  EJJ & ejk & ejl  |  ejj & EJK & ejl  |  ejj & ejk & EJL  |  ejj & ejk & ejl  ;
 FKC <=  ELQ & elr & els  |  elq & ELR & els  |  elq & elr & ELS  |  ELQ & ELR & ELS  ;
 flc <=  ELQ & elr & els  |  elq & ELR & els  |  elq & elr & ELS  |  elq & elr & els  ;
 FKH <=  ELK & ell & elm  |  elk & ELL & elm  |  elk & ell & ELM  |  ELK & ELL & ELM  ;
 flh <=  ELK & ell & elm  |  elk & ELL & elm  |  elk & ell & ELM  |  elk & ell & elm  ;
 FMC <=  ENF & eng & enh  |  enf & ENG & enh  |  enf & eng & ENH  |  ENF & ENG & ENH  ;
 fnc <=  ENF & eng & enh  |  enf & ENG & enh  |  enf & eng & ENH  |  enf & eng & enh  ;
 FMH <=  ENL & enm & enn  |  enl & ENM & enn  |  enl & enm & ENN  |  ENL & ENM & ENN  ;
 fnh <=  ENL & enm & enn  |  enl & ENM & enn  |  enl & enm & ENN  |  enl & enm & enn  ;
 FOC <=  EPS & ept & epu  |  eps & EPT & epu  |  eps & ept & EPU  |  EPS & EPT & EPU  ;
 fpc <=  EPS & ept & epu  |  eps & EPT & epu  |  eps & ept & EPU  |  eps & ept & epu  ;
 FOH <=  EPM & epn & epo  |  epm & EPN & epo  |  epm & epn & EPO  |  EPM & EPN & EPO  ;
 fph <=  EPM & epn & epo  |  epm & EPN & epo  |  epm & epn & EPO  |  epm & epn & epo  ;
 CCE <= ICE ; 
 CFE <= ICE ; 
 cie <= ice ; 
 CCF <= ICF ; 
 CFF <= ICF ; 
 cif <= icf ; 
 CCG <= ICG ; 
 CFG <= ICG ; 
 cig <= icg ; 
 CCH <= ICH ; 
 CFH <= ICH ; 
 cih <= ich ; 
 CCI <= ICI ; 
 CFI <= ICI ; 
 cii <= ici ; 
 CCJ <= ICJ ; 
 CFJ <= ICJ ; 
 cij <= icj ; 
 CCK <= ICK ; 
 CFK <= ICK ; 
 cik <= ick ; 
 CCL <= ICL ; 
 CFL <= ICL ; 
 cil <= icl ; 
 HAE <=  GAB & fam & fan  |  gab & FAM & fan  |  gab & fam & FAN  |  GAB & FAM & FAN  ;
 hbe <=  GAB & fam & fan  |  gab & FAM & fan  |  gab & fam & FAN  |  gab & fam & fan  ;
 HEC <=  GDD & ged & gee  |  gdd & GED & gee  |  gdd & ged & GEE  |  GDD & GED & GEE  ;
 hfc <=  GDD & ged & gee  |  gdd & GED & gee  |  gdd & ged & GEE  |  gdd & ged & gee  ;
 MEA <=  LDA & ldb & leb  |  lda & LDB & leb  |  lda & ldb & LEB  |  LDA & LDB & LEB  ;
 mfa <=  LDA & ldb & leb  |  lda & LDB & leb  |  lda & ldb & LEB  |  lda & ldb & leb  ;
 MEB <= LEA ; 
 HIA <=  GHA & gib & gia  |  gha & GIB & gia  |  gha & gib & GIA  |  GHA & GIB & GIA  ;
 hja <=  GHA & gib & gia  |  gha & GIB & gia  |  gha & gib & GIA  |  gha & gib & gia  ;
 MSA <=  LRA & lsa & ksa  |  lra & LSA & ksa  |  lra & lsa & KSA  |  LRA & LSA & KSA  ;
 mta <=  LRA & lsa & ksa  |  lra & LSA & ksa  |  lra & lsa & KSA  |  lra & lsa & ksa  ;
 MSB <= KRA ; 
 HKD <=  GKD & gkf & gjf  |  gkd & GKF & gjf  |  gkd & gkf & GJF  |  GKD & GKF & GJF  ;
 hld <=  GKD & gkf & gjf  |  gkd & GKF & gjf  |  gkd & gkf & GJF  |  gkd & gkf & gjf  ;
 OMB <= LVA ; 
 KAC <=  IME & imi & imh  |  ime & IMI & imh  |  ime & imi & IMH  |  IME & IMI & IMH  ;
 kbc <=  IME & imi & imh  |  ime & IMI & imh  |  ime & imi & IMH  |  ime & imi & imh  ;
 HOB <=  GNC & gnd & goc  |  gnc & GND & goc  |  gnc & gnd & GOC  |  GNC & GND & GOC  ;
 hpb <=  GNC & gnd & goc  |  gnc & GND & goc  |  gnc & gnd & GOC  |  gnc & gnd & goc  ;
 OPK <=  MKA & mkb & mja  |  mka & MKB & mja  |  mka & mkb & MJA  |  MKA & MKB & MJA  ;
 oqk <=  MKA & mkb & mja  |  mka & MKB & mja  |  mka & mkb & MJA  |  mka & mkb & mja  ;
 KGB <=  JGC & jfc & jgd  |  jgc & JFC & jgd  |  jgc & jfc & JGD  |  JGC & JFC & JGD  ;
 khb <=  JGC & jfc & jgd  |  jgc & JFC & jgd  |  jgc & jfc & JGD  |  jgc & jfc & jgd  ;
 KGC <= JFA ; 
 HSA <=  GRA & gsa & gsb  |  gra & GSA & gsb  |  gra & gsa & GSB  |  GRA & GSA & GSB  ;
 hta <=  GRA & gsa & gsb  |  gra & GSA & gsb  |  gra & gsa & GSB  |  gra & gsa & gsb  ;
 KOB <=  JNC & joc & hoc  |  jnc & JOC & hoc  |  jnc & joc & HOC  |  JNC & JOC & HOC  ;
 kpb <=  JNC & joc & hoc  |  jnc & JOC & hoc  |  jnc & joc & HOC  |  jnc & joc & hoc  ;
 KOD <= JNB ; 
 FQD <=  ERW & erx & qif  |  erw & ERX & qif  |  erw & erx & QIF  |  ERW & ERX & QIF  ;
 frd <=  ERW & erx & qif  |  erw & ERX & qif  |  erw & erx & QIF  |  erw & erx & qif  ;
 FAE <=  EBC & ebd & ebe  |  ebc & EBD & ebe  |  ebc & ebd & EBE  |  EBC & EBD & EBE  ;
 fbe <=  EBC & ebd & ebe  |  ebc & EBD & ebe  |  ebc & ebd & EBE  |  ebc & ebd & ebe  ;
 FAJ <=  EBU & ebv & ebw  |  ebu & EBV & ebw  |  ebu & ebv & EBW  |  EBU & EBV & EBW  ;
 fbj <=  EBU & ebv & ebw  |  ebu & EBV & ebw  |  ebu & ebv & EBW  |  ebu & ebv & ebw  ;
 FAM <= EBX ; 
 FQI <=  ERQ & err & ers  |  erq & ERR & ers  |  erq & err & ERS  |  ERQ & ERR & ERS  ;
 fri <=  ERQ & err & ers  |  erq & ERR & ers  |  erq & err & ERS  |  erq & err & ers  ;
 FCD <=  EDP & edq & edr  |  edp & EDQ & edr  |  edp & edq & EDR  |  EDP & EDQ & EDR  ;
 fdd <=  EDP & edq & edr  |  edp & EDQ & edr  |  edp & edq & EDR  |  edp & edq & edr  ;
 FCI <=  EDS & edt & edu  |  eds & EDT & edu  |  eds & edt & EDU  |  EDS & EDT & EDU  ;
 fdi <=  EDS & edt & edu  |  eds & EDT & edu  |  eds & edt & EDU  |  eds & edt & edu  ;
 FSD <=  ETL & etm & etn  |  etl & ETM & etn  |  etl & etm & ETN  |  ETL & ETM & ETN  ;
 ftd <=  ETL & etm & etn  |  etl & ETM & etn  |  etl & etm & ETN  |  etl & etm & etn  ;
 FED <=  EFQ & efr & efs  |  efq & EFR & efs  |  efq & efr & EFS  |  EFQ & EFR & EFS  ;
 ffd <=  EFQ & efr & efs  |  efq & EFR & efs  |  efq & efr & EFS  |  efq & efr & efs  ;
 FEI <=  EFT & efu & efv  |  eft & EFU & efv  |  eft & efu & EFV  |  EFT & EFU & EFV  ;
 ffi <=  EFT & efu & efv  |  eft & EFU & efv  |  eft & efu & EFV  |  eft & efu & efv  ;
 FUB <=  EVJ & evk & evl  |  evj & EVK & evl  |  evj & evk & EVL  |  EVJ & EVK & EVL  ;
 ogb <=  EVJ & evk & evl  |  evj & EVK & evl  |  evj & evk & EVL  |  evj & evk & evl  ;
 FGD <=  EHR & ehs & eht  |  ehr & EHS & eht  |  ehr & ehs & EHT  |  EHR & EHS & EHT  ;
 fhd <=  EHR & ehs & eht  |  ehr & EHS & eht  |  ehr & ehs & EHT  |  ehr & ehs & eht  ;
 FGI <=  EHU & ehv & ehw  |  ehu & EHV & ehw  |  ehu & ehv & EHW  |  EHU & EHV & EHW  ;
 fhi <=  EHU & ehv & ehw  |  ehu & EHV & ehw  |  ehu & ehv & EHW  |  ehu & ehv & ehw  ;
 FUG <=  EVP & evq & evr  |  evp & EVQ & evr  |  evp & evq & EVR  |  EVP & EVQ & EVR  ;
 ogg <=  EVP & evq & evr  |  evp & EVQ & evr  |  evp & evq & EVR  |  evp & evq & evr  ;
 FID <=  EJS & ejt & eju  |  ejs & EJT & eju  |  ejs & ejt & EJU  |  EJS & EJT & EJU  ;
 fjd <=  EJS & ejt & eju  |  ejs & EJT & eju  |  ejs & ejt & EJU  |  ejs & ejt & eju  ;
 FII <=  EJV & ejw & ejx  |  ejv & EJW & ejx  |  ejv & ejw & EJX  |  EJV & EJW & EJX  ;
 fji <=  EJV & ejw & ejx  |  ejv & EJW & ejx  |  ejv & ejw & EJX  |  ejv & ejw & ejx  ;
 FKD <=  ELT & elu & elv  |  elt & ELU & elv  |  elt & elu & ELV  |  ELT & ELU & ELV  ;
 fld <=  ELT & elu & elv  |  elt & ELU & elv  |  elt & elu & ELV  |  elt & elu & elv  ;
 FKI <=  ELW & elx & qie  |  elw & ELX & qie  |  elw & elx & QIE  |  ELW & ELX & QIE  ;
 fli <=  ELW & elx & qie  |  elw & ELX & qie  |  elw & elx & QIE  |  elw & elx & qie  ;
 FMD <=  ENU & env & enw  |  enu & ENV & enw  |  enu & env & ENW  |  ENU & ENV & ENW  ;
 fnd <=  ENU & env & enw  |  enu & ENV & enw  |  enu & env & ENW  |  enu & env & enw  ;
 FMI <=  ENO & enp & enq  |  eno & ENP & enq  |  eno & enp & ENQ  |  ENO & ENP & ENQ  ;
 fni <=  ENO & enp & enq  |  eno & ENP & enq  |  eno & enp & ENQ  |  eno & enp & enq  ;
 FMK <= ENX ; 
 FOD <=  EPV & epw & epx  |  epv & EPW & epx  |  epv & epw & EPX  |  EPV & EPW & EPX  ;
 fpd <=  EPV & epw & epx  |  epv & EPW & epx  |  epv & epw & EPX  |  epv & epw & epx  ;
 FOI <=  EPP & epq & epr  |  epp & EPQ & epr  |  epp & epq & EPR  |  EPP & EPQ & EPR  ;
 fpi <=  EPP & epq & epr  |  epp & EPQ & epr  |  epp & epq & EPR  |  epp & epq & epr  ;
 CCM <= ICM ; 
 CFM <= ICM ; 
 cim <= icm ; 
 CCN <= ICN ; 
 CFN <= ICN ; 
 cin <= icn ; 
 CCO <= ICO ; 
 CFO <= ICO ; 
 cio <= ico ; 
 CCP <= ICP ; 
 CFP <= ICP ; 
 cip <= icp ; 
 DAL <= IDL ; 
 DAM <= IDM ; 
 DAN <= IDN ; 
 DAO <= IDO ; 
 DDO <= IDO ; 
 DDP <= IDP ; 
 DAP <= IDP ; 
 DBA <= IEA ; 
 DEA <= IEA ; 
 dha <= iea ; 
 DBB <= IEB ; 
 DEB <= IEB ; 
 dhb <= ieb ; 
 HAF <=  GAD & ilf & ilj  |  gad & ILF & ilj  |  gad & ilf & ILJ  |  GAD & ILF & ILJ  ;
 hbf <=  GAD & ilf & ilj  |  gad & ILF & ilj  |  gad & ilf & ILJ  |  gad & ilf & ilj  ;
 HAG <= ILI ; 
 HED <=  GDE & geg & gef  |  gde & GEG & gef  |  gde & geg & GEF  |  GDE & GEG & GEF  ;
 hfd <=  GDE & geg & gef  |  gde & GEG & gef  |  gde & geg & GEF  |  gde & geg & gef  ;
 MGA <=  KFB & kgb & lfb  |  kfb & KGB & lfb  |  kfb & kgb & LFB  |  KFB & KGB & LFB  ;
 mha <=  KFB & kgb & lfb  |  kfb & KGB & lfb  |  kfb & kgb & LFB  |  kfb & kgb & lfb  ;
 MGB <= LFA ; 
 HIB <=  GHB & ghc & gic  |  ghb & GHC & gic  |  ghb & ghc & GIC  |  GHB & GHC & GIC  ;
 hjb <=  GHB & ghc & gic  |  ghb & GHC & gic  |  ghb & ghc & GIC  |  ghb & ghc & gic  ;
 HKE <=  GJG & gke & gkg  |  gjg & GKE & gkg  |  gjg & gke & GKG  |  GJG & GKE & GKG  ;
 hle <=  GJG & gke & gkg  |  gjg & GKE & gkg  |  gjg & gke & GKG  |  gjg & gke & gkg  ;
 OHE <=  GVA & gvb & gvc  |  gva & GVB & gvc  |  gva & gvb & GVC  |  GVA & GVB & GVC  ;
 oie <=  GVA & gvb & gvc  |  gva & GVB & gvc  |  gva & gvb & GVC  |  gva & gvb & gvc  ;
 KAD <=  IMF & jab & hae  |  imf & JAB & hae  |  imf & jab & HAE  |  IMF & JAB & HAE  ;
 kbd <=  IMF & jab & hae  |  imf & JAB & hae  |  imf & jab & HAE  |  imf & jab & hae  ;
 KAE <= IMB ; 
 HOC <=  GOD & gne & goe  |  god & GNE & goe  |  god & gne & GOE  |  GOD & GNE & GOE  ;
 hpc <=  GOD & gne & goe  |  god & GNE & goe  |  god & gne & GOE  |  god & gne & goe  ;
 HOE <= GNG ; 
 OPM <=  MMB & mla & mma  |  mmb & MLA & mma  |  mmb & mla & MMA  |  MMB & MLA & MMA  ;
 oqm <=  MMB & mla & mma  |  mmb & MLA & mma  |  mmb & mla & MMA  |  mmb & mla & mma  ;
 KIA <=  JIA & jha & jhb  |  jia & JHA & jhb  |  jia & jha & JHB  |  JIA & JHA & JHB  ;
 kja <=  JIA & jha & jhb  |  jia & JHA & jhb  |  jia & jha & JHB  |  jia & jha & jhb  ;
 KIC <= JIB ; 
 HSB <=  GRB & grc & gsc  |  grb & GRC & gsc  |  grb & grc & GSC  |  GRB & GRC & GSC  ;
 htb <=  GRB & grc & gsc  |  grb & GRC & gsc  |  grb & grc & GSC  |  grb & grc & gsc  ;
 KQA <=  JPA & jqa & jpb  |  jpa & JQA & jpb  |  jpa & jqa & JPB  |  JPA & JQA & JPB  ;
 kra <=  JPA & jqa & jpb  |  jpa & JQA & jpb  |  jpa & jqa & JPB  |  jpa & jqa & jpb  ;
 FQE <=  ERK & erl & erm  |  erk & ERL & erm  |  erk & erl & ERM  |  ERK & ERL & ERM  ;
 fre <=  ERK & erl & erm  |  erk & ERL & erm  |  erk & erl & ERM  |  erk & erl & erm  ;
 FEE <=  EFE & eff & efg  |  efe & EFF & efg  |  efe & eff & EFG  |  EFE & EFF & EFG  ;
 ffe <=  EFE & eff & efg  |  efe & EFF & efg  |  efe & eff & EFG  |  efe & eff & efg  ;
 FSG <=  ETO & etp & etq  |  eto & ETP & etq  |  eto & etp & ETQ  |  ETO & ETP & ETQ  ;
 ftg <=  ETO & etp & etq  |  eto & ETP & etq  |  eto & etp & ETQ  |  eto & etp & etq  ;
 FAK <=  EBI & ebj & ebk  |  ebi & EBJ & ebk  |  ebi & ebj & EBK  |  EBI & EBJ & EBK  ;
 fbk <=  EBI & ebj & ebk  |  ebi & EBJ & ebk  |  ebi & ebj & EBK  |  ebi & ebj & ebk  ;
 FAN <= QIC ; 
 FAL <=  EAU & eav & eaw  |  eau & EAV & eaw  |  eau & eav & EAW  |  EAU & EAV & EAW  ;
 fbl <=  EAU & eav & eaw  |  eau & EAV & eaw  |  eau & eav & EAW  |  eau & eav & eaw  ;
 FQJ <=  ERE & erf & erg  |  ere & ERF & erg  |  ere & erf & ERG  |  ERE & ERF & ERG  ;
 frj <=  ERE & erf & erg  |  ere & ERF & erg  |  ere & erf & ERG  |  ere & erf & erg  ;
 FCJ <=  EDV & edw & edx  |  edv & EDW & edx  |  edv & edw & EDX  |  EDV & EDW & EDX  ;
 fdj <=  EDV & edw & edx  |  edv & EDW & edx  |  edv & edw & EDX  |  edv & edw & edx  ;
 FCK <=  EDJ & edk & edl  |  edj & EDK & edl  |  edj & edk & EDL  |  EDJ & EDK & EDL  ;
 fdk <=  EDJ & edk & edl  |  edj & EDK & edl  |  edj & edk & EDL  |  edj & edk & edl  ;
 FSE <=  ESX & eta & etb  |  esx & ETA & etb  |  esx & eta & ETB  |  ESX & ETA & ETB  ;
 fte <=  ESX & eta & etb  |  esx & ETA & etb  |  esx & eta & ETB  |  esx & eta & etb  ;
 FSF <=  ETC & etd & ete  |  etc & ETD & ete  |  etc & etd & ETE  |  ETC & ETD & ETE  ;
 ftf <=  ETC & etd & ete  |  etc & ETD & ete  |  etc & etd & ETE  |  etc & etd & ete  ;
 FEJ <=  EFW & efx & qic  |  efw & EFX & qic  |  efw & efx & QIC  |  EFW & EFX & QIC  ;
 ffj <=  EFW & efx & qic  |  efw & EFX & qic  |  efw & efx & QIC  |  efw & efx & qic  ;
 FUC <=  EVV & evw & evx  |  evv & EVW & evx  |  evv & evw & EVX  |  EVV & EVW & EVX  ;
 ogc <=  EVV & evw & evx  |  evv & EVW & evx  |  evv & evw & EVX  |  evv & evw & evx  ;
 FEL <=  EEW & eex & efa  |  eew & EEX & efa  |  eew & eex & EFA  |  EEW & EEX & EFA  ;
 ffl <=  EEW & eex & efa  |  eew & EEX & efa  |  eew & eex & EFA  |  eew & eex & efa  ;
 FGE <=  EHF & ehg & ehh  |  ehf & EHG & ehh  |  ehf & ehg & EHH  |  EHF & EHG & EHH  ;
 fhe <=  EHF & ehg & ehh  |  ehf & EHG & ehh  |  ehf & ehg & EHH  |  ehf & ehg & ehh  ;
 FGJ <=  EHL & ehm & ehn  |  ehl & EHM & ehn  |  ehl & ehm & EHN  |  EHL & EHM & EHN  ;
 fhj <=  EHL & ehm & ehn  |  ehl & EHM & ehn  |  ehl & ehm & EHN  |  ehl & ehm & ehn  ;
 FGL <= EHX ; 
 FUH <=  EVS & evt & evu  |  evs & EVT & evu  |  evs & evt & EVU  |  EVS & EVT & EVU  ;
 ogh <=  EVS & evt & evu  |  evs & EVT & evu  |  evs & evt & EVU  |  evs & evt & evu  ;
 FUI <=  EVG & evh & evi  |  evg & EVH & evi  |  evg & evh & EVI  |  EVG & EVH & EVI  ;
 ogi <=  EVG & evh & evi  |  evg & EVH & evi  |  evg & evh & EVI  |  evg & evh & evi  ;
 FUJ <= QIH ; 
 FIE <=  EJG & ejh & eji  |  ejg & EJH & eji  |  ejg & ejh & EJI  |  EJG & EJH & EJI  ;
 fje <=  EJG & ejh & eji  |  ejg & EJH & eji  |  ejg & ejh & EJI  |  ejg & ejh & eji  ;
 FIK <=  EJA & ejb & ejc  |  eja & EJB & ejc  |  eja & ejb & EJC  |  EJA & EJB & EJC  ;
 fjk <=  EJA & ejb & ejc  |  eja & EJB & ejc  |  eja & ejb & EJC  |  eja & ejb & ejc  ;
 FIL <= QID ; 
 FEK <=  EFK & efl & efm  |  efk & EFL & efm  |  efk & efl & EFM  |  EFK & EFL & EFM  ;
 ffk <=  EFK & efl & efm  |  efk & EFL & efm  |  efk & efl & EFM  |  efk & efl & efm  ;
 FKE <=  ELH & eli & elj  |  elh & ELI & elj  |  elh & eli & ELJ  |  ELH & ELI & ELJ  ;
 fle <=  ELH & eli & elj  |  elh & ELI & elj  |  elh & eli & ELJ  |  elh & eli & elj  ;
 FKK <=  ELB & elc & eld  |  elb & ELC & eld  |  elb & elc & ELD  |  ELB & ELC & ELD  ;
 flk <=  ELB & elc & eld  |  elb & ELC & eld  |  elb & elc & ELD  |  elb & elc & eld  ;
 FME <=  ENI & enj & enk  |  eni & ENJ & enk  |  eni & enj & ENK  |  ENI & ENJ & ENK  ;
 fne <=  ENI & enj & enk  |  eni & ENJ & enk  |  eni & enj & ENK  |  eni & enj & enk  ;
 FMJ <=  ENC & endd & ene  |  enc & ENDD  & ene  |  enc & endd & ENE  |  ENC & ENDD  & ENE  ;
 fnj <=  ENC & endd & ene  |  enc & ENDD  & ene  |  enc & endd & ENE  |  enc & endd & ene  ;
 FML <= QIE ; 
 FOE <=  EPJ & epk & epl  |  epj & EPK & epl  |  epj & epk & EPL  |  EPJ & EPK & EPL  ;
 fpe <=  EPJ & epk & epl  |  epj & EPK & epl  |  epj & epk & EPL  |  epj & epk & epl  ;
 FOJ <=  EPD & epe & epf  |  epd & EPE & epf  |  epd & epe & EPF  |  EPD & EPE & EPF  ;
 fpj <=  EPD & epe & epf  |  epd & EPE & epf  |  epd & epe & EPF  |  epd & epe & epf  ;
 FOK <= QIE ; 
 DBC <= IEC ; 
 DEC <= IEC ; 
 dhc <= iec ; 
 DBD <= IED ; 
 DED <= IED ; 
 dhd <= ied ; 
 DCA <= IFA ; 
 DFA <= IFA ; 
 dia <= ifa ; 
 DBE <= IEE ; 
 DEE <= IEE ; 
 dhe <= iee ; 
 DBF <= IEF ; 
 DEF <= IEF ; 
 dhf <= ief ; 
 DBG <= IEG ; 
 DEG <= IEG ; 
 dhg <= ieg ; 
 DBK <= IEK ; 
 DEK <= IEK ; 
 dhk <= iek ; 
 DBH <= IEH ; 
 DEH <= IEH ; 
 dhh <= ieh ; 
 FKJ <=  ELN & elo & elp  |  eln & ELO & elp  |  eln & elo & ELP  |  ELN & ELO & ELP  ;
 flj <=  ELN & elo & elp  |  eln & ELO & elp  |  eln & elo & ELP  |  eln & elo & elp  ;
 DBI <= IEI ; 
 DEI <= IEI ; 
 dhi <= iei ; 
 DBJ <= IEJ ; 
 DEJ <= IEJ ; 
 dhj <= iej ; 
 HCA <=  GBA & gcc & gcb  |  gba & GCC & gcb  |  gba & gcc & GCB  |  GBA & GCC & GCB  ;
 hda <=  GBA & gcc & gcb  |  gba & GCC & gcb  |  gba & gcc & GCB  |  gba & gcc & gcb  ;
 HEE <=  GDH & gdg & geh  |  gdh & GDG & geh  |  gdh & gdg & GEH  |  GDH & GDG & GEH  ;
 hfe <=  GDH & gdg & geh  |  gdh & GDG & geh  |  gdh & gdg & GEH  |  gdh & gdg & geh  ;
 HEF <= GDF ; 
 MIA <=  LIA & lha & lib  |  lia & LHA & lib  |  lia & lha & LIB  |  LIA & LHA & LIB  ;
 mja <=  LIA & lha & lib  |  lia & LHA & lib  |  lia & lha & LIB  |  lia & lha & lib  ;
 HIC <=  GHD & gid & ghe  |  ghd & GID & ghe  |  ghd & gid & GHE  |  GHD & GID & GHE  ;
 hjc <=  GHD & gid & ghe  |  ghd & GID & ghe  |  ghd & gid & GHE  |  ghd & gid & ghe  ;
 MUA <=  LTA & kub & ktb  |  lta & KUB & ktb  |  lta & kub & KTB  |  LTA & KUB & KTB  ;
 oma <=  LTA & kub & ktb  |  lta & KUB & ktb  |  lta & kub & KTB  |  lta & kub & ktb  ;
 MUB <= LUA ; 
 HMA <=  GLA & glb & gma  |  gla & GLB & gma  |  gla & glb & GMA  |  GLA & GLB & GMA  ;
 hna <=  GLA & glb & gma  |  gla & GLB & gma  |  gla & glb & GMA  |  gla & glb & gma  ;
 OHF <=  GVD & gve & gvf  |  gvd & GVE & gvf  |  gvd & gve & GVF  |  GVD & GVE & GVF  ;
 oif <=  GVD & gve & gvf  |  gvd & GVE & gvf  |  gvd & gve & GVF  |  gvd & gve & gvf  ;
 KCA <=  IMK & jba & jca  |  imk & JBA & jca  |  imk & jba & JCA  |  IMK & JBA & JCA  ;
 kda <=  IMK & jba & jca  |  imk & JBA & jca  |  imk & jba & JCA  |  imk & jba & jca  ;
 HOD <=  GNF & gog & gof  |  gnf & GOG & gof  |  gnf & gog & GOF  |  GNF & GOG & GOF  ;
 hpd <=  GNF & gog & gof  |  gnf & GOG & gof  |  gnf & gog & GOF  |  gnf & gog & gof  ;
 HOF <= GNB ; 
 OPO <=  MOA & mob & mna  |  moa & MOB & mna  |  moa & mob & MNA  |  MOA & MOB & MNA  ;
 oqo <=  MOA & mob & mna  |  moa & MOB & mna  |  moa & mob & MNA  |  moa & mob & mna  ;
 KIB <=  JID & jhd & jic  |  jid & JHD & jic  |  jid & jhd & JIC  |  JID & JHD & JIC  ;
 kjb <=  JID & jhd & jic  |  jid & JHD & jic  |  jid & jhd & JIC  |  jid & jhd & jic  ;
 KID <= JHC ; 
 HSC <=  GRD & gre & gsg  |  grd & GRE & gsg  |  grd & gre & GSG  |  GRD & GRE & GSG  ;
 htc <=  GRD & gre & gsg  |  grd & GRE & gsg  |  grd & gre & GSG  |  grd & gre & gsg  ;
 KQB <=  JQC & jpc & jqb  |  jqc & JPC & jqb  |  jqc & jpc & JQB  |  JQC & JPC & JQB  ;
 krb <=  JQC & jpc & jqb  |  jqc & JPC & jqb  |  jqc & jpc & JQB  |  jqc & jpc & jqb  ;
 DBL <= IEL ; 
 DEL <= IEL ; 
 dhl <= iel ; 
 DBM <= IEM ; 
 DEM <= IEM ; 
 dhm <= iem ; 
 DBN <= IEN ; 
 DEN <= IEN ; 
 dhn <= ien ; 
 DBP <= IEP ; 
 DEP <= IEP ; 
 dhp <= iep ; 
 DCB <= IFB ; 
 DFB <= IFB ; 
 dib <= ifb ; 
 HCB <=  GCD & gbb & gca  |  gcd & GBB & gca  |  gcd & gbb & GCA  |  GCD & GBB & GCA  ;
 hdb <=  GCD & gbb & gca  |  gcd & GBB & gca  |  gcd & gbb & GCA  |  gcd & gbb & gca  ;
 HGA <=  GFA & ggb & gga  |  gfa & GGB & gga  |  gfa & ggb & GGA  |  GFA & GGB & GGA  ;
 hha <=  GFA & ggb & gga  |  gfa & GGB & gga  |  gfa & ggb & GGA  |  gfa & ggb & gga  ;
 MKA <=  LKA & lja & lkb  |  lka & LJA & lkb  |  lka & lja & LKB  |  LKA & LJA & LKB  ;
 mla <=  LKA & lja & lkb  |  lka & LJA & lkb  |  lka & lja & LKB  |  lka & lja & lkb  ;
 MKB <= LJB ; 
 HID <=  GHF & ghg & gif  |  ghf & GHG & gif  |  ghf & ghg & GIF  |  GHF & GHG & GIF  ;
 hjd <=  GHF & ghg & gif  |  ghf & GHG & gif  |  ghf & ghg & GIF  |  ghf & ghg & gif  ;
 HIF <= FHF ; 
 HMB <=  GMB & glc & flj  |  gmb & GLC & flj  |  gmb & glc & FLJ  |  GMB & GLC & FLJ  ;
 hnb <=  GMB & glc & flj  |  gmb & GLC & flj  |  gmb & glc & FLJ  |  gmb & glc & flj  ;
 OKC <=  JVA & jvb & jvc  |  jva & JVB & jvc  |  jva & jvb & JVC  |  JVA & JVB & JVC  ;
 olc <=  JVA & jvb & jvc  |  jva & JVB & jvc  |  jva & jvb & JVC  |  jva & jvb & jvc  ;
 KCB <=  HBE & jcb & iml  |  hbe & JCB & iml  |  hbe & jcb & IML  |  HBE & JCB & IML  ;
 kdb <=  HBE & jcb & iml  |  hbe & JCB & iml  |  hbe & jcb & IML  |  hbe & jcb & iml  ;
 HQA <=  GQA & gpa & gpc  |  gqa & GPA & gpc  |  gqa & gpa & GPC  |  GQA & GPA & GPC  ;
 hra <=  GQA & gpa & gpc  |  gqa & GPA & gpc  |  gqa & gpa & GPC  |  gqa & gpa & gpc  ;
 OPQ <=  MQA & mqb & mpa  |  mqa & MQB & mpa  |  mqa & mqb & MPA  |  MQA & MQB & MPA  ;
 oqq <=  MQA & mqb & mpa  |  mqa & MQB & mpa  |  mqa & mqb & MPA  |  mqa & mqb & mpa  ;
 KKA <=  JJB & jkb & jka  |  jjb & JKB & jka  |  jjb & jkb & JKA  |  JJB & JKB & JKA  ;
 kla <=  JJB & jkb & jka  |  jjb & JKB & jka  |  jjb & jkb & JKA  |  jjb & jkb & jka  ;
 KKC <= JJA ; 
 HSD <=  GSE & gsf & grf  |  gse & GSF & grf  |  gse & gsf & GRF  |  GSE & GSF & GRF  ;
 htd <=  GSE & gsf & grf  |  gse & GSF & grf  |  gse & gsf & GRF  |  gse & gsf & grf  ;
 HSE <= GSD ; 
 KSA <=  HSB & jra & jsa  |  hsb & JRA & jsa  |  hsb & jra & JSA  |  HSB & JRA & JSA  ;
 kta <=  HSB & jra & jsa  |  hsb & JRA & jsa  |  hsb & jra & JSA  |  hsb & jra & jsa  ;
 DBO <= IEO ; 
 DEO <= IEO ; 
 dho <= ieo ; 
 FGK <=  EGX & eha & ehb  |  egx & EHA & ehb  |  egx & eha & EHB  |  EGX & EHA & EHB  ;
 fhk <=  EGX & eha & ehb  |  egx & EHA & ehb  |  egx & eha & EHB  |  egx & eha & ehb  ;
 FGM <= QID ; 
 FIJ <=  EJM & ejn & ejo  |  ejm & EJN & ejo  |  ejm & ejn & EJO  |  EJM & EJN & EJO  ;
 fjj <=  EJM & ejn & ejo  |  ejm & EJN & ejo  |  ejm & ejn & EJO  |  ejm & ejn & ejo  ;
 DCK <= IFK ; 
 DFK <= IFK ; 
 dik <= ifk ; 
 DCC <= IFC ; 
 DFC <= IFC ; 
 dic <= ifc ; 
 DCL <= IFL ; 
 DFL <= IFL ; 
 dil <= ifl ; 
 DCD <= IFD ; 
 DFD <= IFD ; 
 did <= ifd ; 
 DCM <= IFM ; 
 DFM <= IFM ; 
 dim <= ifm ; 
 DCE <= IFE ; 
 DFE <= IFE ; 
 die <= ife ; 
 DCN <= IFN ; 
 DFN <= IFN ; 
 din <= ifn ; 
 DCF <= IFFF  ; 
 DFF <= IFFF  ; 
 dif <= ifff  ; 
 DCO <= IFO ; 
 DFO <= IFO ; 
 dio <= ifo ; 
 DCG <= IFG ; 
 DFG <= IFG ; 
 dig <= ifg ; 
 DCP <= IFP ; 
 DFP <= IFP ; 
 dip <= ifp ; 
 DCH <= IFH ; 
 DFH <= IFH ; 
 dih <= ifh ; 
 DCI <= IFI ; 
 DFI <= IFI ; 
 dii <= ifi ; 
 FCL <=  ECV & ecw & ecx  |  ecv & ECW & ecx  |  ecv & ecw & ECX  |  ECV & ECW & ECX  ;
 fdl <=  ECV & ecw & ecx  |  ecv & ECW & ecx  |  ecv & ecw & ECX  |  ecv & ecw & ecx  ;
 FCM <= QIC ; 
 DCJ <= IFJ ; 
 DFJ <= IFJ ; 
 dij <= ifj ; 
end 
endmodule;
