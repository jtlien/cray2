module am( IZZ,
 IAA, 
 IAB, 
 IAC, 
 IAD, 
 IAE, 
 IAF, 
 IAG, 
 IAH, 
 IAI, 
 IAJ, 
 IAK, 
 IAL, 
 IAM, 
 IAN, 
 IAO, 
 IAP, 
 IBA, 
 IBB, 
 IBC, 
 IBD, 
 IBE, 
 IBF, 
 IBG, 
 IBH, 
 IBI, 
 IBJ, 
 IBK, 
 IBL, 
 IBM, 
 IBN, 
 IBO, 
 IBP, 
 ICA, 
 ICB, 
 ICC, 
 ICD, 
 ICE, 
 ICF, 
 ICG, 
 ICH, 
 ICI, 
 ICJ, 
 ICK, 
 ICL, 
 ICM, 
 ICN, 
 ICO, 
 ICP, 
 IDA, 
 IDB, 
 IDC, 
 IDD, 
 IDE, 
 IDF, 
 IDG, 
 IDH, 
 IDI, 
 IDJ, 
 IDK, 
 IDL, 
 IDM, 
 IDN, 
 IDO, 
 IDP, 
 IEA, 
 IEB, 
 IEC, 
 IED, 
 IEE, 
 IEF, 
 IFA, 
 IFB, 
 IFC, 
 IFD, 
 IFE, 
 IFFF, 
 IFG, 
 IGA, 
 IGB, 
 IGC, 
 IGD, 
 IGE, 
 IGF, 
 IHA, 
 OAA, 
 OAB, 
 OAC, 
 OAD, 
 OAE, 
 OAF, 
 OAG, 
 OAH, 
 OAI, 
 OAJ, 
 OAK, 
 OAL, 
 OAM, 
 OAN, 
 OAO, 
 OAP, 
 OBA, 
 OBB, 
 OBC, 
 OBD, 
 OBE, 
 OBF, 
 OBG, 
 OBH, 
 OBI, 
 OBJ, 
 OBK, 
 OBL, 
 OBM, 
 OBN, 
 OBO, 
 OBP, 
 OEA, 
 OEB, 
 OEC, 
 OED, 
 OEE, 
 OEF, 
 OFA, 
 OFB, 
 OFC, 
 OFD, 
 OFE, 
 OFF, 
 OGA, 
 OGB, 
 OGC, 
 OGD, 
 OGE, 
 OGF, 
 OHA, 
 OHB, 
 OHC, 
 OHD, 
 OHE, 
 OHF, 
 OIA, 
 OIB, 
 OIC, 
 OID, 
 OIE, 
 OIF, 
 OIG, 
 OIH, 
 OIJ, 
 OIK, 
 OIL, 
 OIM, 
 OJA, 
 OJB, 
 OJC, 
 OJD, 
 OJE, 
 OJF, 
 OJG, 
 OJH, 
 OJI, 
 OJJ, 
 OJK, 
 OJL, 
 OJM, 
 OKA, 
 OKB, 
 OKC, 
 OKD, 
 OKE, 
 OKF, 
 OKG, 
 OKH, 
 OKI, 
 OKJ, 
 OKK, 
 OKL, 
 OKM, 
 OLA, 
 OLB, 
 OLC, 
 OLD, 
 OLE, 
 OLF, 
 OLG, 
 OLH, 
 OLI, 
 OLJ, 
 OLK, 
 OLL, 
 OLM, 
 OMA, 
 OMB, 
 OMC, 
 OMD, 
 OME, 
 OMF, 
 OMG, 
 OMH, 
 OMI, 
 OMJ, 
 OMK, 
 OML, 
 ONA, 
 ONB, 
 ONC, 
 OND, 
 ONE, 
 ONF, 
 ONG, 
 ONH, 
 ONI, 
 ONJ, 
 ONK, 
 ONL, 
 ONM, 
 OOA, 
 OOB, 
 OOC, 
 OOD, 
 OOE, 
 OOF, 
 OOG, 
 OOH, 
 OOI, 
 OOJ, 
 OOK, 
 OOL, 
 OOM, 
 OPA, 
 OPB, 
 OPC, 
 OPD, 
 OPE, 
 OPF, 
 OPG, 
 OPH, 
 OPI, 
 OPJ, 
 OPK, 
 OPL, 
OPM ); 
    
 input IZZ; 
 input IAA; 
 input IAB; 
 input IAC; 
 input IAD; 
 input IAE; 
 input IAF; 
 input IAG; 
 input IAH; 
 input IAI; 
 input IAJ; 
 input IAK; 
 input IAL; 
 input IAM; 
 input IAN; 
 input IAO; 
 input IAP; 
 input IBA; 
 input IBB; 
 input IBC; 
 input IBD; 
 input IBE; 
 input IBF; 
 input IBG; 
 input IBH; 
 input IBI; 
 input IBJ; 
 input IBK; 
 input IBL; 
 input IBM; 
 input IBN; 
 input IBO; 
 input IBP; 
 input ICA; 
 input ICB; 
 input ICC; 
 input ICD; 
 input ICE; 
 input ICF; 
 input ICG; 
 input ICH; 
 input ICI; 
 input ICJ; 
 input ICK; 
 input ICL; 
 input ICM; 
 input ICN; 
 input ICO; 
 input ICP; 
 input IDA; 
 input IDB; 
 input IDC; 
 input IDD; 
 input IDE; 
 input IDF; 
 input IDG; 
 input IDH; 
 input IDI; 
 input IDJ; 
 input IDK; 
 input IDL; 
 input IDM; 
 input IDN; 
 input IDO; 
 input IDP; 
 input IEA; 
 input IEB; 
 input IEC; 
 input IED; 
 input IEE; 
 input IEF; 
 input IFA; 
 input IFB; 
 input IFC; 
 input IFD; 
 input IFE; 
 input IIFF; 
 input IFG; 
 input IGA; 
 input IGB; 
 input IGC; 
 input IGD; 
 input IGE; 
 input IGF; 
 input IHA; 
 output OAA; 
 output OAB; 
 output OAC; 
 output OAD; 
 output OAE; 
 output OAF; 
 output OAG; 
 output OAH; 
 output OAI; 
 output OAJ; 
 output OAK; 
 output OAL; 
 output OAM; 
 output OAN; 
 output OAO; 
 output OAP; 
 output OBA; 
 output OBB; 
 output OBC; 
 output OBD; 
 output OBE; 
 output OBF; 
 output OBG; 
 output OBH; 
 output OBI; 
 output OBJ; 
 output OBK; 
 output OBL; 
 output OBM; 
 output OBN; 
 output OBO; 
 output OBP; 
 output OEA; 
 output OEB; 
 output OEC; 
 output OED; 
 output OEE; 
 output OEF; 
 output OFA; 
 output OFB; 
 output OFC; 
 output OFD; 
 output OFE; 
 output OFF; 
 output OGA; 
 output OGB; 
 output OGC; 
 output OGD; 
 output OGE; 
 output OGF; 
 output OHA; 
 output OHB; 
 output OHC; 
 output OHD; 
 output OHE; 
 output OHF; 
 output OIA; 
 output OIB; 
 output OIC; 
 output OID; 
 output OIE; 
 output OIF; 
 output OIG; 
 output OIH; 
 output OIJ; 
 output OIK; 
 output OIL; 
 output OIM; 
 output OJA; 
 output OJB; 
 output OJC; 
 output OJD; 
 output OJE; 
 output OJF; 
 output OJG; 
 output OJH; 
 output OJI; 
 output OJJ; 
 output OJK; 
 output OJL; 
 output OJM; 
 output OKA; 
 output OKB; 
 output OKC; 
 output OKD; 
 output OKE; 
 output OKF; 
 output OKG; 
 output OKH; 
 output OKI; 
 output OKJ; 
 output OKK; 
 output OKL; 
 output OKM; 
 output OLA; 
 output OLB; 
 output OLC; 
 output OLD; 
 output OLE; 
 output OLF; 
 output OLG; 
 output OLH; 
 output OLI; 
 output OLJ; 
 output OLK; 
 output OLL; 
 output OLM; 
 output OMA; 
 output OMB; 
 output OMC; 
 output OMD; 
 output OME; 
 output OMF; 
 output OMG; 
 output OMH; 
 output OMI; 
 output OMJ; 
 output OMK; 
 output OML; 
 output ONA; 
 output ONB; 
 output ONC; 
 output OND; 
 output ONE; 
 output ONF; 
 output ONG; 
 output ONH; 
 output ONI; 
 output ONJ; 
 output ONK; 
 output ONL; 
 output ONM; 
 output OOA; 
 output OOB; 
 output OOC; 
 output OOD; 
 output OOE; 
 output OOF; 
 output OOG; 
 output OOH; 
 output OOI; 
 output OOJ; 
 output OOK; 
 output OOL; 
 output OOM; 
 output OPA; 
 output OPB; 
 output OPC; 
 output OPD; 
 output OPE; 
 output OPF; 
 output OPG; 
 output OPH; 
 output OPI; 
 output OPJ; 
 output OPK; 
 output OPL; 
 output OPM; 
  
  
reg  AAA ;
reg  AAB ;
reg  AAC ;
reg  AAD ;
reg  AAE ;
reg  AAF ;
reg  AAG ;
reg  AAH ;
reg  AAI ;
reg  AAJ ;
reg  AAK ;
reg  AAL ;
reg  AAM ;
reg  AAN ;
reg  AAO ;
reg  AAP ;
reg  AAQ ;
reg  ABA ;
reg  ABB ;
reg  ABC ;
reg  ABD ;
reg  ABE ;
reg  ABF ;
reg  ABG ;
reg  ABH ;
reg  ABI ;
reg  ABJ ;
reg  ABK ;
reg  ABL ;
reg  ABM ;
reg  ABN ;
reg  ABO ;
reg  ABP ;
reg  ACA ;
reg  ACB ;
reg  ACC ;
reg  ACD ;
reg  ACE ;
reg  ACF ;
reg  ACG ;
reg  ACH ;
reg  ACI ;
reg  ACJ ;
reg  ACK ;
reg  ACL ;
reg  ACM ;
reg  ACN ;
reg  ACO ;
reg  ACP ;
reg  ACQ ;
reg  ADA ;
reg  ADB ;
reg  ADC ;
reg  ADD ;
reg  ADE ;
reg  ADF ;
reg  ADG ;
reg  ADH ;
reg  ADI ;
reg  ADJ ;
reg  ADK ;
reg  ADL ;
reg  ADM ;
reg  ADN ;
reg  ADO ;
reg  ADP ;
reg  BAA ;
reg  BAB ;
reg  BAC ;
reg  BAD ;
reg  BAE ;
reg  BAF ;
reg  BAG ;
reg  BAH ;
reg  BAI ;
reg  BAJ ;
reg  BAK ;
reg  BAL ;
reg  BAM ;
reg  BAN ;
reg  BAO ;
reg  BAP ;
reg  BBA ;
reg  BBB ;
reg  BBC ;
reg  BBD ;
reg  BBE ;
reg  BBF ;
reg  BBG ;
reg  BBH ;
reg  BBI ;
reg  BBJ ;
reg  BBK ;
reg  BBL ;
reg  BBM ;
reg  BBN ;
reg  BBO ;
reg  BBP ;
reg  DGA ;
reg  DGB ;
reg  DHA ;
reg  DHB ;
reg  DHC ;
reg  DHD ;
reg  DHE ;
reg  dhf ;
reg  DIA ;
reg  dib ;
reg  DIC ;
reg  did ;
reg  DIE ;
reg  DJA ;
reg  djb ;
reg  DJC ;
reg  DKA ;
reg  dkb ;
reg  DKC ;
reg  DKD ;
reg  DLA ;
reg  dlb ;
reg  DLC ;
reg  DLD ;
reg  DMA ;
reg  dmb ;
reg  DMC ;
reg  dmd ;
reg  DNA ;
reg  dnb ;
reg  DNC ;
reg  dnd ;
reg  DOA ;
reg  dob ;
reg  DOC ;
reg  dod ;
reg  DOE ;
reg  DPA ;
reg  dpb ;
reg  DPC ;
reg  dpd ;
reg  DPE ;
reg  DQA ;
reg  dqb ;
reg  DQC ;
reg  dqd ;
reg  DQE ;
reg  DQF ;
reg  DRA ;
reg  drb ;
reg  DRC ;
reg  drd ;
reg  DRE ;
reg  DRF ;
reg  DSA ;
reg  dsb ;
reg  DSC ;
reg  dsd ;
reg  DSE ;
reg  dsf ;
reg  DTA ;
reg  dtb ;
reg  DTC ;
reg  dtd ;
reg  DTE ;
reg  dtf ;
reg  DUA ;
reg  dub ;
reg  DUC ;
reg  dud ;
reg  DUE ;
reg  duf ;
reg  DUG ;
reg  DVA ;
reg  dvb ;
reg  DVC ;
reg  dvd ;
reg  DVE ;
reg  dvf ;
reg  DVG ;
reg  DWA ;
reg  dwb ;
reg  DWC ;
reg  dwd ;
reg  DWE ;
reg  dwf ;
reg  DWG ;
reg  DWH ;
reg  DXA ;
reg  dxb ;
reg  DXC ;
reg  dxd ;
reg  DXE ;
reg  dxf ;
reg  DXG ;
reg  DXH ;
reg  DYA ;
reg  dyb ;
reg  DYC ;
reg  dyd ;
reg  DYE ;
reg  dyf ;
reg  DYG ;
reg  dyh ;
reg  DZA ;
reg  dzb ;
reg  DZC ;
reg  dzd ;
reg  DZE ;
reg  dzf ;
reg  DZG ;
reg  dzh ;
reg  DZI ;
reg  dzj ;
reg  DZK ;
reg  dzl ;
reg  DZM ;
reg  dzn ;
reg  DZO ;
reg  dzp ;
reg  DZQ ;
reg  FAA ;
reg  FBA ;
reg  FCA ;
reg  FCB ;
reg  FDA ;
reg  FDB ;
reg  FEA ;
reg  FFA ;
reg  FFB ;
reg  FGA ;
reg  FHA ;
reg  FHB ;
reg  FIA ;
reg  fib ;
reg  FJA ;
reg  fjb ;
reg  FMA ;
reg  FMB ;
reg  FNA ;
reg  fnb ;
reg  FOA ;
reg  fob ;
reg  FOC ;
reg  FPA ;
reg  fpb ;
reg  FPC ;
reg  FQA ;
reg  fqb ;
reg  FQC ;
reg  FRA ;
reg  frb ;
reg  FRC ;
reg  FRD ;
reg  FSA ;
reg  fsb ;
reg  FSC ;
reg  FSD ;
reg  FTA ;
reg  ftb ;
reg  FTC ;
reg  FUA ;
reg  fub ;
reg  FUC ;
reg  FUD ;
reg  FVA ;
reg  fvb ;
reg  FVC ;
reg  fvd ;
reg  FWA ;
reg  fwb ;
reg  FWC ;
reg  FWD ;
reg  FXA ;
reg  fxb ;
reg  FXC ;
reg  fxd ;
reg  FXE ;
reg  FYA ;
reg  fyb ;
reg  FYC ;
reg  FYD ;
reg  FYE ;
reg  fyf ;
reg  FYG ;
reg  fyh ;
reg  FYI ;
reg  FYJ ;
reg  fyk ;
reg  FYL ;
reg  fym ;
reg  FYN ;
reg  FYO ;
reg  fyp ;
reg  FYQ ;
reg  fyr ;
reg  FYS ;
reg  FZA ;
reg  fzb ;
reg  FZC ;
reg  fzd ;
reg  FZE ;
reg  fzf ;
reg  FZG ;
reg  FZH ;
reg  FZI ;
reg  fzj ;
reg  FZK ;
reg  fzl ;
reg  FZM ;
reg  fzn ;
reg  FZO ;
reg  fzp ;
reg  FZR ;
reg  fzs ;
reg  FZT ;
reg  fzu ;
reg  FZV ;
reg  FZW ;
reg  fzx ;
reg  FZY ;
reg  fzz ;
reg  GZK ;
reg  HAA ;
reg  HBA ;
reg  HCA ;
reg  HCB ;
reg  HDA ;
reg  HDB ;
reg  HEA ;
reg  HFA ;
reg  HFB ;
reg  HGA ;
reg  HGB ;
reg  HHA ;
reg  HHB ;
reg  HIA ;
reg  HJA ;
reg  HJB ;
reg  HMA ;
reg  HNA ;
reg  HNB ;
reg  HOA ;
reg  HPA ;
reg  HPB ;
reg  HQA ;
reg  HQB ;
reg  HRA ;
reg  hrb ;
reg  HSA ;
reg  hsb ;
reg  HTA ;
reg  HTB ;
reg  HUA ;
reg  hub ;
reg  HVA ;
reg  hvb ;
reg  HWA ;
reg  hwb ;
reg  HXA ;
reg  hxb ;
reg  HXC ;
reg  HYA ;
reg  hyb ;
reg  HYD ;
reg  HZA ;
reg  hzb ;
reg  HZC ;
reg  hzd ;
reg  HZG ;
reg  hzh ;
reg  HZI ;
reg  hzj ;
reg  HZK ;
reg  HZM ;
reg  hzn ;
reg  HZO ;
reg  HZQ ;
reg  hzr ;
reg  HZT ;
reg  hzu ;
reg  HZV ;
reg  HZW ;
reg  hzx ;
reg  HZY ;
reg  hzz ;
reg  KAA ;
reg  KBA ;
reg  KCA ;
reg  KCB ;
reg  KDA ;
reg  KDB ;
reg  KEA ;
reg  KFA ;
reg  KGA ;
reg  KHA ;
reg  khb ;
reg  KIA ;
reg  KJA ;
reg  KJB ;
reg  KMA ;
reg  KNA ;
reg  KNB ;
reg  KOA ;
reg  KPA ;
reg  KPB ;
reg  KQA ;
reg  KQB ;
reg  KRA ;
reg  KSA ;
reg  KSB ;
reg  KTA ;
reg  KTB ;
reg  KUA ;
reg  KUB ;
reg  KVA ;
reg  KVB ;
reg  KWA ;
reg  KWB ;
reg  KXA ;
reg  kxb ;
reg  KYA ;
reg  KYB ;
reg  KZA ;
reg  KZB ;
reg  KZC ;
reg  KZD ;
reg  KZG ;
reg  KZH ;
reg  KZI ;
reg  kzj ;
reg  KZM ;
reg  kzn ;
reg  KZQ ;
reg  KZR ;
reg  KZT ;
reg  KZW ;
reg  KZX ;
reg  KZY ;
reg  MAA ;
reg  MBA ;
reg  MBB ;
reg  MCA ;
reg  MDA ;
reg  mdb ;
reg  MEA ;
reg  MEB ;
reg  MFA ;
reg  MFB ;
reg  MGA ;
reg  MGB ;
reg  MHA ;
reg  MHB ;
reg  MIA ;
reg  mib ;
reg  MJA ;
reg  mjb ;
reg  MKA ;
reg  MKB ;
reg  MLA ;
reg  MLB ;
reg  MMA ;
reg  MMB ;
reg  MNA ;
reg  MNB ;
reg  MOA ;
reg  mob ;
reg  MQA ;
reg  MQB ;
reg  MRA ;
reg  MRB ;
reg  MSA ;
reg  msb ;
reg  MTA ;
reg  mtb ;
reg  MUA ;
reg  mub ;
reg  MVA ;
reg  mvb ;
reg  MWA ;
reg  mwb ;
reg  MXA ;
reg  mxb ;
reg  MYA ;
reg  myb ;
reg  MZA ;
reg  mzb ;
reg  MZD ;
reg  mze ;
reg  MZI ;
reg  mzj ;
reg  MZL ;
reg  mzm ;
reg  MZO ;
reg  mzp ;
reg  MZR ;
reg  mzs ;
reg  MZU ;
reg  mzv ;
reg  MZX ;
reg  mzy ;
reg  NAA ;
reg  NAB ;
reg  NAC ;
reg  NAD ;
reg  NAE ;
reg  NAF ;
reg  NAG ;
reg  NAH ;
reg  NAI ;
reg  NAJ ;
reg  NAK ;
reg  NAL ;
reg  NAM ;
reg  NAN ;
reg  NAO ;
reg  NAP ;
reg  NAQ ;
reg  NBA ;
reg  NBB ;
reg  NBC ;
reg  NBD ;
reg  NBE ;
reg  NBF ;
reg  NBG ;
reg  NBH ;
reg  NBI ;
reg  NBJ ;
reg  NBK ;
reg  NBL ;
reg  NBM ;
reg  NBN ;
reg  NBO ;
reg  NBP ;
reg  NEB ;
reg  NEE ;
reg  NEF ;
reg  NEG ;
reg  NEH ;
reg  NEI ;
reg  NEJ ;
reg  NEK ;
reg  NEL ;
reg  NEM ;
reg  NEN ;
reg  NEO ;
reg  NEP ;
reg  NFB ;
reg  NFC ;
reg  NFD ;
reg  NFE ;
reg  NFF ;
reg  NFG ;
reg  NFH ;
reg  NFI ;
reg  NFJ ;
reg  NFK ;
reg  NFL ;
reg  NFM ;
reg  NFN ;
reg  NFO ;
reg  NFP ;
reg  OAA ;
reg  OAB ;
reg  OAC ;
reg  OAD ;
reg  OAE ;
reg  OAF ;
reg  OAG ;
reg  OAH ;
reg  OAI ;
reg  OAJ ;
reg  OAK ;
reg  OAL ;
reg  OAM ;
reg  OAN ;
reg  OAO ;
reg  OAP ;
reg  OBA ;
reg  OBB ;
reg  OBC ;
reg  OBD ;
reg  OBE ;
reg  OBF ;
reg  OBG ;
reg  OBH ;
reg  OBI ;
reg  OBJ ;
reg  OBK ;
reg  OBL ;
reg  OBM ;
reg  OBN ;
reg  OBO ;
reg  OBP ;
reg  OEA ;
reg  OEB ;
reg  OEC ;
reg  OED ;
reg  OEE ;
reg  OEF ;
reg  OFA ;
reg  OFB ;
reg  OFC ;
reg  OFD ;
reg  OFE ;
reg  OFF ;
reg  oga ;
reg  ogb ;
reg  ogc ;
reg  ogd ;
reg  oge ;
reg  ogf ;
reg  oha ;
reg  ohb ;
reg  ohc ;
reg  ohd ;
reg  ohe ;
reg  ohf ;
reg  oia ;
reg  oib ;
reg  oic ;
reg  oid ;
reg  oie ;
reg  oif ;
reg  oig ;
reg  oih ;
reg  oii ;
reg  oij ;
reg  oik ;
reg  oil ;
reg  oim ;
reg  OJA ;
reg  OJB ;
reg  OJC ;
reg  OJD ;
reg  OJE ;
reg  OJF ;
reg  OJG ;
reg  OJH ;
reg  OJI ;
reg  OJJ ;
reg  OJK ;
reg  OJL ;
reg  OJM ;
reg  oka ;
reg  okb ;
reg  okc ;
reg  okd ;
reg  oke ;
reg  okf ;
reg  okg ;
reg  okh ;
reg  oki ;
reg  okj ;
reg  okk ;
reg  okl ;
reg  okm ;
reg  OLA ;
reg  OLB ;
reg  OLC ;
reg  OLD ;
reg  OLE ;
reg  OLF ;
reg  OLG ;
reg  OLH ;
reg  OLI ;
reg  OLJ ;
reg  OLK ;
reg  OLL ;
reg  OLM ;
reg  oma ;
reg  omb ;
reg  omc ;
reg  omd ;
reg  ome ;
reg  omf ;
reg  omg ;
reg  omh ;
reg  omi ;
reg  omj ;
reg  omk ;
reg  oml ;
reg  omm ;
reg  ONA ;
reg  ONB ;
reg  ONC ;
reg  OND ;
reg  ONE ;
reg  ONF ;
reg  ONG ;
reg  ONH ;
reg  ONI ;
reg  ONJ ;
reg  ONK ;
reg  ONL ;
reg  ONM ;
reg  ooa ;
reg  oob ;
reg  ooc ;
reg  ood ;
reg  ooe ;
reg  oof ;
reg  oog ;
reg  ooh ;
reg  ooi ;
reg  ooj ;
reg  ook ;
reg  ool ;
reg  oom ;
reg  OPA ;
reg  OPB ;
reg  OPC ;
reg  OPD ;
reg  OPE ;
reg  OPF ;
reg  OPG ;
reg  OPH ;
reg  OPI ;
reg  OPJ ;
reg  OPK ;
reg  OPL ;
reg  OPM ;
reg  PAB ;
reg  PAC ;
reg  PAD ;
reg  PAE ;
reg  PAF ;
reg  PAG ;
reg  PAH ;
reg  pai ;
reg  pak ;
reg  PAL ;
reg  PAO ;
reg  PAQ ;
reg  PBA ;
reg  PBB ;
reg  PBC ;
reg  PBD ;
reg  PBE ;
reg  PBF ;
reg  PBG ;
reg  PBH ;
reg  PBI ;
reg  PBJ ;
reg  PBK ;
reg  PBL ;
reg  PBM ;
reg  PBN ;
reg  PBO ;
reg  PBP ;
reg  PCA ;
reg  PCB ;
reg  PCC ;
reg  PCD ;
reg  PCE ;
reg  PCF ;
reg  PCG ;
reg  PCH ;
reg  PCI ;
reg  PCJ ;
reg  PCK ;
reg  PCL ;
reg  PCM ;
reg  PCN ;
reg  PCO ;
reg  PCP ;
reg  PDE ;
reg  PDF ;
reg  PDG ;
reg  PDH ;
reg  PDI ;
reg  PDJ ;
reg  PDK ;
reg  PDL ;
reg  PDM ;
reg  PDN ;
reg  PDO ;
reg  PDP ;
reg  PEA ;
reg  PEB ;
reg  PEC ;
reg  PED ;
reg  PEE ;
reg  PEF ;
reg  PEG ;
reg  PEH ;
reg  PEI ;
reg  PEJ ;
reg  PEK ;
reg  PEL ;
reg  PEM ;
reg  PEN ;
reg  PEO ;
reg  PEP ;
reg  PFA ;
reg  PFB ;
reg  PFC ;
reg  PFD ;
reg  PFE ;
reg  PFF ;
reg  PFG ;
reg  PFH ;
reg  PFI ;
reg  PFJ ;
reg  PFK ;
reg  PFL ;
reg  PFM ;
reg  PFN ;
reg  PFO ;
reg  PFP ;
reg  PGA ;
reg  PGB ;
reg  PGC ;
reg  PGD ;
reg  PGE ;
reg  PGF ;
reg  PGG ;
reg  PGH ;
reg  PGI ;
reg  PGJ ;
reg  PGK ;
reg  PGL ;
reg  PGM ;
reg  PGN ;
reg  PGO ;
reg  PGP ;
reg  QAA ;
reg  QAB ;
reg  QAC ;
reg  QAD ;
reg  QAE ;
reg  QAF ;
reg  QAG ;
reg  QAH ;
reg  QAI ;
reg  QAJ ;
reg  QAK ;
reg  QAL ;
reg  qva ;
reg  QVB ;
reg  qvc ;
reg  QVD ;
reg  qve ;
reg  QVF ;
reg  QVG ;
reg  QXA ;
reg  qxb ;
reg  QXC ;
reg  qxd ;
reg  QXE ;
reg  qxf ;
reg  QXG ;
reg  qxh ;
reg  QXI ;
reg  qxj ;
reg  QXK ;
reg  qxl ;
reg  QXM ;
reg  qxn ;
reg  QXO ;
reg  qxp ;
reg  QXQ ;
reg  qxr ;
reg  QXS ;
reg  qxt ;
reg  QXU ;
reg  QXV ;
reg  qxw ;
reg  QXX ;
reg  qxy ;
reg  QXZ ;
reg  QYA ;
reg  qyb ;
reg  QYC ;
reg  qyd ;
reg  QYE ;
reg  qyf ;
reg  QYG ;
reg  qyh ;
reg  QYI ;
reg  QYJ ;
reg  qyk ;
reg  QYL ;
reg  qym ;
reg  QYN ;
reg  qyo ;
reg  QYP ;
reg  qyq ;
reg  QYR ;
reg  QYS ;
reg  QZA ;
reg  qzb ;
reg  QZC ;
reg  qzd ;
reg  QZE ;
reg  qzf ;
reg  QZG ;
reg  qzh ;
reg  QZI ;
reg  QZJ ;
reg  QZK ;
reg  qzl ;
reg  QZM ;
reg  qzn ;
reg  QZO ;
reg  qzp ;
reg  QZQ ;
reg  qzr ;
reg  QZS ;
reg  qzt ;
reg  TFA ;
reg  TFB ;
reg  TFC ;
reg  TFD ;
wire  aaa ;
wire  aab ;
wire  aac ;
wire  aad ;
wire  aae ;
wire  aaf ;
wire  aag ;
wire  aah ;
wire  aai ;
wire  aaj ;
wire  aak ;
wire  aal ;
wire  aam ;
wire  aan ;
wire  aao ;
wire  aap ;
wire  aaq ;
wire  aba ;
wire  abb ;
wire  abc ;
wire  abd ;
wire  abe ;
wire  abf ;
wire  abg ;
wire  abh ;
wire  abi ;
wire  abj ;
wire  abk ;
wire  abl ;
wire  abm ;
wire  abn ;
wire  abo ;
wire  abp ;
wire  aca ;
wire  acb ;
wire  acc ;
wire  acd ;
wire  ace ;
wire  acf ;
wire  acg ;
wire  ach ;
wire  aci ;
wire  acj ;
wire  ack ;
wire  acl ;
wire  acm ;
wire  acn ;
wire  aco ;
wire  acp ;
wire  acq ;
wire  ada ;
wire  adb ;
wire  adc ;
wire  add ;
wire  ade ;
wire  adf ;
wire  adg ;
wire  adh ;
wire  adi ;
wire  adj ;
wire  adk ;
wire  adl ;
wire  adm ;
wire  adn ;
wire  ado ;
wire  adp ;
wire  baa ;
wire  bab ;
wire  bac ;
wire  bad ;
wire  bae ;
wire  baf ;
wire  bag ;
wire  bah ;
wire  bai ;
wire  baj ;
wire  bak ;
wire  bal ;
wire  bam ;
wire  ban ;
wire  bao ;
wire  bap ;
wire  bba ;
wire  bbb ;
wire  bbc ;
wire  bbd ;
wire  bbe ;
wire  bbf ;
wire  bbg ;
wire  bbh ;
wire  bbi ;
wire  bbj ;
wire  bbk ;
wire  bbl ;
wire  bbm ;
wire  bbn ;
wire  bbo ;
wire  bbp ;
wire  caa ;
wire  CAA ;
wire  cab ;
wire  CAB ;
wire  cac ;
wire  CAC ;
wire  cad ;
wire  CAD ;
wire  cae ;
wire  CAE ;
wire  caf ;
wire  CAF ;
wire  cag ;
wire  CAG ;
wire  cah ;
wire  CAH ;
wire  cai ;
wire  CAI ;
wire  caj ;
wire  CAJ ;
wire  cak ;
wire  CAK ;
wire  cal ;
wire  CAL ;
wire  cam ;
wire  CAM ;
wire  can ;
wire  CAN ;
wire  cao ;
wire  CAO ;
wire  cap ;
wire  CAP ;
wire  cba ;
wire  CBA ;
wire  cbb ;
wire  CBB ;
wire  cbc ;
wire  CBC ;
wire  cbd ;
wire  CBD ;
wire  cbe ;
wire  CBE ;
wire  cbf ;
wire  CBF ;
wire  cbg ;
wire  CBG ;
wire  cbh ;
wire  CBH ;
wire  cbi ;
wire  CBI ;
wire  cbj ;
wire  CBJ ;
wire  cbk ;
wire  CBK ;
wire  cbl ;
wire  CBL ;
wire  cbm ;
wire  CBM ;
wire  cbn ;
wire  CBN ;
wire  cbo ;
wire  CBO ;
wire  cbp ;
wire  CBP ;
wire  cca ;
wire  CCA ;
wire  ccb ;
wire  CCB ;
wire  ccc ;
wire  CCC ;
wire  ccd ;
wire  CCD ;
wire  cce ;
wire  CCE ;
wire  ccf ;
wire  CCF ;
wire  ccg ;
wire  CCG ;
wire  cch ;
wire  CCH ;
wire  cci ;
wire  CCI ;
wire  ccj ;
wire  CCJ ;
wire  cck ;
wire  CCK ;
wire  ccl ;
wire  CCL ;
wire  ccm ;
wire  CCM ;
wire  ccn ;
wire  CCN ;
wire  cco ;
wire  CCO ;
wire  cda ;
wire  CDA ;
wire  cdb ;
wire  CDB ;
wire  cdc ;
wire  CDC ;
wire  cdd ;
wire  CDD ;
wire  cde ;
wire  CDE ;
wire  cdf ;
wire  CDF ;
wire  cdg ;
wire  CDG ;
wire  cdh ;
wire  CDH ;
wire  cdi ;
wire  CDI ;
wire  cdj ;
wire  CDJ ;
wire  cdk ;
wire  CDK ;
wire  cdl ;
wire  CDL ;
wire  cdm ;
wire  CDM ;
wire  cdn ;
wire  CDN ;
wire  cdo ;
wire  CDO ;
wire  cea ;
wire  CEA ;
wire  ceb ;
wire  CEB ;
wire  cec ;
wire  CEC ;
wire  ced ;
wire  CED ;
wire  cee ;
wire  CEE ;
wire  cef ;
wire  CEF ;
wire  ceg ;
wire  CEG ;
wire  ceh ;
wire  CEH ;
wire  cei ;
wire  CEI ;
wire  cej ;
wire  CEJ ;
wire  cek ;
wire  CEK ;
wire  cel ;
wire  CEL ;
wire  cem ;
wire  CEM ;
wire  cen ;
wire  CEN ;
wire  cfa ;
wire  CFA ;
wire  cfb ;
wire  CFB ;
wire  cfc ;
wire  CFC ;
wire  cfd ;
wire  CFD ;
wire  cfe ;
wire  CFE ;
wire  cff ;
wire  CFF ;
wire  cfg ;
wire  CFG ;
wire  cfh ;
wire  CFH ;
wire  cfi ;
wire  CFI ;
wire  cfj ;
wire  CFJ ;
wire  cfk ;
wire  CFK ;
wire  cfl ;
wire  CFL ;
wire  cfm ;
wire  CFM ;
wire  cfn ;
wire  CFN ;
wire  cga ;
wire  CGA ;
wire  cgb ;
wire  CGB ;
wire  cgc ;
wire  CGC ;
wire  cgd ;
wire  CGD ;
wire  cge ;
wire  CGE ;
wire  cgf ;
wire  CGF ;
wire  cgg ;
wire  CGG ;
wire  cgh ;
wire  CGH ;
wire  cgi ;
wire  CGI ;
wire  cgj ;
wire  CGJ ;
wire  cgk ;
wire  CGK ;
wire  cgl ;
wire  CGL ;
wire  cgm ;
wire  CGM ;
wire  cha ;
wire  CHA ;
wire  chb ;
wire  CHB ;
wire  chc ;
wire  CHC ;
wire  chd ;
wire  CHD ;
wire  che ;
wire  CHE ;
wire  chf ;
wire  CHF ;
wire  chg ;
wire  CHG ;
wire  chh ;
wire  CHH ;
wire  chi ;
wire  CHI ;
wire  chj ;
wire  CHJ ;
wire  chk ;
wire  CHK ;
wire  chl ;
wire  CHL ;
wire  chm ;
wire  CHM ;
wire  cia ;
wire  CIA ;
wire  cib ;
wire  CIB ;
wire  cic ;
wire  CIC ;
wire  cid ;
wire  CID ;
wire  cie ;
wire  CIE ;
wire  cif ;
wire  CIF ;
wire  cig ;
wire  CIG ;
wire  cih ;
wire  CIH ;
wire  cii ;
wire  CII ;
wire  cij ;
wire  CIJ ;
wire  cik ;
wire  CIK ;
wire  cil ;
wire  CIL ;
wire  cja ;
wire  CJA ;
wire  cjb ;
wire  CJB ;
wire  cjc ;
wire  CJC ;
wire  cjd ;
wire  CJD ;
wire  cje ;
wire  CJE ;
wire  cjf ;
wire  CJF ;
wire  cjg ;
wire  CJG ;
wire  cjh ;
wire  CJH ;
wire  cji ;
wire  CJI ;
wire  cjj ;
wire  CJJ ;
wire  cjk ;
wire  CJK ;
wire  cjl ;
wire  CJL ;
wire  cka ;
wire  CKA ;
wire  ckb ;
wire  CKB ;
wire  ckc ;
wire  CKC ;
wire  ckd ;
wire  CKD ;
wire  cke ;
wire  CKE ;
wire  ckf ;
wire  CKF ;
wire  ckg ;
wire  CKG ;
wire  ckh ;
wire  CKH ;
wire  cki ;
wire  CKI ;
wire  ckj ;
wire  CKJ ;
wire  ckk ;
wire  CKK ;
wire  cla ;
wire  CLA ;
wire  clb ;
wire  CLB ;
wire  clc ;
wire  CLC ;
wire  cld ;
wire  CLD ;
wire  cle ;
wire  CLE ;
wire  clf ;
wire  CLF ;
wire  clg ;
wire  CLG ;
wire  clh ;
wire  CLH ;
wire  cli ;
wire  CLI ;
wire  clj ;
wire  CLJ ;
wire  clk ;
wire  CLK ;
wire  cma ;
wire  CMA ;
wire  cmb ;
wire  CMB ;
wire  cmc ;
wire  CMC ;
wire  cmd ;
wire  CMD ;
wire  cme ;
wire  CME ;
wire  cmf ;
wire  CMF ;
wire  cmg ;
wire  CMG ;
wire  cmh ;
wire  CMH ;
wire  cmi ;
wire  CMI ;
wire  cmj ;
wire  CMJ ;
wire  cna ;
wire  CNA ;
wire  cnb ;
wire  CNB ;
wire  cnc ;
wire  CNC ;
wire  cnd ;
wire  CND ;
wire  cne ;
wire  CNE ;
wire  cnf ;
wire  CNF ;
wire  cng ;
wire  CNG ;
wire  cnh ;
wire  CNH ;
wire  cni ;
wire  CNI ;
wire  cnj ;
wire  CNJ ;
wire  coa ;
wire  COA ;
wire  cob ;
wire  COB ;
wire  coc ;
wire  COC ;
wire  cod ;
wire  COD ;
wire  coe ;
wire  COE ;
wire  cof ;
wire  COF ;
wire  cog ;
wire  COG ;
wire  coh ;
wire  COH ;
wire  coi ;
wire  COI ;
wire  cpa ;
wire  CPA ;
wire  cpb ;
wire  CPB ;
wire  cpc ;
wire  CPC ;
wire  cpd ;
wire  CPD ;
wire  cpe ;
wire  CPE ;
wire  cpf ;
wire  CPF ;
wire  cpg ;
wire  CPG ;
wire  cph ;
wire  CPH ;
wire  cpi ;
wire  CPI ;
wire  cqa ;
wire  CQA ;
wire  cqb ;
wire  CQB ;
wire  cqc ;
wire  CQC ;
wire  cqd ;
wire  CQD ;
wire  cqe ;
wire  CQE ;
wire  cqf ;
wire  CQF ;
wire  cqg ;
wire  CQG ;
wire  cqh ;
wire  CQH ;
wire  cra ;
wire  CRA ;
wire  crb ;
wire  CRB ;
wire  crc ;
wire  CRC ;
wire  crd ;
wire  CRD ;
wire  cre ;
wire  CRE ;
wire  crf ;
wire  CRF ;
wire  crg ;
wire  CRG ;
wire  crh ;
wire  CRH ;
wire  csa ;
wire  CSA ;
wire  csb ;
wire  CSB ;
wire  csc ;
wire  CSC ;
wire  csd ;
wire  CSD ;
wire  cse ;
wire  CSE ;
wire  csf ;
wire  CSF ;
wire  csg ;
wire  CSG ;
wire  cta ;
wire  CTA ;
wire  ctb ;
wire  CTB ;
wire  ctc ;
wire  CTC ;
wire  ctd ;
wire  CTD ;
wire  cte ;
wire  CTE ;
wire  ctf ;
wire  CTF ;
wire  ctg ;
wire  CTG ;
wire  cua ;
wire  CUA ;
wire  cub ;
wire  CUB ;
wire  cuc ;
wire  CUC ;
wire  cud ;
wire  CUD ;
wire  cue ;
wire  CUE ;
wire  cuf ;
wire  CUF ;
wire  cva ;
wire  CVA ;
wire  cvb ;
wire  CVB ;
wire  cvc ;
wire  CVC ;
wire  cvd ;
wire  CVD ;
wire  cve ;
wire  CVE ;
wire  cvf ;
wire  CVF ;
wire  cwa ;
wire  CWA ;
wire  cwb ;
wire  CWB ;
wire  cwc ;
wire  CWC ;
wire  cwd ;
wire  CWD ;
wire  cwe ;
wire  CWE ;
wire  cxa ;
wire  CXA ;
wire  cxb ;
wire  CXB ;
wire  cxc ;
wire  CXC ;
wire  cxd ;
wire  CXD ;
wire  cxe ;
wire  CXE ;
wire  cya ;
wire  CYA ;
wire  cyb ;
wire  CYB ;
wire  cyc ;
wire  CYC ;
wire  cyd ;
wire  CYD ;
wire  cza ;
wire  CZA ;
wire  czb ;
wire  CZB ;
wire  czc ;
wire  CZC ;
wire  czd ;
wire  CZD ;
wire  daa ;
wire  DAA ;
wire  dab ;
wire  DAB ;
wire  dac ;
wire  DAC ;
wire  dba ;
wire  DBA ;
wire  dbb ;
wire  DBB ;
wire  dbc ;
wire  DBC ;
wire  dca ;
wire  DCA ;
wire  dcb ;
wire  DCB ;
wire  dda ;
wire  DDA ;
wire  ddb ;
wire  DDB ;
wire  dea ;
wire  DEA ;
wire  dfa ;
wire  DFA ;
wire  dga ;
wire  dgb ;
wire  dha ;
wire  dhb ;
wire  dhc ;
wire  dhd ;
wire  dhe ;
wire  DHF ;
wire  dia ;
wire  DIB ;
wire  dic ;
wire  DID ;
wire  die ;
wire  dja ;
wire  DJB ;
wire  djc ;
wire  dka ;
wire  DKB ;
wire  dkc ;
wire  dkd ;
wire  dla ;
wire  DLB ;
wire  dlc ;
wire  dld ;
wire  dma ;
wire  DMB ;
wire  dmc ;
wire  DMD ;
wire  dna ;
wire  DNB ;
wire  dnc ;
wire  DND ;
wire  doa ;
wire  DOB ;
wire  doc ;
wire  DOD ;
wire  doe ;
wire  dpa ;
wire  DPB ;
wire  dpc ;
wire  DPD ;
wire  dpe ;
wire  dqa ;
wire  DQB ;
wire  dqc ;
wire  DQD ;
wire  dqe ;
wire  dqf ;
wire  dra ;
wire  DRB ;
wire  drc ;
wire  DRD ;
wire  dre ;
wire  drf ;
wire  dsa ;
wire  DSB ;
wire  dsc ;
wire  DSD ;
wire  dse ;
wire  DSF ;
wire  dta ;
wire  DTB ;
wire  dtc ;
wire  DTD ;
wire  dte ;
wire  DTF ;
wire  dua ;
wire  DUB ;
wire  duc ;
wire  DUD ;
wire  due ;
wire  DUF ;
wire  dug ;
wire  dva ;
wire  DVB ;
wire  dvc ;
wire  DVD ;
wire  dve ;
wire  DVF ;
wire  dvg ;
wire  dwa ;
wire  DWB ;
wire  dwc ;
wire  DWD ;
wire  dwe ;
wire  DWF ;
wire  dwg ;
wire  dwh ;
wire  dxa ;
wire  DXB ;
wire  dxc ;
wire  DXD ;
wire  dxe ;
wire  DXF ;
wire  dxg ;
wire  dxh ;
wire  dya ;
wire  DYB ;
wire  dyc ;
wire  DYD ;
wire  dye ;
wire  DYF ;
wire  dyg ;
wire  DYH ;
wire  dza ;
wire  DZB ;
wire  dzc ;
wire  DZD ;
wire  dze ;
wire  DZF ;
wire  dzg ;
wire  DZH ;
wire  dzi ;
wire  DZJ ;
wire  dzk ;
wire  DZL ;
wire  dzm ;
wire  DZN ;
wire  dzo ;
wire  DZP ;
wire  dzq ;
wire  eaa ;
wire  EAA ;
wire  eba ;
wire  EBA ;
wire  eca ;
wire  ECA ;
wire  ecb ;
wire  ECB ;
wire  eda ;
wire  EDA ;
wire  edb ;
wire  EDB ;
wire  eea ;
wire  EEA ;
wire  efa ;
wire  EFA ;
wire  efb ;
wire  EFB ;
wire  eia ;
wire  EIA ;
wire  eib ;
wire  EIB ;
wire  eja ;
wire  EJA ;
wire  ejb ;
wire  EJB ;
wire  eka ;
wire  EKA ;
wire  ekb ;
wire  EKB ;
wire  ekc ;
wire  EKC ;
wire  ela ;
wire  ELA ;
wire  elb ;
wire  ELB ;
wire  elc ;
wire  ELC ;
wire  ema ;
wire  EMA ;
wire  emb ;
wire  EMB ;
wire  ena ;
wire  ENA ;
wire  enb ;
wire  ENB ;
wire  enc ;
wire  ENC ;
wire  eoa ;
wire  EOA ;
wire  eob ;
wire  EOB ;
wire  eoc ;
wire  EOC ;
wire  eod ;
wire  EOD ;
wire  epa ;
wire  EPA ;
wire  epb ;
wire  EPB ;
wire  epc ;
wire  EPC ;
wire  epd ;
wire  EPD ;
wire  eqa ;
wire  EQA ;
wire  eqb ;
wire  EQB ;
wire  eqc ;
wire  EQC ;
wire  eqd ;
wire  EQD ;
wire  era ;
wire  ERA ;
wire  erb ;
wire  ERB ;
wire  erc ;
wire  ERC ;
wire  erd ;
wire  ERD ;
wire  ere ;
wire  ERE ;
wire  esa ;
wire  ESA ;
wire  esb ;
wire  ESB ;
wire  esc ;
wire  ESC ;
wire  esd ;
wire  ESD ;
wire  eta ;
wire  ETA ;
wire  etb ;
wire  ETB ;
wire  etc ;
wire  ETC ;
wire  etd ;
wire  ETD ;
wire  eua ;
wire  EUA ;
wire  eub ;
wire  EUB ;
wire  euc ;
wire  EUC ;
wire  eud ;
wire  EUD ;
wire  eue ;
wire  EUE ;
wire  eva ;
wire  EVA ;
wire  evb ;
wire  EVB ;
wire  evc ;
wire  EVC ;
wire  evd ;
wire  EVD ;
wire  eve ;
wire  EVE ;
wire  evf ;
wire  EVF ;
wire  ewa ;
wire  EWA ;
wire  ewb ;
wire  EWB ;
wire  ewc ;
wire  EWC ;
wire  ewd ;
wire  EWD ;
wire  ewe ;
wire  EWE ;
wire  ewf ;
wire  EWF ;
wire  exa ;
wire  EXA ;
wire  exb ;
wire  EXB ;
wire  exc ;
wire  EXC ;
wire  exd ;
wire  EXD ;
wire  exe ;
wire  EXE ;
wire  exf ;
wire  EXF ;
wire  exg ;
wire  EXG ;
wire  exh ;
wire  EXH ;
wire  exi ;
wire  EXI ;
wire  exj ;
wire  EXJ ;
wire  exk ;
wire  EXK ;
wire  exl ;
wire  EXL ;
wire  exm ;
wire  EXM ;
wire  exn ;
wire  EXN ;
wire  exo ;
wire  EXO ;
wire  exp ;
wire  EXP ;
wire  exq ;
wire  EXQ ;
wire  exr ;
wire  EXR ;
wire  exs ;
wire  EXS ;
wire  ext ;
wire  EXT ;
wire  exu ;
wire  EXU ;
wire  eya ;
wire  EYA ;
wire  eyb ;
wire  EYB ;
wire  eyc ;
wire  EYC ;
wire  eyd ;
wire  EYD ;
wire  eye ;
wire  EYE ;
wire  eyf ;
wire  EYF ;
wire  eyg ;
wire  EYG ;
wire  eyh ;
wire  EYH ;
wire  eyi ;
wire  EYI ;
wire  eyj ;
wire  EYJ ;
wire  eyk ;
wire  EYK ;
wire  eyl ;
wire  EYL ;
wire  eym ;
wire  EYM ;
wire  eyn ;
wire  EYN ;
wire  eyo ;
wire  EYO ;
wire  eyp ;
wire  EYP ;
wire  eyq ;
wire  EYQ ;
wire  eyr ;
wire  EYR ;
wire  eys ;
wire  EYS ;
wire  eyt ;
wire  EYT ;
wire  eyu ;
wire  EYU ;
wire  eyv ;
wire  EYV ;
wire  eyw ;
wire  EYW ;
wire  eyx ;
wire  EYX ;
wire  eyy ;
wire  EYY ;
wire  eyz ;
wire  EYZ ;
wire  eza ;
wire  EZA ;
wire  ezb ;
wire  EZB ;
wire  ezc ;
wire  EZC ;
wire  ezd ;
wire  EZD ;
wire  eze ;
wire  EZE ;
wire  ezf ;
wire  EZF ;
wire  ezg ;
wire  EZG ;
wire  ezh ;
wire  EZH ;
wire  ezi ;
wire  EZI ;
wire  ezj ;
wire  EZJ ;
wire  ezk ;
wire  EZK ;
wire  ezl ;
wire  EZL ;
wire  ezm ;
wire  EZM ;
wire  ezn ;
wire  EZN ;
wire  ezo ;
wire  EZO ;
wire  ezp ;
wire  EZP ;
wire  ezq ;
wire  EZQ ;
wire  ezr ;
wire  EZR ;
wire  ezs ;
wire  EZS ;
wire  ezt ;
wire  EZT ;
wire  ezu ;
wire  EZU ;
wire  ezv ;
wire  EZV ;
wire  ezw ;
wire  EZW ;
wire  ezx ;
wire  EZX ;
wire  faa ;
wire  fba ;
wire  fca ;
wire  fcb ;
wire  fda ;
wire  fdb ;
wire  fea ;
wire  ffa ;
wire  ffb ;
wire  fga ;
wire  fha ;
wire  fhb ;
wire  fia ;
wire  FIB ;
wire  fja ;
wire  FJB ;
wire  fma ;
wire  fmb ;
wire  fna ;
wire  FNB ;
wire  foa ;
wire  FOB ;
wire  foc ;
wire  fpa ;
wire  FPB ;
wire  fpc ;
wire  fqa ;
wire  FQB ;
wire  fqc ;
wire  fra ;
wire  FRB ;
wire  frc ;
wire  frd ;
wire  fsa ;
wire  FSB ;
wire  fsc ;
wire  fsd ;
wire  fta ;
wire  FTB ;
wire  ftc ;
wire  fua ;
wire  FUB ;
wire  fuc ;
wire  fud ;
wire  fva ;
wire  FVB ;
wire  fvc ;
wire  FVD ;
wire  fwa ;
wire  FWB ;
wire  fwc ;
wire  fwd ;
wire  fxa ;
wire  FXB ;
wire  fxc ;
wire  FXD ;
wire  fxe ;
wire  fya ;
wire  FYB ;
wire  fyc ;
wire  fyd ;
wire  fye ;
wire  FYF ;
wire  fyg ;
wire  FYH ;
wire  fyi ;
wire  fyj ;
wire  FYK ;
wire  fyl ;
wire  FYM ;
wire  fyn ;
wire  fyo ;
wire  FYP ;
wire  fyq ;
wire  FYR ;
wire  fys ;
wire  fza ;
wire  FZB ;
wire  fzc ;
wire  FZD ;
wire  fze ;
wire  FZF ;
wire  fzg ;
wire  fzh ;
wire  fzi ;
wire  FZJ ;
wire  fzk ;
wire  FZL ;
wire  fzm ;
wire  FZN ;
wire  fzo ;
wire  FZP ;
wire  fzr ;
wire  FZS ;
wire  fzt ;
wire  FZU ;
wire  fzv ;
wire  fzw ;
wire  FZX ;
wire  fzy ;
wire  FZZ ;
wire  gma ;
wire  GMA ;
wire  gmb ;
wire  GMB ;
wire  gna ;
wire  GNA ;
wire  goa ;
wire  GOA ;
wire  gob ;
wire  GOB ;
wire  gpa ;
wire  GPA ;
wire  gpb ;
wire  GPB ;
wire  gqa ;
wire  GQA ;
wire  gqb ;
wire  GQB ;
wire  gra ;
wire  GRA ;
wire  grb ;
wire  GRB ;
wire  grc ;
wire  GRC ;
wire  gsa ;
wire  GSA ;
wire  gsb ;
wire  GSB ;
wire  gsc ;
wire  GSC ;
wire  gta ;
wire  GTA ;
wire  gtb ;
wire  GTB ;
wire  gua ;
wire  GUA ;
wire  gub ;
wire  GUB ;
wire  guc ;
wire  GUC ;
wire  gva ;
wire  GVA ;
wire  gvb ;
wire  GVB ;
wire  gvc ;
wire  GVC ;
wire  gwa ;
wire  GWA ;
wire  gwb ;
wire  GWB ;
wire  gwc ;
wire  GWC ;
wire  gwd ;
wire  GWD ;
wire  gxa ;
wire  GXA ;
wire  gxb ;
wire  GXB ;
wire  gxc ;
wire  GXC ;
wire  gya ;
wire  GYA ;
wire  gyb ;
wire  GYB ;
wire  gyc ;
wire  GYC ;
wire  gye ;
wire  GYE ;
wire  gyf ;
wire  GYF ;
wire  gyg ;
wire  GYG ;
wire  gyh ;
wire  GYH ;
wire  gyi ;
wire  GYI ;
wire  gyj ;
wire  GYJ ;
wire  gyl ;
wire  GYL ;
wire  gza ;
wire  GZA ;
wire  gzb ;
wire  GZB ;
wire  gzc ;
wire  GZC ;
wire  gzd ;
wire  GZD ;
wire  gze ;
wire  GZE ;
wire  gzf ;
wire  GZF ;
wire  gzg ;
wire  GZG ;
wire  gzh ;
wire  GZH ;
wire  gzi ;
wire  GZI ;
wire  gzj ;
wire  GZJ ;
wire  gzk ;
wire  gzm ;
wire  GZM ;
wire  gzn ;
wire  GZN ;
wire  gzo ;
wire  GZO ;
wire  gzp ;
wire  GZP ;
wire  gzq ;
wire  GZQ ;
wire  gzr ;
wire  GZR ;
wire  gzs ;
wire  GZS ;
wire  gzt ;
wire  GZT ;
wire  gzu ;
wire  GZU ;
wire  gzv ;
wire  GZV ;
wire  gzw ;
wire  GZW ;
wire  gzx ;
wire  GZX ;
wire  gzy ;
wire  GZY ;
wire  gzz ;
wire  GZZ ;
wire  haa ;
wire  hba ;
wire  hca ;
wire  hcb ;
wire  hda ;
wire  hdb ;
wire  hea ;
wire  hfa ;
wire  hfb ;
wire  hga ;
wire  hgb ;
wire  hha ;
wire  hhb ;
wire  hia ;
wire  hja ;
wire  hjb ;
wire  hma ;
wire  hna ;
wire  hnb ;
wire  hoa ;
wire  hpa ;
wire  hpb ;
wire  hqa ;
wire  hqb ;
wire  hra ;
wire  HRB ;
wire  hsa ;
wire  HSB ;
wire  hta ;
wire  htb ;
wire  hua ;
wire  HUB ;
wire  hva ;
wire  HVB ;
wire  hwa ;
wire  HWB ;
wire  hxa ;
wire  HXB ;
wire  hxc ;
wire  hya ;
wire  HYB ;
wire  hyd ;
wire  hza ;
wire  HZB ;
wire  hzc ;
wire  HZD ;
wire  hzg ;
wire  HZH ;
wire  hzi ;
wire  HZJ ;
wire  hzk ;
wire  hzm ;
wire  HZN ;
wire  hzo ;
wire  hzq ;
wire  HZR ;
wire  hzt ;
wire  HZU ;
wire  hzv ;
wire  hzw ;
wire  HZX ;
wire  hzy ;
wire  HZZ ;
wire  iaa ;
wire  iab ;
wire  iac ;
wire  iad ;
wire  iae ;
wire  iaf ;
wire  iag ;
wire  iah ;
wire  iai ;
wire  iaj ;
wire  iak ;
wire  ial ;
wire  iam ;
wire  ian ;
wire  iao ;
wire  iap ;
wire  iba ;
wire  ibb ;
wire  ibc ;
wire  ibd ;
wire  ibe ;
wire  ibf ;
wire  ibg ;
wire  ibh ;
wire  ibi ;
wire  ibj ;
wire  ibk ;
wire  ibl ;
wire  ibm ;
wire  ibn ;
wire  ibo ;
wire  ibp ;
wire  ica ;
wire  icb ;
wire  icc ;
wire  icd ;
wire  ice ;
wire  icf ;
wire  icg ;
wire  ich ;
wire  ici ;
wire  icj ;
wire  ick ;
wire  icl ;
wire  icm ;
wire  icn ;
wire  ico ;
wire  icp ;
wire  ida ;
wire  idb ;
wire  idc ;
wire  idd ;
wire  ide ;
wire  idf ;
wire  idg ;
wire  idh ;
wire  idi ;
wire  idj ;
wire  idk ;
wire  idl ;
wire  idm ;
wire  idn ;
wire  ido ;
wire  idp ;
wire  iea ;
wire  ieb ;
wire  iec ;
wire  ied ;
wire  iee ;
wire  ief ;
wire  ifa ;
wire  ifb ;
wire  ifc ;
wire  ifd ;
wire  ife ;
wire  iiff ;
wire  ifg ;
wire  iga ;
wire  igb ;
wire  igc ;
wire  igd ;
wire  ige ;
wire  igf ;
wire  iha ;
wire  jzt ;
wire  JZT ;
wire  jzu ;
wire  JZU ;
wire  jzy ;
wire  JZY ;
wire  jzz ;
wire  JZZ ;
wire  kaa ;
wire  kba ;
wire  kca ;
wire  kcb ;
wire  kda ;
wire  kdb ;
wire  kea ;
wire  kfa ;
wire  kga ;
wire  kha ;
wire  KHB ;
wire  kia ;
wire  kja ;
wire  kjb ;
wire  kma ;
wire  kna ;
wire  knb ;
wire  koa ;
wire  kpa ;
wire  kpb ;
wire  kqa ;
wire  kqb ;
wire  kra ;
wire  ksa ;
wire  ksb ;
wire  kta ;
wire  ktb ;
wire  kua ;
wire  kub ;
wire  kva ;
wire  kvb ;
wire  kwa ;
wire  kwb ;
wire  kxa ;
wire  KXB ;
wire  kya ;
wire  kyb ;
wire  kza ;
wire  kzb ;
wire  kzc ;
wire  kzd ;
wire  kzg ;
wire  kzh ;
wire  kzi ;
wire  KZJ ;
wire  kzm ;
wire  KZN ;
wire  kzq ;
wire  kzr ;
wire  kzt ;
wire  kzw ;
wire  kzx ;
wire  kzy ;
wire  laa ;
wire  LAA ;
wire  lba ;
wire  LBA ;
wire  lbb ;
wire  LBB ;
wire  lca ;
wire  LCA ;
wire  lcb ;
wire  LCB ;
wire  lda ;
wire  LDA ;
wire  ldb ;
wire  LDB ;
wire  ldc ;
wire  LDC ;
wire  lea ;
wire  LEA ;
wire  leb ;
wire  LEB ;
wire  lfa ;
wire  LFA ;
wire  lfb ;
wire  LFB ;
wire  lfc ;
wire  LFC ;
wire  lga ;
wire  LGA ;
wire  lgb ;
wire  LGB ;
wire  lha ;
wire  LHA ;
wire  lhb ;
wire  LHB ;
wire  lia ;
wire  LIA ;
wire  lib ;
wire  LIB ;
wire  lic ;
wire  LIC ;
wire  lid ;
wire  LID ;
wire  lja ;
wire  LJA ;
wire  ljb ;
wire  LJB ;
wire  lka ;
wire  LKA ;
wire  lkb ;
wire  LKB ;
wire  lla ;
wire  LLA ;
wire  llb ;
wire  LLB ;
wire  lma ;
wire  LMA ;
wire  lmb ;
wire  LMB ;
wire  lna ;
wire  LNA ;
wire  lnb ;
wire  LNB ;
wire  loa ;
wire  LOA ;
wire  lob ;
wire  LOB ;
wire  loc ;
wire  LOC ;
wire  lqa ;
wire  LQA ;
wire  lqb ;
wire  LQB ;
wire  lra ;
wire  LRA ;
wire  lrb ;
wire  LRB ;
wire  lsa ;
wire  LSA ;
wire  lsb ;
wire  LSB ;
wire  lsc ;
wire  LSC ;
wire  lta ;
wire  LTA ;
wire  ltb ;
wire  LTB ;
wire  ltc ;
wire  LTC ;
wire  lua ;
wire  LUA ;
wire  lub ;
wire  LUB ;
wire  luc ;
wire  LUC ;
wire  lva ;
wire  LVA ;
wire  lvb ;
wire  LVB ;
wire  lvc ;
wire  LVC ;
wire  lwa ;
wire  LWA ;
wire  lwb ;
wire  LWB ;
wire  lwc ;
wire  LWC ;
wire  lxa ;
wire  LXA ;
wire  lxb ;
wire  LXB ;
wire  lxc ;
wire  LXC ;
wire  lya ;
wire  LYA ;
wire  lyb ;
wire  LYB ;
wire  lyc ;
wire  LYC ;
wire  lza ;
wire  LZA ;
wire  lzb ;
wire  LZB ;
wire  lzc ;
wire  LZC ;
wire  lzd ;
wire  LZD ;
wire  lze ;
wire  LZE ;
wire  lzf ;
wire  LZF ;
wire  lzi ;
wire  LZI ;
wire  lzj ;
wire  LZJ ;
wire  lzk ;
wire  LZK ;
wire  lzl ;
wire  LZL ;
wire  lzm ;
wire  LZM ;
wire  lzn ;
wire  LZN ;
wire  lzo ;
wire  LZO ;
wire  lzp ;
wire  LZP ;
wire  lzq ;
wire  LZQ ;
wire  lzr ;
wire  LZR ;
wire  lzs ;
wire  LZS ;
wire  lzt ;
wire  LZT ;
wire  lzu ;
wire  LZU ;
wire  lzv ;
wire  LZV ;
wire  lzw ;
wire  LZW ;
wire  lzx ;
wire  LZX ;
wire  lzy ;
wire  LZY ;
wire  lzz ;
wire  LZZ ;
wire  maa ;
wire  mba ;
wire  mbb ;
wire  mca ;
wire  mda ;
wire  MDB ;
wire  mea ;
wire  meb ;
wire  mfa ;
wire  mfb ;
wire  mga ;
wire  mgb ;
wire  mha ;
wire  mhb ;
wire  mia ;
wire  MIB ;
wire  mja ;
wire  MJB ;
wire  mka ;
wire  mkb ;
wire  mla ;
wire  mlb ;
wire  mma ;
wire  mmb ;
wire  mna ;
wire  mnb ;
wire  moa ;
wire  MOB ;
wire  mqa ;
wire  mqb ;
wire  mra ;
wire  mrb ;
wire  msa ;
wire  MSB ;
wire  mta ;
wire  MTB ;
wire  mua ;
wire  MUB ;
wire  mva ;
wire  MVB ;
wire  mwa ;
wire  MWB ;
wire  mxa ;
wire  MXB ;
wire  mya ;
wire  MYB ;
wire  mza ;
wire  MZB ;
wire  mzd ;
wire  MZE ;
wire  mzi ;
wire  MZJ ;
wire  mzl ;
wire  MZM ;
wire  mzo ;
wire  MZP ;
wire  mzr ;
wire  MZS ;
wire  mzu ;
wire  MZV ;
wire  mzx ;
wire  MZY ;
wire  naa ;
wire  nab ;
wire  nac ;
wire  nad ;
wire  nae ;
wire  naf ;
wire  nag ;
wire  nah ;
wire  nai ;
wire  naj ;
wire  nak ;
wire  nal ;
wire  nam ;
wire  nan ;
wire  nao ;
wire  nap ;
wire  naq ;
wire  nba ;
wire  nbb ;
wire  nbc ;
wire  nbd ;
wire  nbe ;
wire  nbf ;
wire  nbg ;
wire  nbh ;
wire  nbi ;
wire  nbj ;
wire  nbk ;
wire  nbl ;
wire  nbm ;
wire  nbn ;
wire  nbo ;
wire  nbp ;
wire  neb ;
wire  nee ;
wire  nef ;
wire  neg ;
wire  neh ;
wire  nei ;
wire  nej ;
wire  nek ;
wire  nel ;
wire  nem ;
wire  nen ;
wire  neo ;
wire  nep ;
wire  nfb ;
wire  nfc ;
wire  nfd ;
wire  nfe ;
wire  nff ;
wire  nfg ;
wire  nfh ;
wire  nfi ;
wire  nfj ;
wire  nfk ;
wire  nfl ;
wire  nfm ;
wire  nfn ;
wire  nfo ;
wire  nfp ;
wire  ngd ;
wire  NGD ;
wire  nge ;
wire  NGE ;
wire  nhb ;
wire  NHB ;
wire  nhc ;
wire  NHC ;
wire  nhd ;
wire  NHD ;
wire  nhe ;
wire  NHE ;
wire  nib ;
wire  NIB ;
wire  nic ;
wire  NIC ;
wire  nid ;
wire  NID ;
wire  nie ;
wire  NIE ;
wire  njb ;
wire  NJB ;
wire  njc ;
wire  NJC ;
wire  njd ;
wire  NJD ;
wire  nje ;
wire  NJE ;
wire  nkb ;
wire  NKB ;
wire  nkc ;
wire  NKC ;
wire  nkd ;
wire  NKD ;
wire  nke ;
wire  NKE ;
wire  nlb ;
wire  NLB ;
wire  nlc ;
wire  NLC ;
wire  nld ;
wire  NLD ;
wire  nle ;
wire  NLE ;
wire  nmb ;
wire  NMB ;
wire  nmc ;
wire  NMC ;
wire  nmd ;
wire  NMD ;
wire  nme ;
wire  NME ;
wire  nnb ;
wire  NNB ;
wire  nnc ;
wire  NNC ;
wire  nnd ;
wire  NND ;
wire  nne ;
wire  NNE ;
wire  npb ;
wire  NPB ;
wire  npc ;
wire  NPC ;
wire  npd ;
wire  NPD ;
wire  nqb ;
wire  NQB ;
wire  nqc ;
wire  NQC ;
wire  nqd ;
wire  NQD ;
wire  nrb ;
wire  NRB ;
wire  nrc ;
wire  NRC ;
wire  nrd ;
wire  NRD ;
wire  nsb ;
wire  NSB ;
wire  nsc ;
wire  NSC ;
wire  nsd ;
wire  NSD ;
wire  ntb ;
wire  NTB ;
wire  ntc ;
wire  NTC ;
wire  ntd ;
wire  NTD ;
wire  nub ;
wire  NUB ;
wire  nuc ;
wire  NUC ;
wire  nud ;
wire  NUD ;
wire  nvb ;
wire  NVB ;
wire  nvc ;
wire  NVC ;
wire  nvd ;
wire  NVD ;
wire  nxb ;
wire  NXB ;
wire  nxc ;
wire  NXC ;
wire  nxd ;
wire  NXD ;
wire  nxe ;
wire  NXE ;
wire  nxf ;
wire  NXF ;
wire  nxg ;
wire  NXG ;
wire  nxi ;
wire  NXI ;
wire  nxj ;
wire  NXJ ;
wire  nxk ;
wire  NXK ;
wire  nxl ;
wire  NXL ;
wire  oaa ;
wire  oab ;
wire  oac ;
wire  oad ;
wire  oae ;
wire  oaf ;
wire  oag ;
wire  oah ;
wire  oai ;
wire  oaj ;
wire  oak ;
wire  oal ;
wire  oam ;
wire  oan ;
wire  oao ;
wire  oap ;
wire  oba ;
wire  obb ;
wire  obc ;
wire  obd ;
wire  obe ;
wire  obf ;
wire  obg ;
wire  obh ;
wire  obi ;
wire  obj ;
wire  obk ;
wire  obl ;
wire  obm ;
wire  obn ;
wire  obo ;
wire  obp ;
wire  oea ;
wire  oeb ;
wire  oec ;
wire  oed ;
wire  oee ;
wire  oef ;
wire  ofa ;
wire  ofb ;
wire  ofc ;
wire  ofd ;
wire  ofe ;
wire  off ;
wire  OGA ;
wire  OGB ;
wire  OGC ;
wire  OGD ;
wire  OGE ;
wire  OGF ;
wire  OHA ;
wire  OHB ;
wire  OHC ;
wire  OHD ;
wire  OHE ;
wire  OHF ;
wire  OIA ;
wire  OIB ;
wire  OIC ;
wire  OID ;
wire  OIE ;
wire  OIF ;
wire  OIG ;
wire  OIH ;
wire  OII ;
wire  OIJ ;
wire  OIK ;
wire  OIL ;
wire  OIM ;
wire  oja ;
wire  ojb ;
wire  ojc ;
wire  ojd ;
wire  oje ;
wire  ojf ;
wire  ojg ;
wire  ojh ;
wire  oji ;
wire  ojj ;
wire  ojk ;
wire  ojl ;
wire  ojm ;
wire  OKA ;
wire  OKB ;
wire  OKC ;
wire  OKD ;
wire  OKE ;
wire  OKF ;
wire  OKG ;
wire  OKH ;
wire  OKI ;
wire  OKJ ;
wire  OKK ;
wire  OKL ;
wire  OKM ;
wire  ola ;
wire  olb ;
wire  olc ;
wire  old ;
wire  ole ;
wire  olf ;
wire  olg ;
wire  olh ;
wire  oli ;
wire  olj ;
wire  olk ;
wire  oll ;
wire  olm ;
wire  OMA ;
wire  OMB ;
wire  OMC ;
wire  OMD ;
wire  OME ;
wire  OMF ;
wire  OMG ;
wire  OMH ;
wire  OMI ;
wire  OMJ ;
wire  OMK ;
wire  OML ;
wire  OMM ;
wire  ona ;
wire  onb ;
wire  onc ;
wire  ond ;
wire  one ;
wire  onf ;
wire  ong ;
wire  onh ;
wire  oni ;
wire  onj ;
wire  onk ;
wire  onl ;
wire  onm ;
wire  OOA ;
wire  OOB ;
wire  OOC ;
wire  OOD ;
wire  OOE ;
wire  OOF ;
wire  OOG ;
wire  OOH ;
wire  OOI ;
wire  OOJ ;
wire  OOK ;
wire  OOL ;
wire  OOM ;
wire  opa ;
wire  opb ;
wire  opc ;
wire  opd ;
wire  ope ;
wire  opf ;
wire  opg ;
wire  oph ;
wire  opi ;
wire  opj ;
wire  opk ;
wire  opl ;
wire  opm ;
wire  pab ;
wire  pac ;
wire  pad ;
wire  pae ;
wire  paf ;
wire  pag ;
wire  pah ;
wire  PAI ;
wire  PAK ;
wire  pal ;
wire  pam ;
wire  PAM ;
wire  pao ;
wire  pap ;
wire  PAP ;
wire  paq ;
wire  pba ;
wire  pbb ;
wire  pbc ;
wire  pbd ;
wire  pbe ;
wire  pbf ;
wire  pbg ;
wire  pbh ;
wire  pbi ;
wire  pbj ;
wire  pbk ;
wire  pbl ;
wire  pbm ;
wire  pbn ;
wire  pbo ;
wire  pbp ;
wire  pca ;
wire  pcb ;
wire  pcc ;
wire  pcd ;
wire  pce ;
wire  pcf ;
wire  pcg ;
wire  pch ;
wire  pci ;
wire  pcj ;
wire  pck ;
wire  pcl ;
wire  pcm ;
wire  pcn ;
wire  pco ;
wire  pcp ;
wire  pde ;
wire  pdf ;
wire  pdg ;
wire  pdh ;
wire  pdi ;
wire  pdj ;
wire  pdk ;
wire  pdl ;
wire  pdm ;
wire  pdn ;
wire  pdo ;
wire  pdp ;
wire  pea ;
wire  peb ;
wire  pec ;
wire  ped ;
wire  pee ;
wire  pef ;
wire  peg ;
wire  peh ;
wire  pei ;
wire  pej ;
wire  pek ;
wire  pel ;
wire  pem ;
wire  pen ;
wire  peo ;
wire  pep ;
wire  pfa ;
wire  pfb ;
wire  pfc ;
wire  pfd ;
wire  pfe ;
wire  pff ;
wire  pfg ;
wire  pfh ;
wire  pfi ;
wire  pfj ;
wire  pfk ;
wire  pfl ;
wire  pfm ;
wire  pfn ;
wire  pfo ;
wire  pfp ;
wire  pga ;
wire  pgb ;
wire  pgc ;
wire  pgd ;
wire  pge ;
wire  pgf ;
wire  pgg ;
wire  pgh ;
wire  pgi ;
wire  pgj ;
wire  pgk ;
wire  pgl ;
wire  pgm ;
wire  pgn ;
wire  pgo ;
wire  pgp ;
wire  qaa ;
wire  qab ;
wire  qac ;
wire  qad ;
wire  qae ;
wire  qaf ;
wire  qag ;
wire  qah ;
wire  qai ;
wire  qaj ;
wire  qak ;
wire  qal ;
wire  QVA ;
wire  qvb ;
wire  QVC ;
wire  qvd ;
wire  QVE ;
wire  qvf ;
wire  qvg ;
wire  qxa ;
wire  QXB ;
wire  qxc ;
wire  QXD ;
wire  qxe ;
wire  QXF ;
wire  qxg ;
wire  QXH ;
wire  qxi ;
wire  QXJ ;
wire  qxk ;
wire  QXL ;
wire  qxm ;
wire  QXN ;
wire  qxo ;
wire  QXP ;
wire  qxq ;
wire  QXR ;
wire  qxs ;
wire  QXT ;
wire  qxu ;
wire  qxv ;
wire  QXW ;
wire  qxx ;
wire  QXY ;
wire  qxz ;
wire  qya ;
wire  QYB ;
wire  qyc ;
wire  QYD ;
wire  qye ;
wire  QYF ;
wire  qyg ;
wire  QYH ;
wire  qyi ;
wire  qyj ;
wire  QYK ;
wire  qyl ;
wire  QYM ;
wire  qyn ;
wire  QYO ;
wire  qyp ;
wire  QYQ ;
wire  qyr ;
wire  qys ;
wire  qza ;
wire  QZB ;
wire  qzc ;
wire  QZD ;
wire  qze ;
wire  QZF ;
wire  qzg ;
wire  QZH ;
wire  qzi ;
wire  qzj ;
wire  qzk ;
wire  QZL ;
wire  qzm ;
wire  QZN ;
wire  qzo ;
wire  QZP ;
wire  qzq ;
wire  QZR ;
wire  qzs ;
wire  QZT ;
wire  rae ;
wire  RAE ;
wire  raf ;
wire  RAF ;
wire  rag ;
wire  RAG ;
wire  rah ;
wire  RAH ;
wire  rai ;
wire  RAI ;
wire  raj ;
wire  RAJ ;
wire  rak ;
wire  RAK ;
wire  ral ;
wire  RAL ;
wire  ram ;
wire  RAM ;
wire  ran ;
wire  RAN ;
wire  rao ;
wire  RAO ;
wire  rap ;
wire  RAP ;
wire  rba ;
wire  RBA ;
wire  rbb ;
wire  RBB ;
wire  rbc ;
wire  RBC ;
wire  rbd ;
wire  RBD ;
wire  rbe ;
wire  RBE ;
wire  rbf ;
wire  RBF ;
wire  rbg ;
wire  RBG ;
wire  rbh ;
wire  RBH ;
wire  rbi ;
wire  RBI ;
wire  rbj ;
wire  RBJ ;
wire  rbk ;
wire  RBK ;
wire  rbl ;
wire  RBL ;
wire  rbm ;
wire  RBM ;
wire  rbn ;
wire  RBN ;
wire  rbo ;
wire  RBO ;
wire  rbp ;
wire  RBP ;
wire  tea ;
wire  TEA ;
wire  teb ;
wire  TEB ;
wire  tec ;
wire  TEC ;
wire  ted ;
wire  TED ;
wire  tee ;
wire  TEE ;
wire  tef ;
wire  TEF ;
wire  teg ;
wire  TEG ;
wire  teh ;
wire  TEH ;
wire  tfa ;
wire  tfb ;
wire  tfc ;
wire  tfd ;
wire  ZZI ;
wire  ZZO ;
assign ZZI = 1'b1;
assign ZZO = 1'b0;
assign aal = ~AAL;  //complement 
assign aam = ~AAM;  //complement 
assign aan = ~AAN;  //complement 
assign aao = ~AAO;  //complement 
assign aap = ~AAP;  //complement 
assign RAO =  NAO & neo  ; 
assign rao = ~RAO;  //complement 
assign RAP =  NAP & nep  ; 
assign rap = ~RAP;  //complement 
assign LUC =  KUB  ; 
assign luc = ~LUC;  //complement 
assign dhb = ~DHB;  //complement 
assign qxu = ~QXU;  //complement 
assign ftc = ~FTC;  //complement 
assign pao = ~PAO;  //complement 
assign dhc = ~DHC;  //complement 
assign dhd = ~DHD;  //complement 
assign dkc = ~DKC;  //complement 
assign dkd = ~DKD;  //complement 
assign ojg = ~OJG;  //complement 
assign olg = ~OLG;  //complement 
assign ong = ~ONG;  //complement 
assign opg = ~OPG;  //complement 
assign neb = ~NEB;  //complement 
assign dic = ~DIC;  //complement 
assign DID = ~did;  //complement 
assign dha = ~DHA;  //complement 
assign fyn = ~FYN;  //complement 
assign kcb = ~KCB;  //complement 
assign kdb = ~KDB;  //complement 
assign dga = ~DGA;  //complement 
assign dgb = ~DGB;  //complement 
assign dpe = ~DPE;  //complement 
assign qyi = ~QYI;  //complement 
assign nbc = ~NBC;  //complement 
assign dja = ~DJA;  //complement 
assign DJB = ~djb;  //complement 
assign fza = ~FZA;  //complement 
assign FZB = ~fzb;  //complement 
assign EXE =  DXH  ; 
assign exe = ~EXE;  //complement 
assign EDA =  DHC  ; 
assign eda = ~EDA;  //complement 
assign EFA =  DIA  ; 
assign efa = ~EFA;  //complement 
assign nbb = ~NBB;  //complement 
assign dka = ~DKA;  //complement 
assign DKB = ~dkb;  //complement 
assign dwg = ~DWG;  //complement 
assign dwh = ~DWH;  //complement 
assign dxg = ~DXG;  //complement 
assign dxh = ~DXH;  //complement 
assign die = ~DIE;  //complement 
assign djc = ~DJC;  //complement 
assign dug = ~DUG;  //complement 
assign hea = ~HEA;  //complement 
assign mda = ~MDA;  //complement 
assign MDB = ~mdb;  //complement 
assign dla = ~DLA;  //complement 
assign DLB = ~dlb;  //complement 
assign nfp = ~NFP;  //complement 
assign EZG =  DZI & dzb & dzk  |  dzi & DZB & dzk  |  dzi & dzb & DZK  |  DZI & DZB & DZK  ; 
assign ezg = ~EZG; //complement 
assign ezh =  DZI & dzb & dzk  |  dzi & DZB & dzk  |  dzi & dzb & DZK  |  dzi & dzb & dzk  ; 
assign EZH = ~ezh;  //complement 
assign mzx = ~MZX;  //complement 
assign MZY = ~mzy;  //complement 
assign dma = ~DMA;  //complement 
assign DMB = ~dmb;  //complement 
assign aaa = ~AAA;  //complement 
assign aab = ~AAB;  //complement 
assign aac = ~AAC;  //complement 
assign aad = ~AAD;  //complement 
assign aae = ~AAE;  //complement 
assign aaf = ~AAF;  //complement 
assign RAI =  NAI & nei  ; 
assign rai = ~RAI;  //complement 
assign RAJ =  NAJ & nej  ; 
assign raj = ~RAJ;  //complement 
assign RAK =  NAK & nek  ; 
assign rak = ~RAK;  //complement 
assign aag = ~AAG;  //complement 
assign aah = ~AAH;  //complement 
assign aai = ~AAI;  //complement 
assign aaj = ~AAJ;  //complement 
assign aak = ~AAK;  //complement 
assign RAL =  NAL & nel  ; 
assign ral = ~RAL;  //complement 
assign RAM =  NAM & nem  ; 
assign ram = ~RAM;  //complement 
assign RAN =  NAN & nen  ; 
assign ran = ~RAN;  //complement 
assign dhe = ~DHE;  //complement 
assign DHF = ~dhf;  //complement 
assign dia = ~DIA;  //complement 
assign DIB = ~dib;  //complement 
assign dnc = ~DNC;  //complement 
assign DND = ~dnd;  //complement 
assign abg = ~ABG;  //complement 
assign abh = ~ABH;  //complement 
assign EYO =  QZO & qzq & qzd  |  qzo & QZQ & qzd  |  qzo & qzq & QZD  |  QZO & QZQ & QZD  ; 
assign eyo = ~EYO; //complement 
assign eyp =  QZO & qzq & qzd  |  qzo & QZQ & qzd  |  qzo & qzq & QZD  |  qzo & qzq & qzd  ; 
assign EYP = ~eyp;  //complement 
assign EYQ =  QZS & qzf & qzh  |  qzs & QZF & qzh  |  qzs & qzf & QZH  |  QZS & QZF & QZH  ; 
assign eyq = ~EYQ; //complement 
assign eyr =  QZS & qzf & qzh  |  qzs & QZF & qzh  |  qzs & qzf & QZH  |  qzs & qzf & qzh  ; 
assign EYR = ~eyr;  //complement 
assign doa = ~DOA;  //complement 
assign DOB = ~dob;  //complement 
assign abi = ~ABI;  //complement 
assign abj = ~ABJ;  //complement 
assign abk = ~ABK;  //complement 
assign hja = ~HJA;  //complement 
assign hia = ~HIA;  //complement 
assign hma = ~HMA;  //complement 
assign mba = ~MBA;  //complement 
assign EYU =  QXE & qxg & qzn  |  qxe & QXG & qzn  |  qxe & qxg & QZN  |  QXE & QXG & QZN  ; 
assign eyu = ~EYU; //complement 
assign eyv =  QXE & qxg & qzn  |  qxe & QXG & qzn  |  qxe & qxg & QZN  |  qxe & qxg & qzn  ; 
assign EYV = ~eyv;  //complement 
assign doc = ~DOC;  //complement 
assign DOD = ~dod;  //complement 
assign abl = ~ABL;  //complement 
assign abm = ~ABM;  //complement 
assign abn = ~ABN;  //complement 
assign EYW =  QZP & qzr & qzt  |  qzp & QZR & qzt  |  qzp & qzr & QZT  |  QZP & QZR & QZT  ; 
assign eyw = ~EYW; //complement 
assign eyx =  QZP & qzr & qzt  |  qzp & QZR & qzt  |  qzp & qzr & QZT  |  qzp & qzr & qzt  ; 
assign EYX = ~eyx;  //complement 
assign EZA =  DZA & dyb & dzc  |  dza & DYB & dzc  |  dza & dyb & DZC  |  DZA & DYB & DZC  ; 
assign eza = ~EZA; //complement 
assign ezb =  DZA & dyb & dzc  |  dza & DYB & dzc  |  dza & dyb & DZC  |  dza & dyb & dzc  ; 
assign EZB = ~ezb;  //complement 
assign dpa = ~DPA;  //complement 
assign DPB = ~dpb;  //complement 
assign abo = ~ABO;  //complement 
assign abp = ~ABP;  //complement 
assign EZC =  DZE & dzg & dyd  |  dze & DZG & dyd  |  dze & dzg & DYD  |  DZE & DZG & DYD  ; 
assign ezc = ~EZC; //complement 
assign ezd =  DZE & dzg & dyd  |  dze & DZG & dyd  |  dze & dzg & DYD  |  dze & dzg & dyd  ; 
assign EZD = ~ezd;  //complement 
assign EZE =  DYF  ; 
assign eze = ~EZE;  //complement 
assign EZF =  DYH  ; 
assign ezf = ~EZF;  //complement 
assign LAA =  KAA  ; 
assign laa = ~LAA;  //complement 
assign dpc = ~DPC;  //complement 
assign DPD = ~dpd;  //complement 
assign EZO =  QYE & qyg & dzl  |  qye & QYG & dzl  |  qye & qyg & DZL  |  QYE & QYG & DZL  ; 
assign ezo = ~EZO; //complement 
assign ezp =  QYE & qyg & dzl  |  qye & QYG & dzl  |  qye & qyg & DZL  |  qye & qyg & dzl  ; 
assign EZP = ~ezp;  //complement 
assign EZI =  DZM & dzo & dzd  |  dzm & DZO & dzd  |  dzm & dzo & DZD  |  DZM & DZO & DZD  ; 
assign ezi = ~EZI; //complement 
assign ezj =  DZM & dzo & dzd  |  dzm & DZO & dzd  |  dzm & dzo & DZD  |  dzm & dzo & dzd  ; 
assign EZJ = ~ezj;  //complement 
assign EZK =  DZQ & dzf & dzh  |  dzq & DZF & dzh  |  dzq & dzf & DZH  |  DZQ & DZF & DZH  ; 
assign ezk = ~EZK; //complement 
assign ezl =  DZQ & dzf & dzh  |  dzq & DZF & dzh  |  dzq & dzf & DZH  |  dzq & dzf & dzh  ; 
assign EZL = ~ezl;  //complement 
assign dqa = ~DQA;  //complement 
assign DQB = ~dqb;  //complement 
assign faa = ~FAA;  //complement 
assign fba = ~FBA;  //complement 
assign fca = ~FCA;  //complement 
assign fda = ~FDA;  //complement 
assign EZM =  QYA & qyc & dzj  |  qya & QYC & dzj  |  qya & qyc & DZJ  |  QYA & QYC & DZJ  ; 
assign ezm = ~EZM; //complement 
assign ezn =  QYA & qyc & dzj  |  qya & QYC & dzj  |  qya & qyc & DZJ  |  qya & qyc & dzj  ; 
assign EZN = ~ezn;  //complement 
assign EZQ =  QYI & dzn & dzp  |  qyi & DZN & dzp  |  qyi & dzn & DZP  |  QYI & DZN & DZP  ; 
assign ezq = ~EZQ; //complement 
assign ezr =  QYI & dzn & dzp  |  qyi & DZN & dzp  |  qyi & dzn & DZP  |  qyi & dzn & dzp  ; 
assign EZR = ~ezr;  //complement 
assign dmc = ~DMC;  //complement 
assign DMD = ~dmd;  //complement 
assign aba = ~ABA;  //complement 
assign abb = ~ABB;  //complement 
assign abc = ~ABC;  //complement 
assign LID =  HGB & KHB  ; 
assign lid = ~LID;  //complement 
assign GZF =  FZD & FZH  ; 
assign gzf = ~GZF;  //complement 
assign EYZ =  QXJ & QXO  ; 
assign eyz = ~EYZ;  //complement 
assign dna = ~DNA;  //complement 
assign DNB = ~dnb;  //complement 
assign abd = ~ABD;  //complement 
assign abe = ~ABE;  //complement 
assign abf = ~ABF;  //complement 
assign EYJ =  QZI & qys & qyo  |  qzi & QYS & qyo  |  qzi & qys & QYO  |  QZI & QYS & QYO  ; 
assign eyj = ~EYJ; //complement 
assign eyk =  QZI & qys & qyo  |  qzi & QYS & qyo  |  qzi & qys & QYO  |  qzi & qys & qyo  ; 
assign EYK = ~eyk;  //complement 
assign EYM =  QZK & qzm & qzb  |  qzk & QZM & qzb  |  qzk & qzm & QZB  |  QZK & QZM & QZB  ; 
assign eym = ~EYM; //complement 
assign eyn =  QZK & qzm & qzb  |  qzk & QZM & qzb  |  qzk & qzm & QZB  |  qzk & qzm & qzb  ; 
assign EYN = ~eyn;  //complement 
assign CAA = BAA & ACA ; 
assign caa = ~CAA ; //complement 
assign CAB = BAA & ACC ; 
assign cab = ~CAB ;  //complement 
assign CAC = BAA & ACE ; 
assign cac = ~CAC ;  //complement 
assign CAD = BAA & ACG; 
assign cad = ~CAD; 
assign CPB =  BAP & ACD  ; 
assign cpb = ~CPB;  //complement 
assign CPC =  BAP & ACF  ; 
assign cpc = ~CPC;  //complement 
assign CPD =  BAP & ACH  ; 
assign cpd = ~CPD;  //complement 
assign baa = ~BAA;  //complement 
assign bab = ~BAB;  //complement 
assign bac = ~BAC;  //complement 
assign oaa = ~OAA;  //complement 
assign oab = ~OAB;  //complement 
assign oac = ~OAC;  //complement 
assign CAE = BAA & ACI ; 
assign cae = ~CAE ; //complement 
assign CAF = BAA & ACK ; 
assign caf = ~CAF ;  //complement 
assign CAG = BAA & ACM ; 
assign cag = ~CAG ;  //complement 
assign CAH = BAA & ACO; 
assign cah = ~CAH; 
assign CPE =  BAP & ACJ  ; 
assign cpe = ~CPE;  //complement 
assign CPF =  BAP & ACL  ; 
assign cpf = ~CPF;  //complement 
assign CPG =  BAP & ACN  ; 
assign cpg = ~CPG;  //complement 
assign bad = ~BAD;  //complement 
assign bae = ~BAE;  //complement 
assign baf = ~BAF;  //complement 
assign oad = ~OAD;  //complement 
assign oae = ~OAE;  //complement 
assign oaf = ~OAF;  //complement 
assign CAI = BAA & ADA ; 
assign cai = ~CAI ; //complement 
assign CAJ = BAA & ADC ; 
assign caj = ~CAJ ;  //complement 
assign CAK = BAA & ADE ; 
assign cak = ~CAK ;  //complement 
assign CAL = BAA & ADG; 
assign cal = ~CAL; 
assign CPH =  BAP & ACP  ; 
assign cph = ~CPH;  //complement 
assign CPI =  BAP & ADB  ; 
assign cpi = ~CPI;  //complement 
assign CQA =  BBA & ACA  ; 
assign cqa = ~CQA;  //complement 
assign bai = ~BAI;  //complement 
assign baj = ~BAJ;  //complement 
assign bak = ~BAK;  //complement 
assign oag = ~OAG;  //complement 
assign oah = ~OAH;  //complement 
assign GUC =  FUD  ; 
assign guc = ~GUC;  //complement 
assign GVC =  ZZO  ; 
assign gvc = ~GVC;  //complement 
assign GYJ =  ZZO  ; 
assign gyj = ~GYJ;  //complement 
assign CQB =  BBA & ACC  ; 
assign cqb = ~CQB;  //complement 
assign CQC =  BBA & ACE  ; 
assign cqc = ~CQC;  //complement 
assign CQD =  BBA & ACG  ; 
assign cqd = ~CQD;  //complement 
assign bal = ~BAL;  //complement 
assign bam = ~BAM;  //complement 
assign ban = ~BAN;  //complement 
assign oai = ~OAI;  //complement 
assign oaj = ~OAJ;  //complement 
assign oak = ~OAK;  //complement 
assign CAM = BAA & ADI ; 
assign cam = ~CAM ; //complement 
assign CAN = BAA & ADK ; 
assign can = ~CAN ;  //complement 
assign CAO = BAA & ADM ; 
assign cao = ~CAO ;  //complement 
assign CAP = BAA & ADO; 
assign cap = ~CAP; 
assign CQE =  BBA & ACI  ; 
assign cqe = ~CQE;  //complement 
assign CQF =  BBA & ACK  ; 
assign cqf = ~CQF;  //complement 
assign CQG =  BBA & ACM  ; 
assign cqg = ~CQG;  //complement 
assign bbi = ~BBI;  //complement 
assign bbj = ~BBJ;  //complement 
assign bbk = ~BBK;  //complement 
assign oal = ~OAL;  //complement 
assign oam = ~OAM;  //complement 
assign oan = ~OAN;  //complement 
assign CBA = BAB & ACB ; 
assign cba = ~CBA ; //complement 
assign CBB = BAB & ACD ; 
assign cbb = ~CBB ;  //complement 
assign CBC = BAB & ACF ; 
assign cbc = ~CBC ;  //complement 
assign CBD = BAB & ACH; 
assign cbd = ~CBD; 
assign CQH =  BBA & ACO  ; 
assign cqh = ~CQH;  //complement 
assign CRA =  BBB & ACB  ; 
assign cra = ~CRA;  //complement 
assign CRB =  BBB & ACD  ; 
assign crb = ~CRB;  //complement 
assign bbl = ~BBL;  //complement 
assign bbm = ~BBM;  //complement 
assign bbn = ~BBN;  //complement 
assign oao = ~OAO;  //complement 
assign oap = ~OAP;  //complement 
assign knb = ~KNB;  //complement 
assign kjb = ~KJB;  //complement 
assign paq = ~PAQ;  //complement 
assign CRC =  BBB & ACF  ; 
assign crc = ~CRC;  //complement 
assign CRD =  BBB & ACH  ; 
assign crd = ~CRD;  //complement 
assign CRE =  BBB & ACJ  ; 
assign cre = ~CRE;  //complement 
assign doe = ~DOE;  //complement 
assign pal = ~PAL;  //complement 
assign fpc = ~FPC;  //complement 
assign fga = ~FGA;  //complement 
assign oba = ~OBA;  //complement 
assign obb = ~OBB;  //complement 
assign obc = ~OBC;  //complement 
assign CBE = BAB & ACJ ; 
assign cbe = ~CBE ; //complement 
assign CBF = BAB & ACL ; 
assign cbf = ~CBF ;  //complement 
assign CBG = BAB & ACN ; 
assign cbg = ~CBG ;  //complement 
assign CBH = BAB & ACP; 
assign cbh = ~CBH; 
assign CRF =  BBB & ACL  ; 
assign crf = ~CRF;  //complement 
assign CRG =  BBB & ACN  ; 
assign crg = ~CRG;  //complement 
assign CRH =  BBB & ACP  ; 
assign crh = ~CRH;  //complement 
assign obe = ~OBE;  //complement 
assign obf = ~OBF;  //complement 
assign obg = ~OBG;  //complement 
assign obd = ~OBD;  //complement 
assign NKB =  NAQ  ; 
assign nkb = ~NKB;  //complement 
assign PAP =  PAO & PAK  ; 
assign pap = ~PAP;  //complement 
assign RBA =  NBA & naq  ; 
assign rba = ~RBA;  //complement 
assign RBB =  NBB & nfb  ; 
assign rbb = ~RBB;  //complement 
assign RBC =  NBC & nfc  ; 
assign rbc = ~RBC;  //complement 
assign dvg = ~DVG;  //complement 
assign drc = ~DRC;  //complement 
assign DRD = ~drd;  //complement 
assign RBD =  NBD & nfd  ; 
assign rbd = ~RBD;  //complement 
assign RBE =  NBE & nfe  ; 
assign rbe = ~RBE;  //complement 
assign RBF =  NBF & nff  ; 
assign rbf = ~RBF;  //complement 
assign nah = ~NAH;  //complement 
assign mzd = ~MZD;  //complement 
assign MZE = ~mze;  //complement 
assign dsa = ~DSA;  //complement 
assign DSB = ~dsb;  //complement 
assign EXR =  QVD & qvf & qvg  |  qvd & QVF & qvg  |  qvd & qvf & QVG  |  QVD & QVF & QVG  ; 
assign exr = ~EXR; //complement 
assign exs =  QVD & qvf & qvg  |  qvd & QVF & qvg  |  qvd & qvf & QVG  |  qvd & qvf & qvg  ; 
assign EXS = ~exs;  //complement 
assign neh = ~NEH;  //complement 
assign RBG =  NBG & nfg  ; 
assign rbg = ~RBG;  //complement 
assign RBH =  NBH & nfh  ; 
assign rbh = ~RBH;  //complement 
assign RBI =  NBI & nfi  ; 
assign rbi = ~RBI;  //complement 
assign dsc = ~DSC;  //complement 
assign DSD = ~dsd;  //complement 
assign mkb = ~MKB;  //complement 
assign nei = ~NEI;  //complement 
assign nek = ~NEK;  //complement 
assign dse = ~DSE;  //complement 
assign DSF = ~dsf;  //complement 
assign fzi = ~FZI;  //complement 
assign FZJ = ~fzj;  //complement 
assign fze = ~FZE;  //complement 
assign FZF = ~fzf;  //complement 
assign EXT =  QXP & qxr & qxt  |  qxp & QXR & qxt  |  qxp & qxr & QXT  |  QXP & QXR & QXT  ; 
assign ext = ~EXT; //complement 
assign exu =  QXP & qxr & qxt  |  qxp & QXR & qxt  |  qxp & qxr & QXT  |  qxp & qxr & qxt  ; 
assign EXU = ~exu;  //complement 
assign dta = ~DTA;  //complement 
assign DTB = ~dtb;  //complement 
assign fzg = ~FZG;  //complement 
assign fzh = ~FZH;  //complement 
assign EXF =  DWF  ; 
assign exf = ~EXF;  //complement 
assign ECA =  DHA  ; 
assign eca = ~ECA;  //complement 
assign LFC =  ZZO  ; 
assign lfc = ~LFC;  //complement 
assign EWE =  DWG & dwh & dvf  |  dwg & DWH & dvf  |  dwg & dwh & DVF  |  DWG & DWH & DVF  ; 
assign ewe = ~EWE; //complement 
assign ewf =  DWG & dwh & dvf  |  dwg & DWH & dvf  |  dwg & dwh & DVF  |  dwg & dwh & dvf  ; 
assign EWF = ~ewf;  //complement 
assign dtc = ~DTC;  //complement 
assign DTD = ~dtd;  //complement 
assign nub =  nbi  ; 
assign NUB = ~nub;  //complement 
assign nuc =  nfj & nbi  |  nbj  ; 
assign NUC = ~nuc;  //complement 
assign EXI =  QXQ & qxs & qxd  |  qxq & QXS & qxd  |  qxq & qxs & QXD  |  QXQ & QXS & QXD  ; 
assign exi = ~EXI; //complement 
assign exj =  QXQ & qxs & qxd  |  qxq & QXS & qxd  |  qxq & qxs & QXD  |  qxq & qxs & qxd  ; 
assign EXJ = ~exj;  //complement 
assign EXN =  QXV & qxx & qxl  |  qxv & QXX & qxl  |  qxv & qxx & QXL  |  QXV & QXX & QXL  ; 
assign exn = ~EXN; //complement 
assign exo =  QXV & qxx & qxl  |  qxv & QXX & qxl  |  qxv & qxx & QXL  |  qxv & qxx & qxl  ; 
assign EXO = ~exo;  //complement 
assign EXP =  QXZ & qvb & qxn  |  qxz & QVB & qxn  |  qxz & qvb & QXN  |  QXZ & QVB & QXN  ; 
assign exp = ~EXP; //complement 
assign exq =  QXZ & qvb & qxn  |  qxz & QVB & qxn  |  qxz & qvb & QXN  |  qxz & qvb & qxn  ; 
assign EXQ = ~exq;  //complement 
assign bbd = ~BBD;  //complement 
assign bbe = ~BBE;  //complement 
assign bbf = ~BBF;  //complement 
assign bba = ~BBA;  //complement 
assign bbb = ~BBB;  //complement 
assign bbc = ~BBC;  //complement 
assign dqc = ~DQC;  //complement 
assign DQD = ~dqd;  //complement 
assign dra = ~DRA;  //complement 
assign DRB = ~drb;  //complement 
assign duc = ~DUC;  //complement 
assign DUD = ~dud;  //complement 
assign GZM =  FZR & fzt & fzn  |  fzr & FZT & fzn  |  fzr & fzt & FZN  |  FZR & FZT & FZN  ; 
assign gzm = ~GZM; //complement 
assign gzn =  FZR & fzt & fzn  |  fzr & FZT & fzn  |  fzr & fzt & FZN  |  fzr & fzt & fzn  ; 
assign GZN = ~gzn;  //complement 
assign EZS =  QYJ & qyl & qyb  |  qyj & QYL & qyb  |  qyj & qyl & QYB  |  QYJ & QYL & QYB  ; 
assign ezs = ~EZS; //complement 
assign ezt =  QYJ & qyl & qyb  |  qyj & QYL & qyb  |  qyj & qyl & QYB  |  qyj & qyl & qyb  ; 
assign EZT = ~ezt;  //complement 
assign EZU =  QYN & qyp & qyd  |  qyn & QYP & qyd  |  qyn & qyp & QYD  |  QYN & QYP & QYD  ; 
assign ezu = ~EZU; //complement 
assign ezv =  QYN & qyp & qyd  |  qyn & QYP & qyd  |  qyn & qyp & QYD  |  qyn & qyp & qyd  ; 
assign EZV = ~ezv;  //complement 
assign due = ~DUE;  //complement 
assign DUF = ~duf;  //complement 
assign fea = ~FEA;  //complement 
assign nel = ~NEL;  //complement 
assign EZW =  QYR & qyh & qyf  |  qyr & QYH & qyf  |  qyr & qyh & QYF  |  QYR & QYH & QYF  ; 
assign ezw = ~EZW; //complement 
assign ezx =  QYR & qyh & qyf  |  qyr & QYH & qyf  |  qyr & qyh & QYF  |  qyr & qyh & qyf  ; 
assign EZX = ~ezx;  //complement 
assign qys = ~QYS;  //complement 
assign dva = ~DVA;  //complement 
assign DVB = ~dvb;  //complement 
assign frc = ~FRC;  //complement 
assign nem = ~NEM;  //complement 
assign hna = ~HNA;  //complement 
assign hnb = ~HNB;  //complement 
assign hoa = ~HOA;  //complement 
assign fwc = ~FWC;  //complement 
assign EJA =  DJA & did & djc  |  dja & DID & djc  |  dja & did & DJC  |  DJA & DID & DJC  ; 
assign eja = ~EJA; //complement 
assign ejb =  DJA & did & djc  |  dja & DID & djc  |  dja & did & DJC  |  dja & did & djc  ; 
assign EJB = ~ejb;  //complement 
assign dvc = ~DVC;  //complement 
assign DVD = ~dvd;  //complement 
assign GZZ =  FYH & fyn  |  fyh & FYN  ; 
assign gzz = ~GZZ;  //complement 
assign EKA =  DKA & djb & dkc  |  dka & DJB & dkc  |  dka & djb & DKC  |  DKA & DJB & DKC  ; 
assign eka = ~EKA; //complement 
assign ekb =  DKA & djb & dkc  |  dka & DJB & dkc  |  dka & djb & DKC  |  dka & djb & dkc  ; 
assign EKB = ~ekb;  //complement 
assign ELA =  DLA & dkb & dlc  |  dla & DKB & dlc  |  dla & dkb & DLC  |  DLA & DKB & DLC  ; 
assign ela = ~ELA; //complement 
assign elb =  DLA & dkb & dlc  |  dla & DKB & dlc  |  dla & dkb & DLC  |  dla & dkb & dlc  ; 
assign ELB = ~elb;  //complement 
assign dve = ~DVE;  //complement 
assign DVF = ~dvf;  //complement 
assign kxa = ~KXA;  //complement 
assign KXB = ~kxb;  //complement 
assign EMA =  DMA & dlb & dmc  |  dma & DLB & dmc  |  dma & dlb & DMC  |  DMA & DLB & DMC  ; 
assign ema = ~EMA; //complement 
assign emb =  DMA & dlb & dmc  |  dma & DLB & dmc  |  dma & dlb & DMC  |  dma & dlb & dmc  ; 
assign EMB = ~emb;  //complement 
assign ENA =  DNA & dmb & dnc  |  dna & DMB & dnc  |  dna & dmb & DNC  |  DNA & DMB & DNC  ; 
assign ena = ~ENA; //complement 
assign enb =  DNA & dmb & dnc  |  dna & DMB & dnc  |  dna & dmb & DNC  |  dna & dmb & dnc  ; 
assign ENB = ~enb;  //complement 
assign dwa = ~DWA;  //complement 
assign DWB = ~dwb;  //complement 
assign fzm = ~FZM;  //complement 
assign FZN = ~fzn;  //complement 
assign EOA =  DOA & dnb & doc  |  doa & DNB & doc  |  doa & dnb & DOC  |  DOA & DNB & DOC  ; 
assign eoa = ~EOA; //complement 
assign eob =  DOA & dnb & doc  |  doa & DNB & doc  |  doa & dnb & DOC  |  doa & dnb & doc  ; 
assign EOB = ~eob;  //complement 
assign EPA =  DPA & dob & dpc  |  dpa & DOB & dpc  |  dpa & dob & DPC  |  DPA & DOB & DPC  ; 
assign epa = ~EPA; //complement 
assign epb =  DPA & dob & dpc  |  dpa & DOB & dpc  |  dpa & dob & DPC  |  dpa & dob & dpc  ; 
assign EPB = ~epb;  //complement 
assign dte = ~DTE;  //complement 
assign DTF = ~dtf;  //complement 
assign hzg = ~HZG;  //complement 
assign HZH = ~hzh;  //complement 
assign GZG =  FZI & fzk & fzf  |  fzi & FZK & fzf  |  fzi & fzk & FZF  |  FZI & FZK & FZF  ; 
assign gzg = ~GZG; //complement 
assign gzh =  FZI & fzk & fzf  |  fzi & FZK & fzf  |  fzi & fzk & FZF  |  fzi & fzk & fzf  ; 
assign GZH = ~gzh;  //complement 
assign GZI =  FZM & fzo & fzj  |  fzm & FZO & fzj  |  fzm & fzo & FZJ  |  FZM & FZO & FZJ  ; 
assign gzi = ~GZI; //complement 
assign gzj =  FZM & fzo & fzj  |  fzm & FZO & fzj  |  fzm & fzo & FZJ  |  fzm & fzo & fzj  ; 
assign GZJ = ~gzj;  //complement 
assign dua = ~DUA;  //complement 
assign DUB = ~dub;  //complement 
assign hxc = ~HXC;  //complement 
assign foc = ~FOC;  //complement 
assign fcb = ~FCB;  //complement 
assign GZV =  FYI  ; 
assign gzv = ~GZV;  //complement 
assign GZW =  FZZ  ; 
assign gzw = ~GZW;  //complement 
assign EIA =  DIC & dib & die  |  dic & DIB & die  |  dic & dib & DIE  |  DIC & DIB & DIE  ; 
assign eia = ~EIA; //complement 
assign eib =  DIC & dib & die  |  dic & DIB & die  |  dic & dib & DIE  |  dic & dib & die  ; 
assign EIB = ~eib;  //complement 
assign CBI = BAB & ADB ; 
assign cbi = ~CBI ; //complement 
assign CBJ = BAB & ADD ; 
assign cbj = ~CBJ ;  //complement 
assign CBK = BAB & ADF ; 
assign cbk = ~CBK ;  //complement 
assign CBL = BAB & ADH; 
assign cbl = ~CBL; 
assign CSA =  BBC & ACA  ; 
assign csa = ~CSA;  //complement 
assign CSB =  BBC & ACC  ; 
assign csb = ~CSB;  //complement 
assign CSC =  BBC & ACE  ; 
assign csc = ~CSC;  //complement 
assign frd = ~FRD;  //complement 
assign mbb = ~MBB;  //complement 
assign obh = ~OBH;  //complement 
assign CBM = BAB & ADJ ; 
assign cbm = ~CBM ; //complement 
assign CBN = BAB & ADL ; 
assign cbn = ~CBN ;  //complement 
assign CBO = BAB & ADN ; 
assign cbo = ~CBO ;  //complement 
assign CBP = BAB & ADO; 
assign cbp = ~CBP; 
assign CSD =  BBC & ACG  ; 
assign csd = ~CSD;  //complement 
assign CSE =  BBC & ACI  ; 
assign cse = ~CSE;  //complement 
assign CSF =  BBC & ACK  ; 
assign csf = ~CSF;  //complement 
assign LYA =  HYA & hxb & kza  |  hya & HXB & kza  |  hya & hxb & KZA  |  HYA & HXB & KZA  ; 
assign lya = ~LYA; //complement 
assign lyb =  HYA & hxb & kza  |  hya & HXB & kza  |  hya & hxb & KZA  |  hya & hxb & kza  ; 
assign LYB = ~lyb;  //complement 
assign obi = ~OBI;  //complement 
assign obj = ~OBJ;  //complement 
assign obk = ~OBK;  //complement 
assign fyq = ~FYQ;  //complement 
assign FYR = ~fyr;  //complement 
assign CSG =  BBC & ACM  ; 
assign csg = ~CSG;  //complement 
assign CTA =  BBD & ACB  ; 
assign cta = ~CTA;  //complement 
assign CTB =  BBD & ACD  ; 
assign ctb = ~CTB;  //complement 
assign mja = ~MJA;  //complement 
assign MJB = ~mjb;  //complement 
assign obl = ~OBL;  //complement 
assign obm = ~OBM;  //complement 
assign obn = ~OBN;  //complement 
assign CCA = BAC & ACA ; 
assign cca = ~CCA ; //complement 
assign CCB = BAC & ACC ; 
assign ccb = ~CCB ;  //complement 
assign CCC = BAC & ACE ; 
assign ccc = ~CCC ;  //complement 
assign CCD = BAC & ACG; 
assign ccd = ~CCD; 
assign CTC =  BBD & ACF  ; 
assign ctc = ~CTC;  //complement 
assign CTD =  BBD & ACH  ; 
assign ctd = ~CTD;  //complement 
assign CTE =  BBD & ACJ  ; 
assign cte = ~CTE;  //complement 
assign fqc = ~FQC;  //complement 
assign hzo = ~HZO;  //complement 
assign fwd = ~FWD;  //complement 
assign obo = ~OBO;  //complement 
assign obp = ~OBP;  //complement 
assign CCE = BAC & ACI ; 
assign cce = ~CCE ; //complement 
assign CCF = BAC & ACK ; 
assign ccf = ~CCF ;  //complement 
assign CCG = BAC & ACM ; 
assign ccg = ~CCG ;  //complement 
assign CCH = BAC & ACO; 
assign cch = ~CCH; 
assign CTF =  BBD & ACL  ; 
assign ctf = ~CTF;  //complement 
assign CTG =  BBD & ACN  ; 
assign ctg = ~CTG;  //complement 
assign CUA =  BBE & ACA  ; 
assign cua = ~CUA;  //complement 
assign mma = ~MMA;  //complement 
assign ENC =  DMD  ; 
assign enc = ~ENC;  //complement 
assign CCI = BAC & ADA ; 
assign cci = ~CCI ; //complement 
assign CCJ = BAC & ADC ; 
assign ccj = ~CCJ ;  //complement 
assign CUB =  BBE & ACC  ; 
assign cub = ~CUB;  //complement 
assign CUC =  BBE & ACE  ; 
assign cuc = ~CUC;  //complement 
assign CUD =  BBE & ACG  ; 
assign cud = ~CUD;  //complement 
assign GZQ =  FZW & fzy & fzs  |  fzw & FZY & fzs  |  fzw & fzy & FZS  |  FZW & FZY & FZS  ; 
assign gzq = ~GZQ; //complement 
assign gzr =  FZW & fzy & fzs  |  fzw & FZY & fzs  |  fzw & fzy & FZS  |  fzw & fzy & fzs  ; 
assign GZR = ~gzr;  //complement 
assign nfb = ~NFB;  //complement 
assign CCK = BAC & ADE ; 
assign cck = ~CCK ; //complement 
assign CCL = BAC & ADG ; 
assign ccl = ~CCL ;  //complement 
assign CCM = BAC & ADI ; 
assign ccm = ~CCM ;  //complement 
assign CCN = BAC & ADK; 
assign ccn = ~CCN; 
assign CUE =  BBE & ACI  ; 
assign cue = ~CUE;  //complement 
assign CUF =  BBE & ACK  ; 
assign cuf = ~CUF;  //complement 
assign fdb = ~FDB;  //complement 
assign fzv = ~FZV;  //complement 
assign fyi = ~FYI;  //complement 
assign kba = ~KBA;  //complement 
assign kca = ~KCA;  //complement 
assign CCO =  ADM & BAC  ; 
assign cco = ~CCO;  //complement 
assign CVA = BBF & ACB ; 
assign cva = ~CVA ; //complement 
assign CVB = BBF & ACD ; 
assign cvb = ~CVB ;  //complement 
assign CVC = BBF & ACF ; 
assign cvc = ~CVC ;  //complement 
assign CVD = BBF & ACH; 
assign cvd = ~CVD; 
assign kda = ~KDA;  //complement 
assign nen = ~NEN;  //complement 
assign aaq = ~AAQ;  //complement 
assign foa = ~FOA;  //complement 
assign FOB = ~fob;  //complement 
assign fpa = ~FPA;  //complement 
assign FPB = ~fpb;  //complement 
assign dwc = ~DWC;  //complement 
assign DWD = ~dwd;  //complement 
assign RBN =  NBN & nfn  ; 
assign rbn = ~RBN;  //complement 
assign RBO =  NBO & nfo  ; 
assign rbo = ~RBO;  //complement 
assign RBP =  NBP & nfp  ; 
assign rbp = ~RBP;  //complement 
assign fqa = ~FQA;  //complement 
assign FQB = ~fqb;  //complement 
assign fra = ~FRA;  //complement 
assign FRB = ~frb;  //complement 
assign dwe = ~DWE;  //complement 
assign DWF = ~dwf;  //complement 
assign fyj = ~FYJ;  //complement 
assign FYK = ~fyk;  //complement 
assign fsa = ~FSA;  //complement 
assign FSB = ~fsb;  //complement 
assign fta = ~FTA;  //complement 
assign FTB = ~ftb;  //complement 
assign dxa = ~DXA;  //complement 
assign DXB = ~dxb;  //complement 
assign qzi = ~QZI;  //complement 
assign fua = ~FUA;  //complement 
assign FUB = ~fub;  //complement 
assign fva = ~FVA;  //complement 
assign FVB = ~fvb;  //complement 
assign dxc = ~DXC;  //complement 
assign DXD = ~dxd;  //complement 
assign mka = ~MKA;  //complement 
assign fwa = ~FWA;  //complement 
assign FWB = ~fwb;  //complement 
assign hzy = ~HZY;  //complement 
assign HZZ = ~hzz;  //complement 
assign dxe = ~DXE;  //complement 
assign DXF = ~dxf;  //complement 
assign hra = ~HRA;  //complement 
assign HRB = ~hrb;  //complement 
assign fxa = ~FXA;  //complement 
assign FXB = ~fxb;  //complement 
assign fxc = ~FXC;  //complement 
assign FXD = ~fxd;  //complement 
assign hzq = ~HZQ;  //complement 
assign HZR = ~hzr;  //complement 
assign RBK =  NBK & nfk  ; 
assign rbk = ~RBK;  //complement 
assign RBL =  NBL & nfl  ; 
assign rbl = ~RBL;  //complement 
assign RBM =  NBM & nfm  ; 
assign rbm = ~RBM;  //complement 
assign fia = ~FIA;  //complement 
assign FIB = ~fib;  //complement 
assign kaa = ~KAA;  //complement 
assign fja = ~FJA;  //complement 
assign FJB = ~fjb;  //complement 
assign hzw = ~HZW;  //complement 
assign HZX = ~hzx;  //complement 
assign kzm = ~KZM;  //complement 
assign KZN = ~kzn;  //complement 
assign fma = ~FMA;  //complement 
assign fmb = ~FMB;  //complement 
assign kzt = ~KZT;  //complement 
assign kzy = ~KZY;  //complement 
assign fna = ~FNA;  //complement 
assign FNB = ~fnb;  //complement 
assign dye = ~DYE;  //complement 
assign DYF = ~dyf;  //complement 
assign OIA = ~oia;  //complement 
assign OKA = ~oka;  //complement 
assign OMA = ~oma;  //complement 
assign OOA = ~ooa;  //complement 
assign ERC =  DRF & dqd & dre  |  drf & DQD & dre  |  drf & dqd & DRE  |  DRF & DQD & DRE  ; 
assign erc = ~ERC; //complement 
assign erd =  DRF & dqd & dre  |  drf & DQD & dre  |  drf & dqd & DRE  |  drf & dqd & dre  ; 
assign ERD = ~erd;  //complement 
assign ESA =  DSA & drb & dsc  |  dsa & DRB & dsc  |  dsa & drb & DSC  |  DSA & DRB & DSC  ; 
assign esa = ~ESA; //complement 
assign esb =  DSA & drb & dsc  |  dsa & DRB & dsc  |  dsa & drb & DSC  |  dsa & drb & dsc  ; 
assign ESB = ~esb;  //complement 
assign dyg = ~DYG;  //complement 
assign DYH = ~dyh;  //complement 
assign nep = ~NEP;  //complement 
assign ESC =  DSE  ; 
assign esc = ~ESC;  //complement 
assign ESD =  DRD  ; 
assign esd = ~ESD;  //complement 
assign EYY =  QXI  ; 
assign eyy = ~EYY;  //complement 
assign ETA =  DTA & dsb & dtc  |  dta & DSB & dtc  |  dta & dsb & DTC  |  DTA & DSB & DTC  ; 
assign eta = ~ETA; //complement 
assign etb =  DTA & dsb & dtc  |  dta & DSB & dtc  |  dta & dsb & DTC  |  dta & dsb & dtc  ; 
assign ETB = ~etb;  //complement 
assign dza = ~DZA;  //complement 
assign DZB = ~dzb;  //complement 
assign ntd =  nff & nfg & nbe  |  nfg & nbf  |  nbg  ; 
assign NTD = ~ntd; //complement 
assign ETC =  DTE & dsf & dsd  |  dte & DSF & dsd  |  dte & dsf & DSD  |  DTE & DSF & DSD  ; 
assign etc = ~ETC; //complement 
assign etd =  DTE & dsf & dsd  |  dte & DSF & dsd  |  dte & dsf & DSD  |  dte & dsf & dsd  ; 
assign ETD = ~etd;  //complement 
assign EUA =  DUA & dtb & duc  |  dua & DTB & duc  |  dua & dtb & DUC  |  DUA & DTB & DUC  ; 
assign eua = ~EUA; //complement 
assign eub =  DUA & dtb & duc  |  dua & DTB & duc  |  dua & dtb & DUC  |  dua & dtb & duc  ; 
assign EUB = ~eub;  //complement 
assign dzc = ~DZC;  //complement 
assign DZD = ~dzd;  //complement 
assign GYC =  FXD  ; 
assign gyc = ~GYC;  //complement 
assign EUC =  DUE & dtf & dug  |  due & DTF & dug  |  due & dtf & DUG  |  DUE & DTF & DUG  ; 
assign euc = ~EUC; //complement 
assign eud =  DUE & dtf & dug  |  due & DTF & dug  |  due & dtf & DUG  |  due & dtf & dug  ; 
assign EUD = ~eud;  //complement 
assign EVA =  DVA & dub & dvc  |  dva & DUB & dvc  |  dva & dub & DVC  |  DVA & DUB & DVC  ; 
assign eva = ~EVA; //complement 
assign evb =  DVA & dub & dvc  |  dva & DUB & dvc  |  dva & dub & DVC  |  dva & dub & dvc  ; 
assign EVB = ~evb;  //complement 
assign dze = ~DZE;  //complement 
assign DZF = ~dzf;  //complement 
assign nrc =  nen & nam  |  nan  ; 
assign NRC = ~nrc; //complement 
assign EVC =  DVE & dvg & duf  |  dve & DVG & duf  |  dve & dvg & DUF  |  DVE & DVG & DUF  ; 
assign evc = ~EVC; //complement 
assign evd =  DVE & dvg & duf  |  dve & DVG & duf  |  dve & dvg & DUF  |  dve & dvg & duf  ; 
assign EVD = ~evd;  //complement 
assign EWA =  DWA & dvb & dwb  |  dwa & DVB & dwb  |  dwa & dvb & DWB  |  DWA & DVB & DWB  ; 
assign ewa = ~EWA; //complement 
assign ewb =  DWA & dvb & dwb  |  dwa & DVB & dwb  |  dwa & dvb & DWB  |  dwa & dvb & dwb  ; 
assign EWB = ~ewb;  //complement 
assign dzg = ~DZG;  //complement 
assign DZH = ~dzh;  //complement 
assign mla = ~MLA;  //complement 
assign EWC =  DWC & dwe & dvd  |  dwc & DWE & dvd  |  dwc & dwe & DVD  |  DWC & DWE & DVD  ; 
assign ewc = ~EWC; //complement 
assign ewd =  DWC & dwe & dvd  |  dwc & DWE & dvd  |  dwc & dwe & DVD  |  dwc & dwe & dvd  ; 
assign EWD = ~ewd;  //complement 
assign EXA =  DXA & dwb & dxc  |  dxa & DWB & dxc  |  dxa & dwb & DXC  |  DXA & DWB & DXC  ; 
assign exa = ~EXA; //complement 
assign exb =  DXA & dwb & dxc  |  dxa & DWB & dxc  |  dxa & dwb & DXC  |  dxa & dwb & dxc  ; 
assign EXB = ~exb;  //complement 
assign dya = ~DYA;  //complement 
assign DYB = ~dyb;  //complement 
assign RBJ =  NBJ & nfj  ; 
assign rbj = ~RBJ;  //complement 
assign EPC =  DPE  ; 
assign epc = ~EPC;  //complement 
assign EPD =  DOD  ; 
assign epd = ~EPD;  //complement 
assign EUE =  DTD  ; 
assign eue = ~EUE;  //complement 
assign EQA =  DQA & dpb & dqc  |  dqa & DPB & dqc  |  dqa & dpb & DQC  |  DQA & DPB & DQC  ; 
assign eqa = ~EQA; //complement 
assign eqb =  DQA & dpb & dqc  |  dqa & DPB & dqc  |  dqa & dpb & DQC  |  dqa & dpb & dqc  ; 
assign EQB = ~eqb;  //complement 
assign dyc = ~DYC;  //complement 
assign DYD = ~dyd;  //complement 
assign OIH = ~oih;  //complement 
assign OKH = ~okh;  //complement 
assign OMH = ~omh;  //complement 
assign OOH = ~ooh;  //complement 
assign EQC =  DQF & dqe & dpd  |  dqf & DQE & dpd  |  dqf & dqe & DPD  |  DQF & DQE & DPD  ; 
assign eqc = ~EQC; //complement 
assign eqd =  DQF & dqe & dpd  |  dqf & DQE & dpd  |  dqf & dqe & DPD  |  dqf & dqe & dpd  ; 
assign EQD = ~eqd;  //complement 
assign ERA =  DRA & dqb & drc  |  dra & DQB & drc  |  dra & dqb & DRC  |  DRA & DQB & DRC  ; 
assign era = ~ERA; //complement 
assign erb =  DRA & dqb & drc  |  dra & DQB & drc  |  dra & dqb & DRC  |  dra & dqb & drc  ; 
assign ERB = ~erb;  //complement 
assign CDA = BAD & ACB ; 
assign cda = ~CDA ; //complement 
assign CDB = BAD & ACD ; 
assign cdb = ~CDB ;  //complement 
assign CDC = BAD & ACF ; 
assign cdc = ~CDC ;  //complement 
assign CDD = BAD & ACH; 
assign cdd = ~CDD; 
assign CVE =  ACJ & BBF  ; 
assign cve = ~CVE;  //complement 
assign CVF =  ACL & BBF  ; 
assign cvf = ~CVF;  //complement 
assign EVF =  DUD  ; 
assign evf = ~EVF;  //complement 
assign kea = ~KEA;  //complement 
assign hfa = ~HFA;  //complement 
assign hfb = ~HFB;  //complement 
assign moa = ~MOA;  //complement 
assign MOB = ~mob;  //complement 
assign CDE = BAD & ACJ ; 
assign cde = ~CDE ; //complement 
assign CDF = BAD & ACL ; 
assign cdf = ~CDF ;  //complement 
assign CDG = BAD & ACN ; 
assign cdg = ~CDG ;  //complement 
assign CDH = BAD & ACP; 
assign cdh = ~CDH; 
assign CWA = BBG & ACA ; 
assign cwa = ~CWA ; //complement 
assign CWB = BBG & ACC ; 
assign cwb = ~CWB ;  //complement 
assign CWC = BBG & ACE ; 
assign cwc = ~CWC ;  //complement 
assign CWD = BBG & ACG; 
assign cwd = ~CWD; 
assign kfa = ~KFA;  //complement 
assign kga = ~KGA;  //complement 
assign fzc = ~FZC;  //complement 
assign FZD = ~fzd;  //complement 
assign CDI =  ADB & BAD  ; 
assign cdi = ~CDI;  //complement 
assign CDJ =  ADD & BAD  ; 
assign cdj = ~CDJ;  //complement 
assign nqb =  nai  ; 
assign NQB = ~nqb;  //complement 
assign CWE =  ACI & BBG  ; 
assign cwe = ~CWE;  //complement 
assign CXA =  BBH & ACB  ; 
assign cxa = ~CXA;  //complement 
assign CXB =  BBH & ACD  ; 
assign cxb = ~CXB;  //complement 
assign kia = ~KIA;  //complement 
assign fxe = ~FXE;  //complement 
assign EYE =  DXF  ; 
assign eye = ~EYE;  //complement 
assign CDK =  ADF & BAD  ; 
assign cdk = ~CDK;  //complement 
assign CDL =  ADH & BAD  ; 
assign cdl = ~CDL;  //complement 
assign CDM =  ADJ & BAD  ; 
assign cdm = ~CDM;  //complement 
assign CXC =  BBH & ACF  ; 
assign cxc = ~CXC;  //complement 
assign CXD =  BBH & ACH  ; 
assign cxd = ~CXD;  //complement 
assign CXE =  BBH & ACJ  ; 
assign cxe = ~CXE;  //complement 
assign kja = ~KJA;  //complement 
assign nfc = ~NFC;  //complement 
assign CDN =  ADL & BAD  ; 
assign cdn = ~CDN;  //complement 
assign CDO =  ADN & BAD  ; 
assign cdo = ~CDO;  //complement 
assign nrb =  nam  ; 
assign NRB = ~nrb;  //complement 
assign CYA =  BBI & ACA  ; 
assign cya = ~CYA;  //complement 
assign CYB =  BBI & ACC  ; 
assign cyb = ~CYB;  //complement 
assign CYC =  BBI & ACE  ; 
assign cyc = ~CYC;  //complement 
assign kma = ~KMA;  //complement 
assign kha = ~KHA;  //complement 
assign KHB = ~khb;  //complement 
assign CEA = BAE & ACA ; 
assign cea = ~CEA ; //complement 
assign CEB = BAE & ACC ; 
assign ceb = ~CEB ;  //complement 
assign CEC = BAE & ACE ; 
assign cec = ~CEC ;  //complement 
assign CED = BAE & ACG; 
assign ced = ~CED; 
assign CYD =  BBI & ACG  ; 
assign cyd = ~CYD;  //complement 
assign CZA =  BBJ & ACB  ; 
assign cza = ~CZA;  //complement 
assign CZB =  BBJ & ACD  ; 
assign czb = ~CZB;  //complement 
assign kna = ~KNA;  //complement 
assign koa = ~KOA;  //complement 
assign naq = ~NAQ;  //complement 
assign CEE = BAE & ACI ; 
assign cee = ~CEE ; //complement 
assign CEF = BAE & ACK ; 
assign cef = ~CEF ;  //complement 
assign CEG = BAE & ACM ; 
assign ceg = ~CEG ;  //complement 
assign CEH = BAE & ACO; 
assign ceh = ~CEH; 
assign CZC =  BBJ & ACF  ; 
assign czc = ~CZC;  //complement 
assign CZD =  BBJ & ACH  ; 
assign czd = ~CZD;  //complement 
assign DAA =  BBK & ACA  ; 
assign daa = ~DAA;  //complement 
assign kpa = ~KPA;  //complement 
assign kpb = ~KPB;  //complement 
assign kqa = ~KQA;  //complement 
assign fsd = ~FSD;  //complement 
assign CEI =  ADA & BAE  ; 
assign cei = ~CEI;  //complement 
assign CEJ =  ADC & BAE  ; 
assign cej = ~CEJ;  //complement 
assign EVE =  DVG  ; 
assign eve = ~EVE;  //complement 
assign DAB =  BBK & ACC  ; 
assign dab = ~DAB;  //complement 
assign DAC =  BBK & ACE  ; 
assign dac = ~DAC;  //complement 
assign DBA =  BBL & ACB  ; 
assign dba = ~DBA;  //complement 
assign kqb = ~KQB;  //complement 
assign kra = ~KRA;  //complement 
assign ksa = ~KSA;  //complement 
assign ksb = ~KSB;  //complement 
assign mna = ~MNA;  //complement 
assign nfg = ~NFG;  //complement 
assign nfh = ~NFH;  //complement 
assign nfi = ~NFI;  //complement 
assign kzw = ~KZW;  //complement 
assign nfl = ~NFL;  //complement 
assign PAK = ~pak;  //complement 
assign OIB = ~oib;  //complement 
assign OKB = ~okb;  //complement 
assign OMB = ~omb;  //complement 
assign OOB = ~oob;  //complement 
assign GZE =  FZH & fzd  |  fzh & FZD  ; 
assign gze = ~GZE;  //complement 
assign EDB =  DHD  ; 
assign edb = ~EDB;  //complement 
assign EOC =  DOE  ; 
assign eoc = ~EOC;  //complement 
assign fzk = ~FZK;  //complement 
assign FZL = ~fzl;  //complement 
assign LZW =  KZW  ; 
assign lzw = ~LZW;  //complement 
assign LZT =  KZR  ; 
assign lzt = ~LZT;  //complement 
assign LZZ =  KZY  ; 
assign lzz = ~LZZ;  //complement 
assign mqb = ~MQB;  //complement 
assign GNA =  FNA  ; 
assign gna = ~GNA;  //complement 
assign fzo = ~FZO;  //complement 
assign FZP = ~fzp;  //complement 
assign dlc = ~DLC;  //complement 
assign dld = ~DLD;  //complement 
assign dqe = ~DQE;  //complement 
assign dre = ~DRE;  //complement 
assign JZY =  HZY & hyd & hzx  |  hzy & HYD & hzx  |  hzy & hyd & HZX  |  HZY & HYD & HZX  ; 
assign jzy = ~JZY; //complement 
assign jzz =  HZY & hyd & hzx  |  hzy & HYD & hzx  |  hzy & hyd & HZX  |  hzy & hyd & hzx  ; 
assign JZZ = ~jzz;  //complement 
assign dqf = ~DQF;  //complement 
assign drf = ~DRF;  //complement 
assign fzy = ~FZY;  //complement 
assign FZZ = ~fzz;  //complement 
assign msa = ~MSA;  //complement 
assign MSB = ~msb;  //complement 
assign fha = ~FHA;  //complement 
assign hzk = ~HZK;  //complement 
assign hzv = ~HZV;  //complement 
assign OII = ~oii;  //complement 
assign OKI = ~oki;  //complement 
assign OMI = ~omi;  //complement 
assign OOI = ~ooi;  //complement 
assign GRC =  FRC  ; 
assign grc = ~GRC;  //complement 
assign fya = ~FYA;  //complement 
assign FYB = ~fyb;  //complement 
assign nqc =  nej & nai  |  naj  ; 
assign NQC = ~nqc; //complement 
assign nqd =  nek & nej & nai  |  nek & naj  |  nak  ; 
assign NQD = ~nqd; //complement 
assign EXM =  QXJ & qxo  |  qxj & QXO  ; 
assign exm = ~EXM;  //complement 
assign nff = ~NFF;  //complement 
assign npd =  nef & neg & nae  |  neg & naf  |  nag  ; 
assign NPD = ~npd; //complement 
assign npc =  nef & nae  |  naf  ; 
assign NPC = ~npc; //complement 
assign LZQ =  KZQ  ; 
assign lzq = ~LZQ;  //complement 
assign EYL =  QYQ  ; 
assign eyl = ~EYL;  //complement 
assign GYE =  FYN & FYH  ; 
assign gye = ~GYE;  //complement 
assign GYH =  FYM  ; 
assign gyh = ~GYH;  //complement 
assign dzm = ~DZM;  //complement 
assign DZN = ~dzn;  //complement 
assign OIJ = ~oij;  //complement 
assign OKJ = ~okj;  //complement 
assign OMJ = ~omj;  //complement 
assign OOJ = ~ooj;  //complement 
assign EXC =  DXE & dxg & dwd  |  dxe & DXG & dwd  |  dxe & dxg & DWD  |  DXE & DXG & DWD  ; 
assign exc = ~EXC; //complement 
assign exd =  DXE & dxg & dwd  |  dxe & DXG & dwd  |  dxe & dxg & DWD  |  dxe & dxg & dwd  ; 
assign EXD = ~exd;  //complement 
assign EYA =  DYA & dxb & dyc  |  dya & DXB & dyc  |  dya & dxb & DYC  |  DYA & DXB & DYC  ; 
assign eya = ~EYA; //complement 
assign eyb =  DYA & dxb & dyc  |  dya & DXB & dyc  |  dya & dxb & DYC  |  dya & dxb & dyc  ; 
assign EYB = ~eyb;  //complement 
assign dzo = ~DZO;  //complement 
assign DZP = ~dzp;  //complement 
assign kzx = ~KZX;  //complement 
assign EYC =  DYE & dyg & dxd  |  dye & DYG & dxd  |  dye & dyg & DXD  |  DYE & DYG & DXD  ; 
assign eyc = ~EYC; //complement 
assign eyd =  DYE & dyg & dxd  |  dye & DYG & dxd  |  dye & dyg & DXD  |  dye & dyg & dxd  ; 
assign EYD = ~eyd;  //complement 
assign EYF =  QZA & qyk & qzc  |  qza & QYK & qzc  |  qza & qyk & QZC  |  QZA & QYK & QZC  ; 
assign eyf = ~EYF; //complement 
assign eyg =  QZA & qyk & qzc  |  qza & QYK & qzc  |  qza & qyk & QZC  |  qza & qyk & qzc  ; 
assign EYG = ~eyg;  //complement 
assign qya = ~QYA;  //complement 
assign QYB = ~qyb;  //complement 
assign hyd = ~HYD;  //complement 
assign GSA =  FSA & fsc & fsd  |  fsa & FSC & fsd  |  fsa & fsc & FSD  |  FSA & FSC & FSD  ; 
assign gsa = ~GSA; //complement 
assign gsb =  FSA & fsc & fsd  |  fsa & FSC & fsd  |  fsa & fsc & FSD  |  fsa & fsc & fsd  ; 
assign GSB = ~gsb;  //complement 
assign GTA =  FTA & ftc & fsb  |  fta & FTC & fsb  |  fta & ftc & FSB  |  FTA & FTC & FSB  ; 
assign gta = ~GTA; //complement 
assign gtb =  FTA & ftc & fsb  |  fta & FTC & fsb  |  fta & ftc & FSB  |  fta & ftc & fsb  ; 
assign GTB = ~gtb;  //complement 
assign qyc = ~QYC;  //complement 
assign QYD = ~qyd;  //complement 
assign OIC = ~oic;  //complement 
assign mta = ~MTA;  //complement 
assign MTB = ~mtb;  //complement 
assign OKC = ~okc;  //complement 
assign GUA =  FUA & fuc & ftb  |  fua & FUC & ftb  |  fua & fuc & FTB  |  FUA & FUC & FTB  ; 
assign gua = ~GUA; //complement 
assign gub =  FUA & fuc & ftb  |  fua & FUC & ftb  |  fua & fuc & FTB  |  fua & fuc & ftb  ; 
assign GUB = ~gub;  //complement 
assign GVA =  FVA & fvc & fub  |  fva & FVC & fub  |  fva & fvc & FUB  |  FVA & FVC & FUB  ; 
assign gva = ~GVA; //complement 
assign gvb =  FVA & fvc & fub  |  fva & FVC & fub  |  fva & fvc & FUB  |  fva & fvc & fub  ; 
assign GVB = ~gvb;  //complement 
assign qye = ~QYE;  //complement 
assign QYF = ~qyf;  //complement 
assign OMC = ~omc;  //complement 
assign qvf = ~QVF;  //complement 
assign GWA =  FWA & fwc & fvb  |  fwa & FWC & fvb  |  fwa & fwc & FVB  |  FWA & FWC & FVB  ; 
assign gwa = ~GWA; //complement 
assign gwb =  FWA & fwc & fvb  |  fwa & FWC & fvb  |  fwa & fwc & FVB  |  fwa & fwc & fvb  ; 
assign GWB = ~gwb;  //complement 
assign GXA =  FXA & fxc & fwb  |  fxa & FXC & fwb  |  fxa & fxc & FWB  |  FXA & FXC & FWB  ; 
assign gxa = ~GXA; //complement 
assign gxb =  FXA & fxc & fwb  |  fxa & FXC & fwb  |  fxa & fxc & FWB  |  fxa & fxc & fwb  ; 
assign GXB = ~gxb;  //complement 
assign qyg = ~QYG;  //complement 
assign QYH = ~qyh;  //complement 
assign OOC = ~ooc;  //complement 
assign mfa = ~MFA;  //complement 
assign mwa = ~MWA;  //complement 
assign MWB = ~mwb;  //complement 
assign mxa = ~MXA;  //complement 
assign MXB = ~mxb;  //complement 
assign dzi = ~DZI;  //complement 
assign DZJ = ~dzj;  //complement 
assign hta = ~HTA;  //complement 
assign GOA =  FOA & foc & fnb  |  foa & FOC & fnb  |  foa & foc & FNB  |  FOA & FOC & FNB  ; 
assign goa = ~GOA; //complement 
assign gob =  FOA & foc & fnb  |  foa & FOC & fnb  |  foa & foc & FNB  |  foa & foc & fnb  ; 
assign GOB = ~gob;  //complement 
assign GPA =  FPA & fpc & fob  |  fpa & FPC & fob  |  fpa & fpc & FOB  |  FPA & FPC & FOB  ; 
assign gpa = ~GPA; //complement 
assign gpb =  FPA & fpc & fob  |  fpa & FPC & fob  |  fpa & fpc & FOB  |  fpa & fpc & fob  ; 
assign GPB = ~gpb;  //complement 
assign dzk = ~DZK;  //complement 
assign DZL = ~dzl;  //complement 
assign mrb = ~MRB;  //complement 
assign GQA =  FQA & fqc & fpb  |  fqa & FQC & fpb  |  fqa & fqc & FPB  |  FQA & FQC & FPB  ; 
assign gqa = ~GQA; //complement 
assign gqb =  FQA & fqc & fpb  |  fqa & FQC & fpb  |  fqa & fqc & FPB  |  fqa & fqc & fpb  ; 
assign GQB = ~gqb;  //complement 
assign GRA =  FRA & fqb & frd  |  fra & FQB & frd  |  fra & fqb & FRD  |  FRA & FQB & FRD  ; 
assign gra = ~GRA; //complement 
assign grb =  FRA & fqb & frd  |  fra & FQB & frd  |  fra & fqb & FRD  |  fra & fqb & frd  ; 
assign GRB = ~grb;  //complement 
assign CEK =  ADE & BAE  ; 
assign cek = ~CEK;  //complement 
assign CEL =  ADG & BAE  ; 
assign cel = ~CEL;  //complement 
assign CEM =  ADI & BAE  ; 
assign cem = ~CEM;  //complement 
assign DBB =  BBL & ACD  ; 
assign dbb = ~DBB;  //complement 
assign DBC =  BBL & ACF  ; 
assign dbc = ~DBC;  //complement 
assign DCA =  BBM & ACA  ; 
assign dca = ~DCA;  //complement 
assign kua = ~KUA;  //complement 
assign GZT =  FYE & fyg & fzx  |  fye & FYG & fzx  |  fye & fyg & FZX  |  FYE & FYG & FZX  ; 
assign gzt = ~GZT; //complement 
assign gzu =  FYE & fyg & fzx  |  fye & FYG & fzx  |  fye & fyg & FZX  |  fye & fyg & fzx  ; 
assign GZU = ~gzu;  //complement 
assign CEN =  ADK & BAE  ; 
assign cen = ~CEN;  //complement 
assign GZS =  FZU  ; 
assign gzs = ~GZS;  //complement 
assign GZP =  FZP & FZV  ; 
assign gzp = ~GZP;  //complement 
assign DCB =  BBM & ACC  ; 
assign dcb = ~DCB;  //complement 
assign DDA =  BBN & ACB  ; 
assign dda = ~DDA;  //complement 
assign DDB =  BBN & ACD  ; 
assign ddb = ~DDB;  //complement 
assign kwa = ~KWA;  //complement 
assign OIK = ~oik;  //complement 
assign OKK = ~okk;  //complement 
assign OMK = ~omk;  //complement 
assign OOK = ~ook;  //complement 
assign CFA = BAF & ACB ; 
assign cfa = ~CFA ; //complement 
assign CFB = BAF & ACD ; 
assign cfb = ~CFB ;  //complement 
assign CFC = BAF & ACF ; 
assign cfc = ~CFC ;  //complement 
assign CFD = BAF & ACH; 
assign cfd = ~CFD; 
assign DEA =  BBO & ACA  ; 
assign dea = ~DEA;  //complement 
assign DFA =  BBP & ACB  ; 
assign dfa = ~DFA;  //complement 
assign pab = ~PAB;  //complement 
assign OIE = ~oie;  //complement 
assign OKE = ~oke;  //complement 
assign OME = ~ome;  //complement 
assign OOE = ~ooe;  //complement 
assign CFE = BAF & ACJ ; 
assign cfe = ~CFE ; //complement 
assign CFF = BAF & ACL ; 
assign cff = ~CFF ;  //complement 
assign CFG = BAF & ACN ; 
assign cfg = ~CFG ;  //complement 
assign CFH = BAF & ACP; 
assign cfh = ~CFH; 
assign EXK =  QXU & qxf & qxh  |  qxu & QXF & qxh  |  qxu & qxf & QXH  |  QXU & QXF & QXH  ; 
assign exk = ~EXK; //complement 
assign exl =  QXU & qxf & qxh  |  qxu & QXF & qxh  |  qxu & qxf & QXH  |  qxu & qxf & qxh  ; 
assign EXL = ~exl;  //complement 
assign nsb =  nba  ; 
assign NSB = ~nsb;  //complement 
assign nsc =  nfb & nba  |  nbb  ; 
assign NSC = ~nsc;  //complement 
assign nsd =  nfb & nfc & nba  |  nfc & nbb  |  nbc  ; 
assign NSD = ~nsd; //complement 
assign CFI =  ADB & BAF  ; 
assign cfi = ~CFI;  //complement 
assign CFJ =  ADD & BAF  ; 
assign cfj = ~CFJ;  //complement 
assign CFK =  ADF & BAF  ; 
assign cfk = ~CFK;  //complement 
assign GMA =  FMA & fmb & fjb  |  fma & FMB & fjb  |  fma & fmb & FJB  |  FMA & FMB & FJB  ; 
assign gma = ~GMA; //complement 
assign gmb =  FMA & fmb & fjb  |  fma & FMB & fjb  |  fma & fmb & FJB  |  fma & fmb & fjb  ; 
assign GMB = ~gmb;  //complement 
assign pad = ~PAD;  //complement 
assign pae = ~PAE;  //complement 
assign CFL =  ADH & BAF  ; 
assign cfl = ~CFL;  //complement 
assign CFM =  ADJ & BAF  ; 
assign cfm = ~CFM;  //complement 
assign CFN =  ADL & BAF  ; 
assign cfn = ~CFN;  //complement 
assign kzi = ~KZI;  //complement 
assign KZJ = ~kzj;  //complement 
assign ntb =  nbe  ; 
assign NTB = ~ntb;  //complement 
assign ntc =  nff & nbe  |  nbf  ; 
assign NTC = ~ntc;  //complement 
assign nxb =  nae  |  naf  |  nag  |  nah  ;
assign NXB = ~nxb;  //complement 
assign CGA = BAG & ACA ; 
assign cga = ~CGA ; //complement 
assign CGB = BAG & ACC ; 
assign cgb = ~CGB ;  //complement 
assign CGC = BAG & ACE ; 
assign cgc = ~CGC ;  //complement 
assign CGD = BAG & ACG; 
assign cgd = ~CGD; 
assign haa = ~HAA;  //complement 
assign hba = ~HBA;  //complement 
assign hca = ~HCA;  //complement 
assign hda = ~HDA;  //complement 
assign GSC =  FRB  ; 
assign gsc = ~GSC;  //complement 
assign EEA =  DHE  ; 
assign eea = ~EEA;  //complement 
assign hzc = ~HZC;  //complement 
assign HZD = ~hzd;  //complement 
assign CGE = BAG & ACI ; 
assign cge = ~CGE ; //complement 
assign CGF = BAG & ACK ; 
assign cgf = ~CGF ;  //complement 
assign CGG = BAG & ACM ; 
assign cgg = ~CGG ;  //complement 
assign CGH = BAG & ACO; 
assign cgh = ~CGH; 
assign pfb = ~PFB;  //complement 
assign pfc = ~PFC;  //complement 
assign pfd = ~PFD;  //complement 
assign pfa = ~PFA;  //complement 
assign mea = ~MEA;  //complement 
assign OID = ~oid;  //complement 
assign OKD = ~okd;  //complement 
assign OMD = ~omd;  //complement 
assign OOD = ~ood;  //complement 
assign qzj = ~QZJ;  //complement 
assign NNB =  NFM  ; 
assign nnb = ~NNB;  //complement 
assign OIF = ~oif;  //complement 
assign OKF = ~okf;  //complement 
assign OMF = ~omf;  //complement 
assign OOF = ~oof;  //complement 
assign fyc = ~FYC;  //complement 
assign pdf = ~PDF;  //complement 
assign pdg = ~PDG;  //complement 
assign pdh = ~PDH;  //complement 
assign fye = ~FYE;  //complement 
assign FYF = ~fyf;  //complement 
assign pdk = ~PDK;  //complement 
assign pdl = ~PDL;  //complement 
assign pdj = ~PDJ;  //complement 
assign pdn = ~PDN;  //complement 
assign fyg = ~FYG;  //complement 
assign FYH = ~fyh;  //complement 
assign pdp = ~PDP;  //complement 
assign pdo = ~PDO;  //complement 
assign fyl = ~FYL;  //complement 
assign FYM = ~fym;  //complement 
assign OIL = ~oil;  //complement 
assign OKL = ~okl;  //complement 
assign OML = ~oml;  //complement 
assign OOL = ~ool;  //complement 
assign fsc = ~FSC;  //complement 
assign peb = ~PEB;  //complement 
assign mfb = ~MFB;  //complement 
assign pec = ~PEC;  //complement 
assign hua = ~HUA;  //complement 
assign HUB = ~hub;  //complement 
assign ped = ~PED;  //complement 
assign mqa = ~MQA;  //complement 
assign pac = ~PAC;  //complement 
assign nxc =  nai  |  naj  |  nak  |  nal  ;
assign NXC = ~nxc;  //complement 
assign nxd =  nam  |  nan  |  nao  |  nap  ;
assign NXD = ~nxd;  //complement 
assign nxe =  nba  |  nbb  |  nbc  |  nbd  ;
assign NXE = ~nxe;  //complement 
assign nxf =  nbe  |  nbf  |  nbg  |  nbh  ;
assign NXF = ~nxf;  //complement 
assign NNC =  NFM & NBN  |  NFN  ; 
assign nnc = ~NNC;  //complement 
assign kta = ~KTA;  //complement 
assign kzq = ~KZQ;  //complement 
assign qyn = ~QYN;  //complement 
assign QYO = ~qyo;  //complement 
assign pej = ~PEJ;  //complement 
assign mlb = ~MLB;  //complement 
assign GYA =  FYA & fyc & fxb  |  fya & FYC & fxb  |  fya & fyc & FXB  |  FYA & FYC & FXB  ; 
assign gya = ~GYA; //complement 
assign gyb =  FYA & fyc & fxb  |  fya & FYC & fxb  |  fya & fyc & FXB  |  fya & fyc & fxb  ; 
assign GYB = ~gyb;  //complement 
assign qyp = ~QYP;  //complement 
assign QYQ = ~qyq;  //complement 
assign pek = ~PEK;  //complement 
assign mra = ~MRA;  //complement 
assign GYF =  FYO & fyq & fyk  |  fyo & FYQ & fyk  |  fyo & fyq & FYK  |  FYO & FYQ & FYK  ; 
assign gyf = ~GYF; //complement 
assign gyg =  FYO & fyq & fyk  |  fyo & FYQ & fyk  |  fyo & fyq & FYK  |  fyo & fyq & fyk  ; 
assign GYG = ~gyg;  //complement 
assign qza = ~QZA;  //complement 
assign QZB = ~qzb;  //complement 
assign pep = ~PEP;  //complement 
assign GYI =  FYS  ; 
assign gyi = ~GYI;  //complement 
assign GYL =  FYD  ; 
assign gyl = ~GYL;  //complement 
assign LFB =  KFA & HEA  ; 
assign lfb = ~LFB;  //complement 
assign LZC =  KZB  ; 
assign lzc = ~LZC;  //complement 
assign LDC =  KDB  ; 
assign ldc = ~LDC;  //complement 
assign npb =  nae  ; 
assign NPB = ~npb;  //complement 
assign qzc = ~QZC;  //complement 
assign QZD = ~qzd;  //complement 
assign pel = ~PEL;  //complement 
assign LBA =  HAA  ; 
assign lba = ~LBA;  //complement 
assign LBB =  KBA  ; 
assign lbb = ~LBB;  //complement 
assign nfe = ~NFE;  //complement 
assign qze = ~QZE;  //complement 
assign QZF = ~qzf;  //complement 
assign OIM = ~oim;  //complement 
assign OKM = ~okm;  //complement 
assign OMM = ~omm;  //complement 
assign OOM = ~oom;  //complement 
assign LCA =  HBA & kca & kcb  |  hba & KCA & kcb  |  hba & kca & KCB  |  HBA & KCA & KCB  ; 
assign lca = ~LCA; //complement 
assign lcb =  HBA & kca & kcb  |  hba & KCA & kcb  |  hba & kca & KCB  |  hba & kca & kcb  ; 
assign LCB = ~lcb;  //complement 
assign kzr = ~KZR;  //complement 
assign qzg = ~QZG;  //complement 
assign QZH = ~qzh;  //complement 
assign nfk = ~NFK;  //complement 
assign LDA =  KDA & hca & hcb  |  kda & HCA & hcb  |  kda & hca & HCB  |  KDA & HCA & HCB  ; 
assign lda = ~LDA; //complement 
assign ldb =  KDA & hca & hcb  |  kda & HCA & hcb  |  kda & hca & HCB  |  kda & hca & hcb  ; 
assign LDB = ~ldb;  //complement 
assign kva = ~KVA;  //complement 
assign qyj = ~QYJ;  //complement 
assign QYK = ~qyk;  //complement 
assign peg = ~PEG;  //complement 
assign LEA =  KEA & hda & hdb  |  kea & HDA & hdb  |  kea & hda & HDB  |  KEA & HDA & HDB  ; 
assign lea = ~LEA; //complement 
assign leb =  KEA & hda & hdb  |  kea & HDA & hdb  |  kea & hda & HDB  |  kea & hda & hdb  ; 
assign LEB = ~leb;  //complement 
assign mua = ~MUA;  //complement 
assign MUB = ~mub;  //complement 
assign qyl = ~QYL;  //complement 
assign QYM = ~qym;  //complement 
assign peh = ~PEH;  //complement 
assign LFA =  KFA & hea  |  kfa & HEA  ; 
assign lfa = ~LFA;  //complement 
assign LGA =  KGA & hfa & hfb  |  kga & HFA & hfb  |  kga & hfa & HFB  |  KGA & HFA & HFB  ; 
assign lga = ~LGA; //complement 
assign lgb =  KGA & hfa & hfb  |  kga & HFA & hfb  |  kga & hfa & HFB  |  kga & hfa & hfb  ; 
assign LGB = ~lgb;  //complement 
assign CGI =  ADA & BAG  ; 
assign cgi = ~CGI;  //complement 
assign EYH =  QZE & qzg & qym  |  qze & QZG & qym  |  qze & qzg & QYM  |  QZE & QZG & QYM  ; 
assign eyh = ~EYH; //complement 
assign eyi =  QZE & qzg & qym  |  qze & QZG & qym  |  qze & qzg & QYM  |  qze & qzg & qym  ; 
assign EYI = ~eyi;  //complement 
assign naa = ~NAA;  //complement 
assign nac = ~NAC;  //complement 
assign qvg = ~QVG;  //complement 
assign OHF = ~ohf;  //complement 
assign CGJ =  ADC & BAG  ; 
assign cgj = ~CGJ;  //complement 
assign CGK =  ADE & BAG  ; 
assign cgk = ~CGK;  //complement 
assign CGL =  ADG & BAG  ; 
assign cgl = ~CGL;  //complement 
assign oja = ~OJA;  //complement 
assign ola = ~OLA;  //complement 
assign ona = ~ONA;  //complement 
assign opa = ~OPA;  //complement 
assign nad = ~NAD;  //complement 
assign nae = ~NAE;  //complement 
assign CGM =  ADI & BAG  ; 
assign cgm = ~CGM;  //complement 
assign ERE =  ZZO  ; 
assign ere = ~ERE;  //complement 
assign fuc = ~FUC;  //complement 
assign ojb = ~OJB;  //complement 
assign olb = ~OLB;  //complement 
assign onb = ~ONB;  //complement 
assign opb = ~OPB;  //complement 
assign nag = ~NAG;  //complement 
assign CHA = BAH & ACB ; 
assign cha = ~CHA ; //complement 
assign CHB = BAH & ACD ; 
assign chb = ~CHB ;  //complement 
assign CHC = BAH & ACF ; 
assign chc = ~CHC ;  //complement 
assign CHD = BAH & ACH; 
assign chd = ~CHD; 
assign nab = ~NAB;  //complement 
assign naj = ~NAJ;  //complement 
assign nai = ~NAI;  //complement 
assign CHE = BAH & ACJ ; 
assign che = ~CHE ; //complement 
assign CHF = BAH & ACL ; 
assign chf = ~CHF ;  //complement 
assign CHG = BAH & ACN ; 
assign chg = ~CHG ;  //complement 
assign CHH = BAH & ACP; 
assign chh = ~CHH; 
assign nak = ~NAK;  //complement 
assign nal = ~NAL;  //complement 
assign nam = ~NAM;  //complement 
assign CHI =  ADB & BAH  ; 
assign chi = ~CHI;  //complement 
assign CHJ =  ADD & BAH  ; 
assign chj = ~CHJ;  //complement 
assign CHK =  ADF & BAH  ; 
assign chk = ~CHK;  //complement 
assign nan = ~NAN;  //complement 
assign nao = ~NAO;  //complement 
assign nap = ~NAP;  //complement 
assign CHL =  ADH & BAH  ; 
assign chl = ~CHL;  //complement 
assign CHM =  ADJ & BAH  ; 
assign chm = ~CHM;  //complement 
assign GXC =  FXE  ; 
assign gxc = ~GXC;  //complement 
assign nbj = ~NBJ;  //complement 
assign nbk = ~NBK;  //complement 
assign nbm = ~NBM;  //complement 
assign CIA = BAI & ACA ; 
assign cia = ~CIA ; //complement 
assign CIB = BAI & ACC ; 
assign cib = ~CIB ;  //complement 
assign CIC = BAI & ACE ; 
assign cic = ~CIC ;  //complement 
assign CID = BAI & ACG; 
assign cid = ~CID; 
assign nbl = ~NBL;  //complement 
assign nbn = ~NBN;  //complement 
assign nbo = ~NBO;  //complement 
assign nbd = ~NBD;  //complement 
assign fyo = ~FYO;  //complement 
assign FYP = ~fyp;  //complement 
assign GZC =  FZE & fzg & fzb  |  fze & FZG & fzb  |  fze & fzg & FZB  |  FZE & FZG & FZB  ; 
assign gzc = ~GZC; //complement 
assign gzd =  FZE & fzg & fzb  |  fze & FZG & fzb  |  fze & fzg & FZB  |  fze & fzg & fzb  ; 
assign GZD = ~gzd;  //complement 
assign LHA =  HGA & kha  |  hga & KHA  ; 
assign lha = ~LHA;  //complement 
assign kzc = ~KZC;  //complement 
assign nbf = ~NBF;  //complement 
assign LIA =  KIA & hha & hhb  |  kia & HHA & hhb  |  kia & hha & HHB  |  KIA & HHA & HHB  ; 
assign lia = ~LIA; //complement 
assign lib =  KIA & hha & hhb  |  kia & HHA & hhb  |  kia & hha & HHB  |  kia & hha & hhb  ; 
assign LIB = ~lib;  //complement 
assign LJA =  KJA & kjb & hia  |  kja & KJB & hia  |  kja & kjb & HIA  |  KJA & KJB & HIA  ; 
assign lja = ~LJA; //complement 
assign ljb =  KJA & kjb & hia  |  kja & KJB & hia  |  kja & kjb & HIA  |  kja & kjb & hia  ; 
assign LJB = ~ljb;  //complement 
assign LZU =  HZT & hzv & hzr  |  hzt & HZV & hzr  |  hzt & hzv & HZR  |  HZT & HZV & HZR  ; 
assign lzu = ~LZU; //complement 
assign lzv =  HZT & hzv & hzr  |  hzt & HZV & hzr  |  hzt & hzv & HZR  |  hzt & hzv & hzr  ; 
assign LZV = ~lzv;  //complement 
assign nbh = ~NBH;  //complement 
assign LKA =  KMA & hja & hjb  |  kma & HJA & hjb  |  kma & hja & HJB  |  KMA & HJA & HJB  ; 
assign lka = ~LKA; //complement 
assign lkb =  KMA & hja & hjb  |  kma & HJA & hjb  |  kma & hja & HJB  |  kma & hja & hjb  ; 
assign LKB = ~lkb;  //complement 
assign LLA =  KNA & knb & hma  |  kna & KNB & hma  |  kna & knb & HMA  |  KNA & KNB & HMA  ; 
assign lla = ~LLA; //complement 
assign llb =  KNA & knb & hma  |  kna & KNB & hma  |  kna & knb & HMA  |  kna & knb & hma  ; 
assign LLB = ~llb;  //complement 
assign nfn = ~NFN;  //complement 
assign kwb = ~KWB;  //complement 
assign LMA =  KOA & hna & hnb  |  koa & HNA & hnb  |  koa & hna & HNB  |  KOA & HNA & HNB  ; 
assign lma = ~LMA; //complement 
assign lmb =  KOA & hna & hnb  |  koa & HNA & hnb  |  koa & hna & HNB  |  koa & hna & hnb  ; 
assign LMB = ~lmb;  //complement 
assign LNA =  HOA & kpa & kpb  |  hoa & KPA & kpb  |  hoa & kpa & KPB  |  HOA & KPA & KPB  ; 
assign lna = ~LNA; //complement 
assign lnb =  HOA & kpa & kpb  |  hoa & KPA & kpb  |  hoa & kpa & KPB  |  hoa & kpa & kpb  ; 
assign LNB = ~lnb;  //complement 
assign kyb = ~KYB;  //complement 
assign nbi = ~NBI;  //complement 
assign LOA =  HPA & hpb & kqa  |  hpa & HPB & kqa  |  hpa & hpb & KQA  |  HPA & HPB & KQA  ; 
assign loa = ~LOA; //complement 
assign lob =  HPA & hpb & kqa  |  hpa & HPB & kqa  |  hpa & hpb & KQA  |  hpa & hpb & kqa  ; 
assign LOB = ~lob;  //complement 
assign nfd = ~NFD;  //complement 
assign kvb = ~KVB;  //complement 
assign GWC =  FWD & fvd  |  fwd & FVD  ; 
assign gwc = ~GWC;  //complement 
assign LQA =  KRA & hqa & hqb  |  kra & HQA & hqb  |  kra & hqa & HQB  |  KRA & HQA & HQB  ; 
assign lqa = ~LQA; //complement 
assign lqb =  KRA & hqa & hqb  |  kra & HQA & hqb  |  kra & hqa & HQB  |  kra & hqa & hqb  ; 
assign LQB = ~lqb;  //complement 
assign GWD =  FWD & FVD  ; 
assign gwd = ~GWD;  //complement 
assign LHB =  HGA & KHA  ; 
assign lhb = ~LHB;  //complement 
assign nba = ~NBA;  //complement 
assign nfo = ~NFO;  //complement 
assign LSA =  KTA & hsa & hrb  |  kta & HSA & hrb  |  kta & hsa & HRB  |  KTA & HSA & HRB  ; 
assign lsa = ~LSA; //complement 
assign lsb =  KTA & hsa & hrb  |  kta & HSA & hrb  |  kta & hsa & HRB  |  kta & hsa & hrb  ; 
assign LSB = ~lsb;  //complement 
assign LTA =  KUA & hta & hsb  |  kua & HTA & hsb  |  kua & hta & HSB  |  KUA & HTA & HSB  ; 
assign lta = ~LTA; //complement 
assign ltb =  KUA & hta & hsb  |  kua & HTA & hsb  |  kua & hta & HSB  |  kua & hta & hsb  ; 
assign LTB = ~ltb;  //complement 
assign nfj = ~NFJ;  //complement 
assign LUA =  KVA & htb & hua  |  kva & HTB & hua  |  kva & htb & HUA  |  KVA & HTB & HUA  ; 
assign lua = ~LUA; //complement 
assign lub =  KVA & htb & hua  |  kva & HTB & hua  |  kva & htb & HUA  |  kva & htb & hua  ; 
assign LUB = ~lub;  //complement 
assign kzd = ~KZD;  //complement 
assign LVA =  HVA & hub & kwa  |  hva & HUB & kwa  |  hva & hub & KWA  |  HVA & HUB & KWA  ; 
assign lva = ~LVA; //complement 
assign lvb =  HVA & hub & kwa  |  hva & HUB & kwa  |  hva & hub & KWA  |  hva & hub & kwa  ; 
assign LVB = ~lvb;  //complement 
assign qzo = ~QZO;  //complement 
assign QZP = ~qzp;  //complement 
assign fzr = ~FZR;  //complement 
assign FZS = ~fzs;  //complement 
assign LRA =  KSA & ksb & hra  |  ksa & KSB & hra  |  ksa & ksb & HRA  |  KSA & KSB & HRA  ; 
assign lra = ~LRA; //complement 
assign lrb =  KSA & ksb & hra  |  ksa & KSB & hra  |  ksa & ksb & HRA  |  ksa & ksb & hra  ; 
assign LRB = ~lrb;  //complement 
assign EXG =  QXK & qxm & qxb  |  qxk & QXM & qxb  |  qxk & qxm & QXB  |  QXK & QXM & QXB  ; 
assign exg = ~EXG; //complement 
assign exh =  QXK & qxm & qxb  |  qxk & QXM & qxb  |  qxk & qxm & QXB  |  qxk & qxm & qxb  ; 
assign EXH = ~exh;  //complement 
assign qzq = ~QZQ;  //complement 
assign QZR = ~qzr;  //complement 
assign ojc = ~OJC;  //complement 
assign olc = ~OLC;  //complement 
assign onc = ~ONC;  //complement 
assign opc = ~OPC;  //complement 
assign NHC =  NEE & NAF  |  NEF  ; 
assign nhc = ~NHC;  //complement 
assign NHD =  NEE & NAF & NAG  |  NEF & NAG  |  NEG  ; 
assign nhd = ~NHD; //complement 
assign qzs = ~QZS;  //complement 
assign QZT = ~qzt;  //complement 
assign NHE =  NEE & NAF & NAG & NAH  |  NEF & NAG & NAH  |  NEG & NAH  |  NEH  ; 
assign nhe = ~NHE;  //complement 
assign NIC =  NEI & NAJ  |  NEJ  ; 
assign nic = ~NIC;  //complement 
assign NID =  NEI & NAJ & NAK  |  NEJ & NAK  |  NEK  ; 
assign nid = ~NID; //complement 
assign qxa = ~QXA;  //complement 
assign QXB = ~qxb;  //complement 
assign NIE =  NEI & NAJ & NAK & NAL  |  NEJ & NAK & NAL  |  NEK & NAL  |  NEL  ; 
assign nie = ~NIE;  //complement 
assign NJC =  NEM & NAN  |  NEN  ; 
assign njc = ~NJC;  //complement 
assign NJD =  NEM & NAN & NAO  |  NEN & NAO  |  NEO  ; 
assign njd = ~NJD; //complement 
assign qxc = ~QXC;  //complement 
assign QXD = ~qxd;  //complement 
assign NJE =  NEM & NAN & NAO & NAP  |  NEN & NAO & NAP  |  NEO & NAP  |  NEP  ; 
assign nje = ~NJE;  //complement 
assign NKC =  NAQ & NBB  |  NFB  ; 
assign nkc = ~NKC;  //complement 
assign NKD =  NAQ & NBB & NBC  |  NFB & NBC  |  NFC  ; 
assign nkd = ~NKD; //complement 
assign qxe = ~QXE;  //complement 
assign QXF = ~qxf;  //complement 
assign NKE =  NAQ & NBB & NBC & NBD  |  NFB & NBC & NBD  |  NFC & NBD  |  NFD  ; 
assign nke = ~NKE;  //complement 
assign NLC =  NFE & NBF  |  NFF  ; 
assign nlc = ~NLC;  //complement 
assign NLD =  NFE & NBF & NBG  |  NFF & NBG  |  NFG  ; 
assign nld = ~NLD; //complement 
assign qzk = ~QZK;  //complement 
assign QZL = ~qzl;  //complement 
assign nbp = ~NBP;  //complement 
assign nbe = ~NBE;  //complement 
assign NLE =  NFE & NBF & NBG & NBH  |  NFF & NBG & NBH  |  NFG & NBH  |  NFH  ; 
assign nle = ~NLE;  //complement 
assign qzm = ~QZM;  //complement 
assign QZN = ~qzn;  //complement 
assign nbg = ~NBG;  //complement 
assign mia = ~MIA;  //complement 
assign MIB = ~mib;  //complement 
assign ojh = ~OJH;  //complement 
assign olh = ~OLH;  //complement 
assign onh = ~ONH;  //complement 
assign oph = ~OPH;  //complement 
assign CIE = BAI & ACI ; 
assign cie = ~CIE ; //complement 
assign CIF = BAI & ACK ; 
assign cif = ~CIF ;  //complement 
assign CIG = BAI & ACM ; 
assign cig = ~CIG ;  //complement 
assign CIH = BAI & ACO; 
assign cih = ~CIH; 
assign LZX =  HZW & kzx & hzu  |  hzw & KZX & hzu  |  hzw & kzx & HZU  |  HZW & KZX & HZU  ; 
assign lzx = ~LZX; //complement 
assign lzy =  HZW & kzx & hzu  |  hzw & KZX & hzu  |  hzw & kzx & HZU  |  hzw & kzx & hzu  ; 
assign LZY = ~lzy;  //complement 
assign hxa = ~HXA;  //complement 
assign HXB = ~hxb;  //complement 
assign nfm = ~NFM;  //complement 
assign CJA =  BAJ & ACB  ; 
assign cja = ~CJA;  //complement 
assign LVC =  KVB  ; 
assign lvc = ~LVC;  //complement 
assign LZF =  HZB  ; 
assign lzf = ~LZF;  //complement 
assign mzu = ~MZU;  //complement 
assign MZV = ~mzv;  //complement 
assign mza = ~MZA;  //complement 
assign MZB = ~mzb;  //complement 
assign mzl = ~MZL;  //complement 
assign MZM = ~mzm;  //complement 
assign CII = BAI & ADA ; 
assign cii = ~CII ; //complement 
assign CIJ = BAI & ADC ; 
assign cij = ~CIJ ;  //complement 
assign CIK = BAI & ADE ; 
assign cik = ~CIK ;  //complement 
assign CIL = BAI & ADG; 
assign cil = ~CIL; 
assign mya = ~MYA;  //complement 
assign MYB = ~myb;  //complement 
assign kzg = ~KZG;  //complement 
assign mzi = ~MZI;  //complement 
assign MZJ = ~mzj;  //complement 
assign CJB =  BAJ & ACD  ; 
assign cjb = ~CJB;  //complement 
assign CJC =  BAJ & ACF  ; 
assign cjc = ~CJC;  //complement 
assign CJD =  BAJ & ACH  ; 
assign cjd = ~CJD;  //complement 
assign mzo = ~MZO;  //complement 
assign MZP = ~mzp;  //complement 
assign LZR =  KZT & hzq & hzn  |  kzt & HZQ & hzn  |  kzt & hzq & HZN  |  KZT & HZQ & HZN  ; 
assign lzr = ~LZR; //complement 
assign lzs =  KZT & hzq & hzn  |  kzt & HZQ & hzn  |  kzt & hzq & HZN  |  kzt & hzq & hzn  ; 
assign LZS = ~lzs;  //complement 
assign mzr = ~MZR;  //complement 
assign MZS = ~mzs;  //complement 
assign CJE =  BAJ & ACJ  ; 
assign cje = ~CJE;  //complement 
assign CJF =  BAJ & ACL  ; 
assign cjf = ~CJF;  //complement 
assign CJG =  BAJ & ACN  ; 
assign cjg = ~CJG;  //complement 
assign pbd = ~PBD;  //complement 
assign kub = ~KUB;  //complement 
assign ktb = ~KTB;  //complement 
assign CJH =  BAJ & ACP  ; 
assign cjh = ~CJH;  //complement 
assign CJI =  BAJ & ADB  ; 
assign cji = ~CJI;  //complement 
assign CJJ =  BAJ & ADD  ; 
assign cjj = ~CJJ;  //complement 
assign htb = ~HTB;  //complement 
assign mva = ~MVA;  //complement 
assign MVB = ~mvb;  //complement 
assign kya = ~KYA;  //complement 
assign CJK =  BAJ & ADF  ; 
assign cjk = ~CJK;  //complement 
assign CJL =  BAJ & ADH  ; 
assign cjl = ~CJL;  //complement 
assign CKA =  BAK & ACA  ; 
assign cka = ~CKA;  //complement 
assign NMC =  NFI & NBJ  |  NFJ  ; 
assign nmc = ~NMC;  //complement 
assign NMD =  NFI & NBJ & NBK  |  NFJ & NBK  |  NFK  ; 
assign nmd = ~NMD; //complement 
assign hva = ~HVA;  //complement 
assign HVB = ~hvb;  //complement 
assign CKB =  BAK & ACC  ; 
assign ckb = ~CKB;  //complement 
assign CKC =  BAK & ACE  ; 
assign ckc = ~CKC;  //complement 
assign CKD =  BAK & ACG  ; 
assign ckd = ~CKD;  //complement 
assign mmb = ~MMB;  //complement 
assign hwa = ~HWA;  //complement 
assign HWB = ~hwb;  //complement 
assign NME =  NFI & NBJ & NBK & NBL  |  NFJ & NBK & NBL  |  NFK & NBL  |  NFL  ; 
assign nme = ~NME;  //complement 
assign oji = ~OJI;  //complement 
assign oli = ~OLI;  //complement 
assign oni = ~ONI;  //complement 
assign opi = ~OPI;  //complement 
assign pbf = ~PBF;  //complement 
assign LWA =  HWA & hvb & kxa  |  hwa & HVB & kxa  |  hwa & hvb & KXA  |  HWA & HVB & KXA  ; 
assign lwa = ~LWA; //complement 
assign lwb =  HWA & hvb & kxa  |  hwa & HVB & kxa  |  hwa & hvb & KXA  |  hwa & hvb & kxa  ; 
assign LWB = ~lwb;  //complement 
assign LXA =  HXA & hwb & kya  |  hxa & HWB & kya  |  hxa & hwb & KYA  |  HXA & HWB & KYA  ; 
assign lxa = ~LXA; //complement 
assign lxb =  HXA & hwb & kya  |  hxa & HWB & kya  |  hxa & hwb & KYA  |  hxa & hwb & kya  ; 
assign LXB = ~lxb;  //complement 
assign LZI =  KZI & hzd & hzg  |  kzi & HZD & hzg  |  kzi & hzd & HZG  |  KZI & HZD & HZG  ; 
assign lzi = ~LZI; //complement 
assign lzj =  KZI & hzd & hzg  |  kzi & HZD & hzg  |  kzi & hzd & HZG  |  kzi & hzd & hzg  ; 
assign LZJ = ~lzj;  //complement 
assign pbg = ~PBG;  //complement 
assign meb = ~MEB;  //complement 
assign LZA =  HZA & hyb & kzc  |  hza & HYB & kzc  |  hza & hyb & KZC  |  HZA & HYB & KZC  ; 
assign lza = ~LZA; //complement 
assign lzb =  HZA & hyb & kzc  |  hza & HYB & kzc  |  hza & hyb & KZC  |  hza & hyb & kzc  ; 
assign LZB = ~lzb;  //complement 
assign mga = ~MGA;  //complement 
assign fvc = ~FVC;  //complement 
assign FVD = ~fvd;  //complement 
assign ojd = ~OJD;  //complement 
assign old = ~OLD;  //complement 
assign ond = ~OND;  //complement 
assign opd = ~OPD;  //complement 
assign LZD =  KZD & kzg & hzc  |  kzd & KZG & hzc  |  kzd & kzg & HZC  |  KZD & KZG & HZC  ; 
assign lzd = ~LZD; //complement 
assign lze =  KZD & kzg & hzc  |  kzd & KZG & hzc  |  kzd & kzg & HZC  |  kzd & kzg & hzc  ; 
assign LZE = ~lze;  //complement 
assign mgb = ~MGB;  //complement 
assign hzm = ~HZM;  //complement 
assign HZN = ~hzn;  //complement 
assign NLB =  NFE  ; 
assign nlb = ~NLB;  //complement 
assign LTC =  KTB  ; 
assign ltc = ~LTC;  //complement 
assign LWC =  KWB  ; 
assign lwc = ~LWC;  //complement 
assign oje = ~OJE;  //complement 
assign ole = ~OLE;  //complement 
assign one = ~ONE;  //complement 
assign ope = ~OPE;  //complement 
assign NND =  NFM & NBN & NBO  |  NFN & NBO  |  NFO  ; 
assign nnd = ~NND; //complement 
assign NNE =  NFM & NBN & NBO & NBP  |  NFN & NBO & NBP  |  NFO & NBP  |  NFP  ; 
assign nne = ~NNE;  //complement 
assign hzi = ~HZI;  //complement 
assign HZJ = ~hzj;  //complement 
assign mha = ~MHA;  //complement 
assign NJB =  NEM  ; 
assign njb = ~NJB;  //complement 
assign NHB =  NEE  ; 
assign nhb = ~NHB;  //complement 
assign NGD =  NEB & NAC  ; 
assign ngd = ~NGD;  //complement 
assign pbh = ~PBH;  //complement 
assign fzw = ~FZW;  //complement 
assign FZX = ~fzx;  //complement 
assign NGE =  NEB & NAC & NAD  ; 
assign nge = ~NGE;  //complement 
assign LXC =  KXB  ; 
assign lxc = ~LXC;  //complement 
assign LZN =  KZM  ; 
assign lzn = ~LZN;  //complement 
assign ffa = ~FFA;  //complement 
assign hya = ~HYA;  //complement 
assign HYB = ~hyb;  //complement 
assign ffb = ~FFB;  //complement 
assign fys = ~FYS;  //complement 
assign nud =  nfj & nfk & nbi  |  nfk & nbj  |  nbk  ; 
assign NUD = ~nud; //complement 
assign GZA =  FZA & fzc & fyb  |  fza & FZC & fyb  |  fza & fzc & FYB  |  FZA & FZC & FYB  ; 
assign gza = ~GZA; //complement 
assign gzb =  FZA & fzc & fyb  |  fza & FZC & fyb  |  fza & fzc & FYB  |  fza & fzc & fyb  ; 
assign GZB = ~gzb;  //complement 
assign kza = ~KZA;  //complement 
assign kzb = ~KZB;  //complement 
assign qxk = ~QXK;  //complement 
assign QXL = ~qxl;  //complement 
assign qyr = ~QYR;  //complement 
assign pfk = ~PFK;  //complement 
assign pfl = ~PFL;  //complement 
assign pfm = ~PFM;  //complement 
assign pfn = ~PFN;  //complement 
assign qxm = ~QXM;  //complement 
assign QXN = ~qxn;  //complement 
assign pbj = ~PBJ;  //complement 
assign pfo = ~PFO;  //complement 
assign pfp = ~PFP;  //complement 
assign pga = ~PGA;  //complement 
assign pgb = ~PGB;  //complement 
assign qxo = ~QXO;  //complement 
assign QXP = ~qxp;  //complement 
assign pgc = ~PGC;  //complement 
assign pgd = ~PGD;  //complement 
assign pge = ~PGE;  //complement 
assign pgf = ~PGF;  //complement 
assign pgg = ~PGG;  //complement 
assign pgh = ~PGH;  //complement 
assign qxq = ~QXQ;  //complement 
assign QXR = ~qxr;  //complement 
assign pbk = ~PBK;  //complement 
assign pgi = ~PGI;  //complement 
assign pgk = ~PGK;  //complement 
assign qxs = ~QXS;  //complement 
assign QXT = ~qxt;  //complement 
assign pgm = ~PGM;  //complement 
assign pgo = ~PGO;  //complement 
assign pbl = ~PBL;  //complement 
assign qxv = ~QXV;  //complement 
assign QXW = ~qxw;  //complement 
assign pbn = ~PBN;  //complement 
assign pbo = ~PBO;  //complement 
assign pbp = ~PBP;  //complement 
assign qxg = ~QXG;  //complement 
assign QXH = ~qxh;  //complement 
assign mhb = ~MHB;  //complement 
assign mnb = ~MNB;  //complement 
assign qxi = ~QXI;  //complement 
assign QXJ = ~qxj;  //complement 
assign pfe = ~PFE;  //complement 
assign pff = ~PFF;  //complement 
assign pfg = ~PFG;  //complement 
assign pfh = ~PFH;  //complement 
assign pfi = ~PFI;  //complement 
assign pfj = ~PFJ;  //complement 
assign CKE =  BAK & ACI  ; 
assign cke = ~CKE;  //complement 
assign CKF =  BAK & ACK  ; 
assign ckf = ~CKF;  //complement 
assign CKG =  BAK & ACM  ; 
assign ckg = ~CKG;  //complement 
assign GZX =  FYJ & fyl & fyf  |  fyj & FYL & fyf  |  fyj & fyl & FYF  |  FYJ & FYL & FYF  ; 
assign gzx = ~GZX; //complement 
assign gzy =  FYJ & fyl & fyf  |  fyj & FYL & fyf  |  fyj & fyl & FYF  |  fyj & fyl & fyf  ; 
assign GZY = ~gzy;  //complement 
assign LYC =  KYB  ; 
assign lyc = ~LYC;  //complement 
assign hjb = ~HJB;  //complement 
assign hpb = ~HPB;  //complement 
assign hpa = ~HPA;  //complement 
assign hqa = ~HQA;  //complement 
assign CKH =  BAK & ACO  ; 
assign ckh = ~CKH;  //complement 
assign CKI =  BAK & ADA  ; 
assign cki = ~CKI;  //complement 
assign CKJ =  BAK & ADC  ; 
assign ckj = ~CKJ;  //complement 
assign dzq = ~DZQ;  //complement 
assign ELC = DLD; 
assign elc = ~ELC; //complement 
assign EBA =  DGB  ; 
assign eba = ~EBA;  //complement 
assign EAA =  DGA  ; 
assign eaa = ~EAA;  //complement 
assign EOD =  DND  ; 
assign eod = ~EOD;  //complement 
assign CKK =  BAK & ADE  ; 
assign ckk = ~CKK;  //complement 
assign CLA =  BAL & ACB  ; 
assign cla = ~CLA;  //complement 
assign CLB =  BAL & ACD  ; 
assign clb = ~CLB;  //complement 
assign fhb = ~FHB;  //complement 
assign hqb = ~HQB;  //complement 
assign fud = ~FUD;  //complement 
assign LZL =  KZJ & hzi & hzh  |  kzj & HZI & hzh  |  kzj & hzi & HZH  |  KZJ & HZI & HZH  ; 
assign lzl = ~LZL; //complement 
assign lzm =  KZJ & hzi & hzh  |  kzj & HZI & hzh  |  kzj & hzi & HZH  |  kzj & hzi & hzh  ; 
assign LZM = ~lzm;  //complement 
assign hsa = ~HSA;  //complement 
assign HSB = ~hsb;  //complement 
assign CLC =  BAL & ACF  ; 
assign clc = ~CLC;  //complement 
assign CLD =  BAL & ACH  ; 
assign cld = ~CLD;  //complement 
assign CLE =  BAL & ACJ  ; 
assign cle = ~CLE;  //complement 
assign LOC = KQB; 
assign loc = ~LOC; //complement 
assign LSC = ZZO; 
assign lsc = ~LSC; //complement 
assign kzh = ~KZH;  //complement 
assign CLF =  BAL & ACL  ; 
assign clf = ~CLF;  //complement 
assign CLG =  BAL & ACN  ; 
assign clg = ~CLG;  //complement 
assign CLH =  BAL & ACP  ; 
assign clh = ~CLH;  //complement 
assign pba = ~PBA;  //complement 
assign pbb = ~PBB;  //complement 
assign pbe = ~PBE;  //complement 
assign pbi = ~PBI;  //complement 
assign pbm = ~PBM;  //complement 
assign pca = ~PCA;  //complement 
assign pce = ~PCE;  //complement 
assign pci = ~PCI;  //complement 
assign pcm = ~PCM;  //complement 
assign pde = ~PDE;  //complement 
assign CLI =  BAL & ADB  ; 
assign cli = ~CLI;  //complement 
assign CLJ =  BAL & ADD  ; 
assign clj = ~CLJ;  //complement 
assign CLK =  BAL & ADF  ; 
assign clk = ~CLK;  //complement 
assign pdi = ~PDI;  //complement 
assign pdm = ~PDM;  //complement 
assign pea = ~PEA;  //complement 
assign pee = ~PEE;  //complement 
assign pei = ~PEI;  //complement 
assign pem = ~PEM;  //complement 
assign paf = ~PAF;  //complement 
assign CMA =  BAM & ACA  ; 
assign cma = ~CMA;  //complement 
assign CMB =  BAM & ACC  ; 
assign cmb = ~CMB;  //complement 
assign CMC =  BAM & ACE  ; 
assign cmc = ~CMC;  //complement 
assign pcb = ~PCB;  //complement 
assign pcc = ~PCC;  //complement 
assign pcd = ~PCD;  //complement 
assign CMD =  BAM & ACG  ; 
assign cmd = ~CMD;  //complement 
assign CME =  BAM & ACI  ; 
assign cme = ~CME;  //complement 
assign CMF =  BAM & ACK  ; 
assign cmf = ~CMF;  //complement 
assign pcf = ~PCF;  //complement 
assign pcg = ~PCG;  //complement 
assign pch = ~PCH;  //complement 
assign peo = ~PEO;  //complement 
assign pen = ~PEN;  //complement 
assign pah = ~PAH;  //complement 
assign neo = ~NEO;  //complement 
assign qaa = ~QAA;  //complement 
assign qab = ~QAB;  //complement 
assign qac = ~QAC;  //complement 
assign qad = ~QAD;  //complement 
assign TEA = QAB; 
assign tea = ~TEA; //complement 
assign TEB = QAB; 
assign teb = ~TEB;  //complement 
assign TEC = QAB; 
assign tec = ~TEC;  //complement 
assign TED = QAB; 
assign ted = ~TED;  //complement 
assign qae = ~QAE;  //complement 
assign qaf = ~QAF;  //complement 
assign qag = ~QAG;  //complement 
assign qah = ~QAH;  //complement 
assign nee = ~NEE;  //complement 
assign oea = ~OEA;  //complement 
assign oeb = ~OEB;  //complement 
assign oec = ~OEC;  //complement 
assign oed = ~OED;  //complement 
assign oee = ~OEE;  //complement 
assign oef = ~OEF;  //complement 
assign ofa = ~OFA;  //complement 
assign ofb = ~OFB;  //complement 
assign ofc = ~OFC;  //complement 
assign ofd = ~OFD;  //complement 
assign ofe = ~OFE;  //complement 
assign off = ~OFF;  //complement 
assign fyd = ~FYD;  //complement 
assign OHC = ~ohc;  //complement 
assign OHD = ~ohd;  //complement 
assign OHE = ~ohe;  //complement 
assign OGA = ~oga;  //complement 
assign OGB = ~ogb;  //complement 
assign OGC = ~ogc;  //complement 
assign OGD = ~ogd;  //complement 
assign OGE = ~oge;  //complement 
assign OGF = ~ogf;  //complement 
assign OHA = ~oha;  //complement 
assign OHB = ~ohb;  //complement 
assign LIC =  HGB & khb  |  hgb & KHB  ; 
assign lic = ~LIC;  //complement 
assign OIG = ~oig;  //complement 
assign OKG = ~okg;  //complement 
assign OMG = ~omg;  //complement 
assign OOG = ~oog;  //complement 
assign qai = ~QAI;  //complement 
assign qaj = ~QAJ;  //complement 
assign qak = ~QAK;  //complement 
assign qal = ~QAL;  //complement 
assign TEE =  QAA  |  QAB  |  QAC  ; 
assign tee = ~TEE;  //complement 
assign TEF =  QAA  |  QAB  |  QAC  ; 
assign tef = ~TEF; //complement 
assign TEG =  QAA  |  QAB  |  QAC  ; 
assign teg = ~TEG;  //complement 
assign TEH =  QAA  |  QAB  |  QAC  ; 
assign teh = ~TEH;  //complement 
assign ace = ~ACE;  //complement 
assign acf = ~ACF;  //complement 
assign acg = ~ACG;  //complement 
assign ach = ~ACH;  //complement 
assign aci = ~ACI;  //complement 
assign acj = ~ACJ;  //complement 
assign ack = ~ACK;  //complement 
assign acl = ~ACL;  //complement 
assign acm = ~ACM;  //complement 
assign acn = ~ACN;  //complement 
assign aco = ~ACO;  //complement 
assign acp = ~ACP;  //complement 
assign nej = ~NEJ;  //complement 
assign pcj = ~PCJ;  //complement 
assign pck = ~PCK;  //complement 
assign pcl = ~PCL;  //complement 
assign pcn = ~PCN;  //complement 
assign pco = ~PCO;  //complement 
assign pcp = ~PCP;  //complement 
assign pbc = ~PBC;  //complement 
assign RAE =  NAE & nee  ; 
assign rae = ~RAE;  //complement 
assign RAF =  NAF & nef  ; 
assign raf = ~RAF;  //complement 
assign RAG =  NAG & neg  ; 
assign rag = ~RAG;  //complement 
assign qvb = ~QVB;  //complement 
assign QVC = ~qvc;  //complement 
assign bag = ~BAG;  //complement 
assign bah = ~BAH;  //complement 
assign bao = ~BAO;  //complement 
assign bap = ~BAP;  //complement 
assign bbo = ~BBO;  //complement 
assign bbp = ~BBP;  //complement 
assign qvd = ~QVD;  //complement 
assign QVE = ~qve;  //complement 
assign bbg = ~BBG;  //complement 
assign bbh = ~BBH;  //complement 
assign ECB =  DHB  ; 
assign ecb = ~ECB;  //complement 
assign EKC =  DKD  ; 
assign ekc = ~EKC;  //complement 
assign RAH =  NAH & neh  ; 
assign rah = ~RAH;  //complement 
assign nxg =  nbi  |  nbj  |  nbk  |  nbl  ;
assign NXG = ~nxg;  //complement 
assign EYS =  QXA & qxc & qzl  |  qxa & QXC & qzl  |  qxa & qxc & QZL  |  QXA & QXC & QZL  ; 
assign eys = ~EYS; //complement 
assign eyt =  QXA & qxc & qzl  |  qxa & QXC & qzl  |  qxa & qxc & QZL  |  qxa & qxc & qzl  ; 
assign EYT = ~eyt;  //complement 
assign nxi =  nae  |  naf  |  nag  |  nah  |  nai  ;
assign NXI = ~nxi;  //complement 
assign nxj =  naj  |  nak  |  nal  |  nam  |  nan  ;
assign NXJ = ~nxj;  //complement 
assign nxk =  nao  |  nap  |  nba  |  nbb  |  nbc  ;
assign NXK = ~nxk;  //complement 
assign hcb = ~HCB;  //complement 
assign hdb = ~HDB;  //complement 
assign nxl =  nbd  |  nbe  |  nbf  |  nbg  |  nbh  ;
assign NXL = ~nxl;  //complement 
assign NIB =  NEI  ; 
assign nib = ~NIB;  //complement 
assign NMB =  NFI  ; 
assign nmb = ~NMB;  //complement 
assign ojk = ~OJK;  //complement 
assign olk = ~OLK;  //complement 
assign onk = ~ONK;  //complement 
assign opk = ~OPK;  //complement 
assign LZO =  HZM & kzn & hzj  |  hzm & KZN & hzj  |  hzm & kzn & HZJ  |  HZM & KZN & HZJ  ; 
assign lzo = ~LZO; //complement 
assign lzp =  HZM & kzn & hzj  |  hzm & KZN & hzj  |  hzm & kzn & HZJ  |  hzm & kzn & hzj  ; 
assign LZP = ~lzp;  //complement 
assign ojl = ~OJL;  //complement 
assign oll = ~OLL;  //complement 
assign onl = ~ONL;  //complement 
assign opl = ~OPL;  //complement 
assign ojf = ~OJF;  //complement 
assign olf = ~OLF;  //complement 
assign onf = ~ONF;  //complement 
assign opf = ~OPF;  //complement 
assign hga = ~HGA;  //complement 
assign hgb = ~HGB;  //complement 
assign naf = ~NAF;  //complement 
assign hha = ~HHA;  //complement 
assign hhb = ~HHB;  //complement 
assign ojj = ~OJJ;  //complement 
assign olj = ~OLJ;  //complement 
assign onj = ~ONJ;  //complement 
assign opj = ~OPJ;  //complement 
assign qxx = ~QXX;  //complement 
assign QXY = ~qxy;  //complement 
assign acq = ~ACQ;  //complement 
assign pgn = ~PGN;  //complement 
assign pgp = ~PGP;  //complement 
assign qxz = ~QXZ;  //complement 
assign QVA = ~qva;  //complement 
assign tfa = ~TFA;  //complement 
assign tfb = ~TFB;  //complement 
assign tfc = ~TFC;  //complement 
assign tfd = ~TFD;  //complement 
assign hzt = ~HZT;  //complement 
assign HZU = ~hzu;  //complement 
assign neg = ~NEG;  //complement 
assign CMG =  BAM & ACM  ; 
assign cmg = ~CMG;  //complement 
assign CMH =  BAM & ACO  ; 
assign cmh = ~CMH;  //complement 
assign CMI =  BAM & ADA  ; 
assign cmi = ~CMI;  //complement 
assign fzt = ~FZT;  //complement 
assign FZU = ~fzu;  //complement 
assign GZO =  FZP & fzv  |  fzp & FZV  ; 
assign gzo = ~GZO;  //complement 
assign CMJ =  BAM & ADC  ; 
assign cmj = ~CMJ;  //complement 
assign CNA =  BAN & ACB  ; 
assign cna = ~CNA;  //complement 
assign CNB =  BAN & ACD  ; 
assign cnb = ~CNB;  //complement 
assign JZT =  HZT & hzv & hzr  |  hzt & HZV & hzr  |  hzt & hzv & HZR  |  HZT & HZV & HZR  ; 
assign jzt = ~JZT; //complement 
assign jzu =  HZT & hzv & hzr  |  hzt & HZV & hzr  |  hzt & hzv & HZR  |  hzt & hzv & hzr  ; 
assign JZU = ~jzu;  //complement 
assign LZK =  KZH  ; 
assign lzk = ~LZK;  //complement 
assign hza = ~HZA;  //complement 
assign HZB = ~hzb;  //complement 
assign gzk = ~GZK;  //complement 
assign CNC =  BAN & ACF  ; 
assign cnc = ~CNC;  //complement 
assign CND =  BAN & ACH  ; 
assign cnd = ~CND;  //complement 
assign CNE =  BAN & ACJ  ; 
assign cne = ~CNE;  //complement 
assign nvb =  nbm  ; 
assign NVB = ~nvb;  //complement 
assign nvc =  nfn & nbm  |  nbn  ; 
assign NVC = ~nvc;  //complement 
assign pag = ~PAG;  //complement 
assign ada = ~ADA;  //complement 
assign adb = ~ADB;  //complement 
assign adc = ~ADC;  //complement 
assign add = ~ADD;  //complement 
assign CNF =  BAN & ACL  ; 
assign cnf = ~CNF;  //complement 
assign CNG =  BAN & ACN  ; 
assign cng = ~CNG;  //complement 
assign CNH =  BAN & ACP  ; 
assign cnh = ~CNH;  //complement 
assign nvd =  nfn & nfo & nbm  |  nfo & nbn  |  nbo  ; 
assign NVD = ~nvd; //complement 
assign ade = ~ADE;  //complement 
assign adf = ~ADF;  //complement 
assign adg = ~ADG;  //complement 
assign adh = ~ADH;  //complement 
assign PAI = ~pai;  //complement 
assign CNI =  BAN & ADB  ; 
assign cni = ~CNI;  //complement 
assign CNJ =  BAN & ADD  ; 
assign cnj = ~CNJ;  //complement 
assign COA =  BAO & ACA  ; 
assign coa = ~COA;  //complement 
assign adi = ~ADI;  //complement 
assign adj = ~ADJ;  //complement 
assign adk = ~ADK;  //complement 
assign adl = ~ADL;  //complement 
assign nrd =  neo & nen & nam  |  neo & nan  |  nao  ; 
assign NRD = ~nrd; //complement 
assign nef = ~NEF;  //complement 
assign COB =  BAO & ACC  ; 
assign cob = ~COB;  //complement 
assign COC =  BAO & ACE  ; 
assign coc = ~COC;  //complement 
assign COD =  BAO & ACG  ; 
assign cod = ~COD;  //complement 
assign pef = ~PEF;  //complement 
assign adm = ~ADM;  //complement 
assign adn = ~ADN;  //complement 
assign ado = ~ADO;  //complement 
assign adp = ~ADP;  //complement 
assign aca = ~ACA;  //complement 
assign acb = ~ACB;  //complement 
assign acc = ~ACC;  //complement 
assign acd = ~ACD;  //complement 
assign COE =  BAO & ACI  ; 
assign coe = ~COE;  //complement 
assign COF =  BAO & ACK  ; 
assign cof = ~COF;  //complement 
assign COG =  BAO & ACM  ; 
assign cog = ~COG;  //complement 
assign EFB =  DHF  ; 
assign efb = ~EFB;  //complement 
assign PAM =  PAO & PAI & PAL  |  PAQ & PAI  ; 
assign pam = ~PAM;  //complement 
assign maa = ~MAA;  //complement 
assign mca = ~MCA;  //complement 
assign COH =  BAO & ACO  ; 
assign coh = ~COH;  //complement 
assign COI =  BAO & ADA  ; 
assign coi = ~COI;  //complement 
assign CPA =  BAP & ACB  ; 
assign cpa = ~CPA;  //complement 
assign pgj = ~PGJ;  //complement 
assign pgl = ~PGL;  //complement 
assign ojm = ~OJM;  //complement 
assign olm = ~OLM;  //complement 
assign onm = ~ONM;  //complement 
assign opm = ~OPM;  //complement 
assign iaa = ~IAA; //complement 
assign iab = ~IAB; //complement 
assign iac = ~IAC; //complement 
assign iad = ~IAD; //complement 
assign iae = ~IAE; //complement 
assign iaf = ~IAF; //complement 
assign iag = ~IAG; //complement 
assign iah = ~IAH; //complement 
assign iai = ~IAI; //complement 
assign iaj = ~IAJ; //complement 
assign iak = ~IAK; //complement 
assign ial = ~IAL; //complement 
assign iam = ~IAM; //complement 
assign ian = ~IAN; //complement 
assign iao = ~IAO; //complement 
assign iap = ~IAP; //complement 
assign iba = ~IBA; //complement 
assign ibb = ~IBB; //complement 
assign ibc = ~IBC; //complement 
assign ibd = ~IBD; //complement 
assign ibe = ~IBE; //complement 
assign ibf = ~IBF; //complement 
assign ibg = ~IBG; //complement 
assign ibh = ~IBH; //complement 
assign ibi = ~IBI; //complement 
assign ibj = ~IBJ; //complement 
assign ibk = ~IBK; //complement 
assign ibl = ~IBL; //complement 
assign ibm = ~IBM; //complement 
assign ibn = ~IBN; //complement 
assign ibo = ~IBO; //complement 
assign ibp = ~IBP; //complement 
assign ica = ~ICA; //complement 
assign icb = ~ICB; //complement 
assign icc = ~ICC; //complement 
assign icd = ~ICD; //complement 
assign ice = ~ICE; //complement 
assign icf = ~ICF; //complement 
assign icg = ~ICG; //complement 
assign ich = ~ICH; //complement 
assign ici = ~ICI; //complement 
assign icj = ~ICJ; //complement 
assign ick = ~ICK; //complement 
assign icl = ~ICL; //complement 
assign icm = ~ICM; //complement 
assign icn = ~ICN; //complement 
assign ico = ~ICO; //complement 
assign icp = ~ICP; //complement 
assign ida = ~IDA; //complement 
assign idb = ~IDB; //complement 
assign idc = ~IDC; //complement 
assign idd = ~IDD; //complement 
assign ide = ~IDE; //complement 
assign idf = ~IDF; //complement 
assign idg = ~IDG; //complement 
assign idh = ~IDH; //complement 
assign idi = ~IDI; //complement 
assign idj = ~IDJ; //complement 
assign idk = ~IDK; //complement 
assign idl = ~IDL; //complement 
assign idm = ~IDM; //complement 
assign idn = ~IDN; //complement 
assign ido = ~IDO; //complement 
assign idp = ~IDP; //complement 
assign iea = ~IEA; //complement 
assign ieb = ~IEB; //complement 
assign iec = ~IEC; //complement 
assign ied = ~IED; //complement 
assign iee = ~IEE; //complement 
assign ief = ~IEF; //complement 
assign ifa = ~IFA; //complement 
assign ifb = ~IFB; //complement 
assign ifc = ~IFC; //complement 
assign ifd = ~IFD; //complement 
assign ife = ~IFE; //complement 
assign iiff = ~IIFF; //complement 
assign ifg = ~IFG; //complement 
assign iga = ~IGA; //complement 
assign igb = ~IGB; //complement 
assign igc = ~IGC; //complement 
assign igd = ~IGD; //complement 
assign ige = ~IGE; //complement 
assign igf = ~IGF; //complement 
assign iha = ~IHA; //complement 
always@(posedge IZZ )
   begin 
 AAL <= IAL & teb |  AAM & TEB ; 
 AAM <= IAM & teb |  AAN & TEB ; 
 AAN <= IAN & teb |  AAO & TEB ; 
 AAO <= IAO & teb |  AAP & TEB ; 
 AAP <= IAP & teb |  ABA & TEB ; 
 DHB <= CCA ; 
 QXU <= DEA ; 
 FTC <= ZZO ; 
 PAO <= NGE ; 
 DHC <= CBB ; 
 DHD <= CDA ; 
 DKC <= CGB ; 
 DKD <= CIA ; 
 OJG <= IFG ; 
 OLG <= IFG ; 
 ONG <= IFG ; 
 OPG <= IFG ; 
 NEB <= MBB & MBA ; 
 DIC <=  CAD & ccc & ceb  |  cad & CCC & ceb  |  cad & ccc & CEB  |  CAD & CCC & CEB  ;
 did <=  CAD & ccc & ceb  |  cad & CCC & ceb  |  cad & ccc & CEB  |  cad & ccc & ceb  ;
 DHA <= CAB ; 
 FYN <= EYX ; 
 KCB <= HCB ; 
 KDB <= HDB ; 
 DGA <= CAA ; 
 DGB <= CBA ; 
 DPE <= CNA ; 
 QYI <= CZA ; 
 NBC <=  MTA  |  MSB  ; 
 DJA <=  CBD & cdc & cfb  |  cbd & CDC & cfb  |  cbd & cdc & CFB  |  CBD & CDC & CFB  ;
 djb <=  CBD & cdc & cfb  |  cbd & CDC & cfb  |  cbd & cdc & CFB  |  cbd & cdc & cfb  ;
 FZA <=  EZA & ezc & eze  |  eza & EZC & eze  |  eza & ezc & EZE  |  EZA & EZC & EZE  ;
 fzb <=  EZA & ezc & eze  |  eza & EZC & eze  |  eza & ezc & EZE  |  eza & ezc & eze  ;
 NBB <=  MSA  |  MRB  ; 
 DKA <=  CAE & ccd & cec  |  cae & CCD & cec  |  cae & ccd & CEC  |  CAE & CCD & CEC  ;
 dkb <=  CAE & ccd & cec  |  cae & CCD & cec  |  cae & ccd & CEC  |  cae & ccd & cec  ;
 DWG <= CSB ; 
 DWH <= CUA ; 
 DXG <= CTB ; 
 DXH <= CVA ; 
 DIE <= CGA ; 
 DJC <= CHA ; 
 DUG <= CSA ; 
 HEA <= FEA ; 
 MDA <=  LDA & ldc & lcb  |  lda & LDC & lcb  |  lda & ldc & LCB  |  LDA & LDC & LCB  ;
 mdb <=  LDA & ldc & lcb  |  lda & LDC & lcb  |  lda & ldc & LCB  |  lda & ldc & lcb  ;
 DLA <=  CBE & cdd & cfc  |  cbe & CDD & cfc  |  cbe & cdd & CFC  |  CBE & CDD & CFC  ;
 dlb <=  CBE & cdd & cfc  |  cbe & CDD & cfc  |  cbe & cdd & CFC  |  cbe & cdd & cfc  ;
 NFP <= MZV & MZX ; 
 MZX <=  LZX & lzz & lzv  |  lzx & LZZ & lzv  |  lzx & lzz & LZV  |  LZX & LZZ & LZV  ;
 mzy <=  LZX & lzz & lzv  |  lzx & LZZ & lzv  |  lzx & lzz & LZV  |  lzx & lzz & lzv  ;
 DMA <=  CAF & cce & ced  |  caf & CCE & ced  |  caf & cce & CED  |  CAF & CCE & CED  ;
 dmb <=  CAF & cce & ced  |  caf & CCE & ced  |  caf & cce & CED  |  caf & cce & ced  ;
 AAA <= IAA & tea |  AAB & TEA ; 
 AAB <= IAB & tea |  AAC & TEA ; 
 AAC <= IAC & tea |  AAD & TEA ; 
 AAD <= IAD & tea |  AAE & TEA ; 
 AAE <= IAE & tea |  AAF & TEA ; 
 AAF <= IAF & tea |  AAG & TEA ; 
 AAG <= IAG & tea |  AAH & TEA ; 
 AAH <= IAH & tea |  AAI & TEA ; 
 AAI <= IAI & teb |  AAJ & TEB ; 
 AAJ <= IAJ & teb |  AAK & TEB ; 
 AAK <= IAK & teb |  AAL & TEB ; 
 DHE <=  CAC & ccb & cea  |  cac & CCB & cea  |  cac & ccb & CEA  |  CAC & CCB & CEA  ;
 dhf <=  CAC & ccb & cea  |  cac & CCB & cea  |  cac & ccb & CEA  |  cac & ccb & cea  ;
 DIA <=  CBC & cdb & cfa  |  cbc & CDB & cfa  |  cbc & cdb & CFA  |  CBC & CDB & CFA  ;
 dib <=  CBC & cdb & cfa  |  cbc & CDB & cfa  |  cbc & cdb & CFA  |  cbc & cdb & cfa  ;
 DNC <=  CHC & cjb & cla  |  chc & CJB & cla  |  chc & cjb & CLA  |  CHC & CJB & CLA  ;
 dnd <=  CHC & cjb & cla  |  chc & CJB & cla  |  chc & cjb & CLA  |  chc & cjb & cla  ;
 ABG <= IBG & tec |  ABH & TEC ; 
 ABH <= IBH & tec |  ABI & TEC ; 
 DOA <=  CAG & ccf & cee  |  cag & CCF & cee  |  cag & ccf & CEE  |  CAG & CCF & CEE  ;
 dob <=  CAG & ccf & cee  |  cag & CCF & cee  |  cag & ccf & CEE  |  cag & ccf & cee  ;
 ABI <= IBI & ted |  ABJ & TED ; 
 ABJ <= IBJ & ted |  ABK & TED ; 
 ABK <= IBK & ted |  ABL & TED ; 
 HJA <= FJA ; 
 HIA <= FIA ; 
 HMA <= GMA ; 
 MBA <= LBA ; 
 DOC <=  CGD & cic & ckb  |  cgd & CIC & ckb  |  cgd & cic & CKB  |  CGD & CIC & CKB  ;
 dod <=  CGD & cic & ckb  |  cgd & CIC & ckb  |  cgd & cic & CKB  |  cgd & cic & ckb  ;
 ABL <= IBL & ted |  ABM & TED ; 
 ABM <= IBM & ted |  ABN & TED ; 
 ABN <= IBN & ted |  ABO & TED ; 
 DPA <=  CBG & cdf & cfe  |  cbg & CDF & cfe  |  cbg & cdf & CFE  |  CBG & CDF & CFE  ;
 dpb <=  CBG & cdf & cfe  |  cbg & CDF & cfe  |  cbg & cdf & CFE  |  cbg & cdf & cfe  ;
 ABO <= IBO & ted |  ABP & TED ; 
 ABP <= IBP & ted |  ZZO & TED ; 
 DPC <=  CHD & cjc & clb  |  chd & CJC & clb  |  chd & cjc & CLB  |  CHD & CJC & CLB  ;
 dpd <=  CHD & cjc & clb  |  chd & CJC & clb  |  chd & cjc & CLB  |  chd & cjc & clb  ;
 DQA <=  CAH & ccg & cef  |  cah & CCG & cef  |  cah & ccg & CEF  |  CAH & CCG & CEF  ;
 dqb <=  CAH & ccg & cef  |  cah & CCG & cef  |  cah & ccg & CEF  |  cah & ccg & cef  ;
 FAA <= EAA ; 
 FBA <= EBA ; 
 FCA <= ECA ; 
 FDA <= EDA ; 
 DMC <=  CGC & cib & cka  |  cgc & CIB & cka  |  cgc & cib & CKA  |  CGC & CIB & CKA  ;
 dmd <=  CGC & cib & cka  |  cgc & CIB & cka  |  cgc & cib & CKA  |  cgc & cib & cka  ;
 ABA <= IBA & tec |  ABB & TEC ; 
 ABB <= IBB & tec |  ABC & TEC ; 
 ABC <= IBC & tec |  ABD & TEC ; 
 DNA <=  CBF & cde & cfd  |  cbf & CDE & cfd  |  cbf & cde & CFD  |  CBF & CDE & CFD  ;
 dnb <=  CBF & cde & cfd  |  cbf & CDE & cfd  |  cbf & cde & CFD  |  cbf & cde & cfd  ;
 ABD <= IBD & tec |  ABE & TEC ; 
 ABE <= IBE & tec |  ABF & TEC ; 
 ABF <= IBF & tec |  ABG & TEC ; 
 BAA <= IAA & tee |  BAA & TEE ; 
 BAB <= IAB & tee |  BAB & TEE ; 
 BAC <= IAC & tee |  BAC & TEE ; 
 OAA <= PFA & TFA |  ICA & tfa ; 
 OAB <= PFB & TFA |  ICB & tfa ; 
 OAC <= PFC & TFA |  ICC & tfa ; 
 BAD <= IAD & tee |  BAD & TEE ; 
 BAE <= IAE & tee |  BAE & TEE ; 
 BAF <= IAF & tee |  BAF & TEE ; 
 OAD <= PFD & TFA |  ICD & tfa ; 
 OAE <= PFE & TFA |  ICE & tfa ; 
 OAF <= PFF & TFA |  ICF & tfa ; 
 BAI <= IAI & tef |  BAI & TEF ; 
 BAJ <= IAJ & tef |  BAJ & TEF ; 
 BAK <= IAK & tef |  BAK & TEF ; 
 OAG <= PFG & TFA |  ICG & tfa ; 
 OAH <= PFH & TFA |  ICH & tfa ; 
 BAL <= IAL & tef |  BAL & TEF ; 
 BAM <= IAM & tef |  BAM & TEF ; 
 BAN <= IAN & tef |  BAN & TEF ; 
 OAI <= PFI & TFB |  ICI & tfb ; 
 OAJ <= PFJ & TFB |  ICJ & tfb ; 
 OAK <= PFK & TFB |  ICK & tfb ; 
 BBI <= IBI & teh |  BBI & TEH ; 
 BBJ <= IBJ & teh |  BBJ & TEH ; 
 BBK <= IBK & teh |  BBK & TEH ; 
 OAL <= PFL & TFB |  ICL & tfb ; 
 OAM <= PFM & TFB |  ICM & tfb ; 
 OAN <= PFN & TFB |  ICN & tfb ; 
 BBL <= IBL & teh |  BBL & TEH ; 
 BBM <= IBM & teh |  BBM & TEH ; 
 BBN <= IBN & teh |  BBN & TEH ; 
 OAO <= PFO & TFB |  ICO & tfb ; 
 OAP <= PFP & TFB |  ICP & tfb ; 
 KNB <= HNB ; 
 KJB <= HJB ; 
 PAQ <= NHE ; 
 DOE <= CMA ; 
 PAL <= NXB ; 
 FPC <= EPD ; 
 FGA <= EIA ; 
 OBA <= PGA & TFC |  IDA & tfc ; 
 OBB <= PGB & TFC |  IDB & tfc ; 
 OBC <= PGC & TFC |  IDC & tfc ; 
 OBE <= PGE & TFC |  IDE & tfc ; 
 OBF <= PGF & TFC |  IDF & tfc ; 
 OBG <= PGG & TFC |  IDG & tfc ; 
 OBD <= PGD & TFC |  IDD & tfc ; 
 DVG <= CTA ; 
 DRC <=  CHE & cjd & clc  |  che & CJD & clc  |  che & cjd & CLC  |  CHE & CJD & CLC  ;
 drd <=  CHE & cjd & clc  |  che & CJD & clc  |  che & cjd & CLC  |  che & cjd & clc  ;
 NAH <=  MHA  |  MGB  ; 
 MZD <=  LZD & lzf & lzb  |  lzd & LZF & lzb  |  lzd & lzf & LZB  |  LZD & LZF & LZB  ;
 mze <=  LZD & lzf & lzb  |  lzd & LZF & lzb  |  lzd & lzf & LZB  |  lzd & lzf & lzb  ;
 DSA <=  CAI & cch & ceg  |  cai & CCH & ceg  |  cai & cch & CEG  |  CAI & CCH & CEG  ;
 dsb <=  CAI & cch & ceg  |  cai & CCH & ceg  |  cai & cch & CEG  |  cai & cch & ceg  ;
 NEH <= MGB & MHA ; 
 DSC <=  CGF & cie & ckd  |  cgf & CIE & ckd  |  cgf & cie & CKD  |  CGF & CIE & CKD  ;
 dsd <=  CGF & cie & ckd  |  cgf & CIE & ckd  |  cgf & cie & CKD  |  cgf & cie & ckd  ;
 MKB <= LKA & LJB ; 
 NEI <= MHB & MIA ; 
 NEK <= MJB & MKA ; 
 DSE <=  CMC & cob & cqa  |  cmc & COB & cqa  |  cmc & cob & CQA  |  CMC & COB & CQA  ;
 dsf <=  CMC & cob & cqa  |  cmc & COB & cqa  |  cmc & cob & CQA  |  cmc & cob & cqa  ;
 FZI <=  EZM & ezo & ezq  |  ezm & EZO & ezq  |  ezm & ezo & EZQ  |  EZM & EZO & EZQ  ;
 fzj <=  EZM & ezo & ezq  |  ezm & EZO & ezq  |  ezm & ezo & EZQ  |  ezm & ezo & ezq  ;
 FZE <=  EZG & ezi & ezk  |  ezg & EZI & ezk  |  ezg & ezi & EZK  |  EZG & EZI & EZK  ;
 fzf <=  EZG & ezi & ezk  |  ezg & EZI & ezk  |  ezg & ezi & EZK  |  ezg & ezi & ezk  ;
 DTA <=  CBI & cdh & cfg  |  cbi & CDH & cfg  |  cbi & cdh & CFG  |  CBI & CDH & CFG  ;
 dtb <=  CBI & cdh & cfg  |  cbi & CDH & cfg  |  cbi & cdh & CFG  |  cbi & cdh & cfg  ;
 FZG <= EZB ; 
 FZH <= EZD ; 
 DTC <=  CHF & cje & cld  |  chf & CJE & cld  |  chf & cje & CLD  |  CHF & CJE & CLD  ;
 dtd <=  CHF & cje & cld  |  chf & CJE & cld  |  chf & cje & CLD  |  chf & cje & cld  ;
 BBD <= IBD & teg |  BBD & TEG ; 
 BBE <= IBE & teg |  BBE & TEG ; 
 BBF <= IBF & teg |  BBF & TEG ; 
 BBA <= IBA & teg |  BBA & TEG ; 
 BBB <= IBB & teg |  BBB & TEG ; 
 BBC <= IBC & teg |  BBC & TEG ; 
 DQC <=  CGE & cid & ckc  |  cge & CID & ckc  |  cge & cid & CKC  |  CGE & CID & CKC  ;
 dqd <=  CGE & cid & ckc  |  cge & CID & ckc  |  cge & cid & CKC  |  cge & cid & ckc  ;
 DRA <=  CBH & cdg & cff  |  cbh & CDG & cff  |  cbh & cdg & CFF  |  CBH & CDG & CFF  ;
 drb <=  CBH & cdg & cff  |  cbh & CDG & cff  |  cbh & cdg & CFF  |  cbh & cdg & cff  ;
 DUC <=  CGG & cif & cke  |  cgg & CIF & cke  |  cgg & cif & CKE  |  CGG & CIF & CKE  ;
 dud <=  CGG & cif & cke  |  cgg & CIF & cke  |  cgg & cif & CKE  |  cgg & cif & cke  ;
 DUE <=  CMD & coc & cqb  |  cmd & COC & cqb  |  cmd & coc & CQB  |  CMD & COC & CQB  ;
 duf <=  CMD & coc & cqb  |  cmd & COC & cqb  |  cmd & coc & CQB  |  cmd & coc & cqb  ;
 FEA <= EEA ; 
 NEL <= MKB & MLA ; 
 QYS <= CYB & DAA ; 
 DVA <=  CBJ & cdi & cfh  |  cbj & CDI & cfh  |  cbj & cdi & CFH  |  CBJ & CDI & CFH  ;
 dvb <=  CBJ & cdi & cfh  |  cbj & CDI & cfh  |  cbj & cdi & CFH  |  cbj & cdi & cfh  ;
 FRC <= ERE ; 
 NEM <= MLB & MMA ; 
 HNA <= GNA ; 
 HNB <= GMB ; 
 HOA <= GOA ; 
 FWC <= EWE ; 
 DVC <=  CHG & cjf & cle  |  chg & CJF & cle  |  chg & cjf & CLE  |  CHG & CJF & CLE  ;
 dvd <=  CHG & cjf & cle  |  chg & CJF & cle  |  chg & cjf & CLE  |  chg & cjf & cle  ;
 DVE <=  CND & cpc & crb  |  cnd & CPC & crb  |  cnd & cpc & CRB  |  CND & CPC & CRB  ;
 dvf <=  CND & cpc & crb  |  cnd & CPC & crb  |  cnd & cpc & CRB  |  cnd & cpc & crb  ;
 KXA <=  HXA & hxc & hwb  |  hxa & HXC & hwb  |  hxa & hxc & HWB  |  HXA & HXC & HWB  ;
 kxb <=  HXA & hxc & hwb  |  hxa & HXC & hwb  |  hxa & hxc & HWB  |  hxa & hxc & hwb  ;
 DWA <=  CAK & ccj & cei  |  cak & CCJ & cei  |  cak & ccj & CEI  |  CAK & CCJ & CEI  ;
 dwb <=  CAK & ccj & cei  |  cak & CCJ & cei  |  cak & ccj & CEI  |  cak & ccj & cei  ;
 FZM <=  EZS & ezu & ezw  |  ezs & EZU & ezw  |  ezs & ezu & EZW  |  EZS & EZU & EZW  ;
 fzn <=  EZS & ezu & ezw  |  ezs & EZU & ezw  |  ezs & ezu & EZW  |  ezs & ezu & ezw  ;
 DTE <=  CNC & cpb & cra  |  cnc & CPB & cra  |  cnc & cpb & CRA  |  CNC & CPB & CRA  ;
 dtf <=  CNC & cpb & cra  |  cnc & CPB & cra  |  cnc & cpb & CRA  |  cnc & cpb & cra  ;
 HZG <=  GZG & gzf & gzd  |  gzg & GZF & gzd  |  gzg & gzf & GZD  |  GZG & GZF & GZD  ;
 hzh <=  GZG & gzf & gzd  |  gzg & GZF & gzd  |  gzg & gzf & GZD  |  gzg & gzf & gzd  ;
 DUA <=  CAJ & cci & ceh  |  caj & CCI & ceh  |  caj & cci & CEH  |  CAJ & CCI & CEH  ;
 dub <=  CAJ & cci & ceh  |  caj & CCI & ceh  |  caj & cci & CEH  |  caj & cci & ceh  ;
 HXC <= GWD ; 
 FOC <= EOD ; 
 FCB <= ECB ; 
 FRD <= EQD ; 
 MBB <= LBB ; 
 OBH <= PGH & TFC |  IDH & tfc ; 
 OBI <= PGI & TFD |  IDI & tfd ; 
 OBJ <= PGJ & TFD |  IDJ & tfd ; 
 OBK <= PGK & TFD |  IDK & tfd ; 
 FYQ <=  EXT & exh & exj  |  ext & EXH & exj  |  ext & exh & EXJ  |  EXT & EXH & EXJ  ;
 fyr <=  EXT & exh & exj  |  ext & EXH & exj  |  ext & exh & EXJ  |  ext & exh & exj  ;
 MJA <=  LJA & lib & lid  |  lja & LIB & lid  |  lja & lib & LID  |  LJA & LIB & LID  ;
 mjb <=  LJA & lib & lid  |  lja & LIB & lid  |  lja & lib & LID  |  lja & lib & lid  ;
 OBL <= PGL & TFD |  IDL & tfd ; 
 OBM <= PGM & TFD |  IDM & tfd ; 
 OBN <= PGN & TFD |  IDN & tfd ; 
 FQC <= ZZO ; 
 HZO <= ZZO ; 
 FWD <= EVD ; 
 OBO <= PGO & TFD |  IDO & tfd ; 
 OBP <= PGP & TFD |  IDP & tfd ; 
 MMA <= LMA & llb |  lma & LLB ; 
 NFB <= MSA & MRB ; 
 FDB <= EDB ; 
 FZV <= EZX ; 
 FYI <= EYR ; 
 KBA <= HBA ; 
 KCA <= HCA ; 
 KDA <= HDA ; 
 NEN <= MMB & MNA ; 
 AAQ <= TEB & AAA ; 
 FOA <=  EOA & enb & eoc  |  eoa & ENB & eoc  |  eoa & enb & EOC  |  EOA & ENB & EOC  ;
 fob <=  EOA & enb & eoc  |  eoa & ENB & eoc  |  eoa & enb & EOC  |  eoa & enb & eoc  ;
 FPA <=  EPA & epc & eob  |  epa & EPC & eob  |  epa & epc & EOB  |  EPA & EPC & EOB  ;
 fpb <=  EPA & epc & eob  |  epa & EPC & eob  |  epa & epc & EOB  |  epa & epc & eob  ;
 DWC <=  CGH & cig & ckf  |  cgh & CIG & ckf  |  cgh & cig & CKF  |  CGH & CIG & CKF  ;
 dwd <=  CGH & cig & ckf  |  cgh & CIG & ckf  |  cgh & cig & CKF  |  cgh & cig & ckf  ;
 FQA <=  EQA & eqc & epb  |  eqa & EQC & epb  |  eqa & eqc & EPB  |  EQA & EQC & EPB  ;
 fqb <=  EQA & eqc & epb  |  eqa & EQC & epb  |  eqa & eqc & EPB  |  eqa & eqc & epb  ;
 FRA <=  ERA & erc & eqb  |  era & ERC & eqb  |  era & erc & EQB  |  ERA & ERC & EQB  ;
 frb <=  ERA & erc & eqb  |  era & ERC & eqb  |  era & erc & EQB  |  era & erc & eqb  ;
 DWE <=  CME & cod & cqc  |  cme & COD & cqc  |  cme & cod & CQC  |  CME & COD & CQC  ;
 dwf <=  CME & cod & cqc  |  cme & COD & cqc  |  cme & cod & CQC  |  cme & cod & cqc  ;
 FYJ <=  EXG & exi & exk  |  exg & EXI & exk  |  exg & exi & EXK  |  EXG & EXI & EXK  ;
 fyk <=  EXG & exi & exk  |  exg & EXI & exk  |  exg & exi & EXK  |  exg & exi & exk  ;
 FSA <=  ESA & esc & erb  |  esa & ESC & erb  |  esa & esc & ERB  |  ESA & ESC & ERB  ;
 fsb <=  ESA & esc & erb  |  esa & ESC & erb  |  esa & esc & ERB  |  esa & esc & erb  ;
 FTA <=  ETA & etc & esb  |  eta & ETC & esb  |  eta & etc & ESB  |  ETA & ETC & ESB  ;
 ftb <=  ETA & etc & esb  |  eta & ETC & esb  |  eta & etc & ESB  |  eta & etc & esb  ;
 DXA <=  CBK & cdj & cfi  |  cbk & CDJ & cfi  |  cbk & cdj & CFI  |  CBK & CDJ & CFI  ;
 dxb <=  CBK & cdj & cfi  |  cbk & CDJ & cfi  |  cbk & cdj & CFI  |  cbk & cdj & cfi  ;
 QZI <= CZB & dba |  czb & DBA ; 
 FUA <=  EUA & euc & etb  |  eua & EUC & etb  |  eua & euc & ETB  |  EUA & EUC & ETB  ;
 fub <=  EUA & euc & etb  |  eua & EUC & etb  |  eua & euc & ETB  |  eua & euc & etb  ;
 FVA <=  EVA & evc & eub  |  eva & EVC & eub  |  eva & evc & EUB  |  EVA & EVC & EUB  ;
 fvb <=  EVA & evc & eub  |  eva & EVC & eub  |  eva & evc & EUB  |  eva & evc & eub  ;
 DXC <=  CHH & cjg & clf  |  chh & CJG & clf  |  chh & cjg & CLF  |  CHH & CJG & CLF  ;
 dxd <=  CHH & cjg & clf  |  chh & CJG & clf  |  chh & cjg & CLF  |  chh & cjg & clf  ;
 MKA <= LKA & ljb |  lka & LJB ; 
 FWA <=  EWA & ewc & evb  |  ewa & EWC & evb  |  ewa & ewc & EVB  |  EWA & EWC & EVB  ;
 fwb <=  EWA & ewc & evb  |  ewa & EWC & evb  |  ewa & ewc & EVB  |  ewa & ewc & evb  ;
 HZY <=  GYF & gyh & gzy  |  gyf & GYH & gzy  |  gyf & gyh & GZY  |  GYF & GYH & GZY  ;
 hzz <=  GYF & gyh & gzy  |  gyf & GYH & gzy  |  gyf & gyh & GZY  |  gyf & gyh & gzy  ;
 DXE <=  CNE & cpd & crc  |  cne & CPD & crc  |  cne & cpd & CRC  |  CNE & CPD & CRC  ;
 dxf <=  CNE & cpd & crc  |  cne & CPD & crc  |  cne & cpd & CRC  |  cne & cpd & crc  ;
 HRA <=  GRA & grc & gqb  |  gra & GRC & gqb  |  gra & grc & GQB  |  GRA & GRC & GQB  ;
 hrb <=  GRA & grc & gqb  |  gra & GRC & gqb  |  gra & grc & GQB  |  gra & grc & gqb  ;
 FXA <=  EXA & exc & ewb  |  exa & EXC & ewb  |  exa & exc & EWB  |  EXA & EXC & EWB  ;
 fxb <=  EXA & exc & ewb  |  exa & EXC & ewb  |  exa & exc & EWB  |  exa & exc & ewb  ;
 FXC <=  EXE & exf & ewd  |  exe & EXF & ewd  |  exe & exf & EWD  |  EXE & EXF & EWD  ;
 fxd <=  EXE & exf & ewd  |  exe & EXF & ewd  |  exe & exf & EWD  |  exe & exf & ewd  ;
 HZQ <=  GZQ & gzs & gzn  |  gzq & GZS & gzn  |  gzq & gzs & GZN  |  GZQ & GZS & GZN  ;
 hzr <=  GZQ & gzs & gzn  |  gzq & GZS & gzn  |  gzq & gzs & GZN  |  gzq & gzs & gzn  ;
 FIA <=  EKA & ekc & ejb  |  eka & EKC & ejb  |  eka & ekc & EJB  |  EKA & EKC & EJB  ;
 fib <=  EKA & ekc & ejb  |  eka & EKC & ejb  |  eka & ekc & EJB  |  eka & ekc & ejb  ;
 KAA <= HAA ; 
 FJA <=  ELA & elc & ekb  |  ela & ELC & ekb  |  ela & elc & EKB  |  ELA & ELC & EKB  ;
 fjb <=  ELA & elc & ekb  |  ela & ELC & ekb  |  ela & elc & EKB  |  ela & elc & ekb  ;
 HZW <=  GZX & gzz & gzu  |  gzx & GZZ & gzu  |  gzx & gzz & GZU  |  GZX & GZZ & GZU  ;
 hzx <=  GZX & gzz & gzu  |  gzx & GZZ & gzu  |  gzx & gzz & GZU  |  gzx & gzz & gzu  ;
 KZM <=  HZM & hzo & hzj  |  hzm & HZO & hzj  |  hzm & hzo & HZJ  |  HZM & HZO & HZJ  ;
 kzn <=  HZM & hzo & hzj  |  hzm & HZO & hzj  |  hzm & hzo & HZJ  |  hzm & hzo & hzj  ;
 FMA <= EMA ; 
 FMB <= ELB ; 
 KZT <= JZT ; 
 KZY <= JZY ; 
 FNA <=  ENA & enc & emb  |  ena & ENC & emb  |  ena & enc & EMB  |  ENA & ENC & EMB  ;
 fnb <=  ENA & enc & emb  |  ena & ENC & emb  |  ena & enc & EMB  |  ena & enc & emb  ;
 DYE <=  CMF & coe & cqd  |  cmf & COE & cqd  |  cmf & coe & CQD  |  CMF & COE & CQD  ;
 dyf <=  CMF & coe & cqd  |  cmf & COE & cqd  |  cmf & coe & CQD  |  cmf & coe & cqd  ;
 oia <= ifa ; 
 oka <= ifa ; 
 oma <= ifa ; 
 ooa <= ifa ; 
 DYG <=  CSC & cub & cwa  |  csc & CUB & cwa  |  csc & cub & CWA  |  CSC & CUB & CWA  ;
 dyh <=  CSC & cub & cwa  |  csc & CUB & cwa  |  csc & cub & CWA  |  csc & cub & cwa  ;
 NEP <= MOB & MQA ; 
 DZA <=  CBL & cdk & cfj  |  cbl & CDK & cfj  |  cbl & cdk & CFJ  |  CBL & CDK & CFJ  ;
 dzb <=  CBL & cdk & cfj  |  cbl & CDK & cfj  |  cbl & cdk & CFJ  |  cbl & cdk & cfj  ;
 DZC <=  CHI & cjh & clg  |  chi & CJH & clg  |  chi & cjh & CLG  |  CHI & CJH & CLG  ;
 dzd <=  CHI & cjh & clg  |  chi & CJH & clg  |  chi & cjh & CLG  |  chi & cjh & clg  ;
 DZE <=  CNF & cpe & crd  |  cnf & CPE & crd  |  cnf & cpe & CRD  |  CNF & CPE & CRD  ;
 dzf <=  CNF & cpe & crd  |  cnf & CPE & crd  |  cnf & cpe & CRD  |  cnf & cpe & crd  ;
 DZG <=  CTC & cvb & cxa  |  ctc & CVB & cxa  |  ctc & cvb & CXA  |  CTC & CVB & CXA  ;
 dzh <=  CTC & cvb & cxa  |  ctc & CVB & cxa  |  ctc & cvb & CXA  |  ctc & cvb & cxa  ;
 MLA <= LLA & lkb |  lla & LKB ; 
 DYA <=  CAL & cck & cej  |  cal & CCK & cej  |  cal & cck & CEJ  |  CAL & CCK & CEJ  ;
 dyb <=  CAL & cck & cej  |  cal & CCK & cej  |  cal & cck & CEJ  |  cal & cck & cej  ;
 DYC <=  CGI & cih & ckg  |  cgi & CIH & ckg  |  cgi & cih & CKG  |  CGI & CIH & CKG  ;
 dyd <=  CGI & cih & ckg  |  cgi & CIH & ckg  |  cgi & cih & CKG  |  cgi & cih & ckg  ;
 oih <= iga ; 
 okh <= iga ; 
 omh <= iga ; 
 ooh <= iga ; 
 KEA <= HEA ; 
 HFA <= FFA ; 
 HFB <= ZZO ; 
 MOA <=  LOA & loc & lnb  |  loa & LOC & lnb  |  loa & loc & LNB  |  LOA & LOC & LNB  ;
 mob <=  LOA & loc & lnb  |  loa & LOC & lnb  |  loa & loc & LNB  |  loa & loc & lnb  ;
 KFA <= HFA ; 
 KGA <= HGA ; 
 FZC <=  EZF & eyb & eyd  |  ezf & EYB & eyd  |  ezf & eyb & EYD  |  EZF & EYB & EYD  ;
 fzd <=  EZF & eyb & eyd  |  ezf & EYB & eyd  |  ezf & eyb & EYD  |  ezf & eyb & eyd  ;
 KIA <= HIA ; 
 FXE <= EWF ; 
 KJA <= HJA ; 
 NFC <= MSB & MTA ; 
 KMA <= HMA ; 
 KHA <=  HHA & hhb & hgb  |  hha & HHB & hgb  |  hha & hhb & HGB  |  HHA & HHB & HGB  ;
 khb <=  HHA & hhb & hgb  |  hha & HHB & hgb  |  hha & hhb & HGB  |  hha & hhb & hgb  ;
 KNA <= HNA ; 
 KOA <= HOA ; 
 NAQ <= MQB & MRA ; 
 KPA <= HPA ; 
 KPB <= HPB ; 
 KQA <= HQA ; 
 FSD <= ESD ; 
 KQB <= HQB ; 
 KRA <= HRA ; 
 KSA <= HSA ; 
 KSB <= HRB ; 
 MNA <= LNA & lmb |  lna & LMB ; 
 NFG <= MWB & MXA ; 
 NFH <= MXB & MYA ; 
 NFI <= MYB & MZA ; 
 KZW <= HZW & hzu |  hzw & HZU ; 
 NFL <= MZJ & MZL ; 
 pak <=  nxi  |  nxj  |  nxk  |  nxl  ; 
 oib <= ifb ; 
 okb <= ifb ; 
 omb <= ifb ; 
 oob <= ifb ; 
 FZK <=  EZH & ezj & ezl  |  ezh & EZJ & ezl  |  ezh & ezj & EZL  |  EZH & EZJ & EZL  ;
 fzl <=  EZH & ezj & ezl  |  ezh & EZJ & ezl  |  ezh & ezj & EZL  |  ezh & ezj & ezl  ;
 MQB <= LQA & LOB ; 
 FZO <=  EZR & ezn & ezp  |  ezr & EZN & ezp  |  ezr & ezn & EZP  |  EZR & EZN & EZP  ;
 fzp <=  EZR & ezn & ezp  |  ezr & EZN & ezp  |  ezr & ezn & EZP  |  ezr & ezn & ezp  ;
 DLC <= CHB ; 
 DLD <= CJA ; 
 DQE <= CMB ; 
 DRE <= CNB ; 
 DQF <= COA ; 
 DRF <= CPA ; 
 FZY <=  EYG & eyi & eyk  |  eyg & EYI & eyk  |  eyg & eyi & EYK  |  EYG & EYI & EYK  ;
 fzz <=  EYG & eyi & eyk  |  eyg & EYI & eyk  |  eyg & eyi & EYK  |  eyg & eyi & eyk  ;
 MSA <=  LSA & lsc & lrb  |  lsa & LSC & lrb  |  lsa & lsc & LRB  |  LSA & LSC & LRB  ;
 msb <=  LSA & lsc & lrb  |  lsa & LSC & lrb  |  lsa & lsc & LRB  |  lsa & lsc & lrb  ;
 FHA <= EJA ; 
 HZK <= ZZO ; 
 HZV <= GZW ; 
 oii <= igb ; 
 oki <= igb ; 
 omi <= igb ; 
 ooi <= igb ; 
 FYA <=  EYA & eyc & exb  |  eya & EYC & exb  |  eya & eyc & EXB  |  EYA & EYC & EXB  ;
 fyb <=  EYA & eyc & exb  |  eya & EYC & exb  |  eya & eyc & EXB  |  eya & eyc & exb  ;
 NFF <= MVB & MWA ; 
 DZM <=  CMG & cof & cqe  |  cmg & COF & cqe  |  cmg & cof & CQE  |  CMG & COF & CQE  ;
 dzn <=  CMG & cof & cqe  |  cmg & COF & cqe  |  cmg & cof & CQE  |  cmg & cof & cqe  ;
 oij <= igc ; 
 okj <= igc ; 
 omj <= igc ; 
 ooj <= igc ; 
 DZO <=  CSD & cuc & cwb  |  csd & CUC & cwb  |  csd & cuc & CWB  |  CSD & CUC & CWB  ;
 dzp <=  CSD & cuc & cwb  |  csd & CUC & cwb  |  csd & cuc & CWB  |  csd & cuc & cwb  ;
 KZX <= HZU & HZW ; 
 QYA <=  CBM & cdl & cfk  |  cbm & CDL & cfk  |  cbm & cdl & CFK  |  CBM & CDL & CFK  ;
 qyb <=  CBM & cdl & cfk  |  cbm & CDL & cfk  |  cbm & cdl & CFK  |  cbm & cdl & cfk  ;
 HYD <= GYI & gye |  gyi & GYE ; 
 QYC <=  CHJ & cji & clh  |  chj & CJI & clh  |  chj & cji & CLH  |  CHJ & CJI & CLH  ;
 qyd <=  CHJ & cji & clh  |  chj & CJI & clh  |  chj & cji & CLH  |  chj & cji & clh  ;
 oic <= ifc ; 
 MTA <=  LTA & ltc & lsb  |  lta & LTC & lsb  |  lta & ltc & LSB  |  LTA & LTC & LSB  ;
 mtb <=  LTA & ltc & lsb  |  lta & LTC & lsb  |  lta & ltc & LSB  |  lta & ltc & lsb  ;
 okc <= ifc ; 
 QYE <=  CNG & cpf & cre  |  cng & CPF & cre  |  cng & cpf & CRE  |  CNG & CPF & CRE  ;
 qyf <=  CNG & cpf & cre  |  cng & CPF & cre  |  cng & cpf & CRE  |  cng & cpf & cre  ;
 omc <= ifc ; 
 QVF <= DBC ; 
 QYG <=  CTD & cvc & cxb  |  ctd & CVC & cxb  |  ctd & cvc & CXB  |  CTD & CVC & CXB  ;
 qyh <=  CTD & cvc & cxb  |  ctd & CVC & cxb  |  ctd & cvc & CXB  |  ctd & cvc & cxb  ;
 ooc <= ifc ; 
 MFA <= LFA & leb |  lfa & LEB ; 
 MWA <=  LWA & lwc & lvb  |  lwa & LWC & lvb  |  lwa & lwc & LVB  |  LWA & LWC & LVB  ;
 mwb <=  LWA & lwc & lvb  |  lwa & LWC & lvb  |  lwa & lwc & LVB  |  lwa & lwc & lvb  ;
 MXA <=  LXA & lxc & lwb  |  lxa & LXC & lwb  |  lxa & lxc & LWB  |  LXA & LXC & LWB  ;
 mxb <=  LXA & lxc & lwb  |  lxa & LXC & lwb  |  lxa & lxc & LWB  |  lxa & lxc & lwb  ;
 DZI <=  CAM & ccl & cek  |  cam & CCL & cek  |  cam & ccl & CEK  |  CAM & CCL & CEK  ;
 dzj <=  CAM & ccl & cek  |  cam & CCL & cek  |  cam & ccl & CEK  |  cam & ccl & cek  ;
 HTA <= GTA & gsb |  gta & GSB ; 
 DZK <=  CGJ & cii & ckh  |  cgj & CII & ckh  |  cgj & cii & CKH  |  CGJ & CII & CKH  ;
 dzl <=  CGJ & cii & ckh  |  cgj & CII & ckh  |  cgj & cii & CKH  |  cgj & cii & ckh  ;
 MRB <= LQB & LRA ; 
 KUA <= HUA & htb |  hua & HTB ; 
 KWA <= HWA & hvb |  hwa & HVB ; 
 oik <= igd ; 
 okk <= igd ; 
 omk <= igd ; 
 ook <= igd ; 
 PAB <=  NGE  ; 
 oie <= ife ; 
 oke <= ife ; 
 ome <= ife ; 
 ooe <= ife ; 
 PAD <=  NGE & NXB & NXC  |  NHE & NXC  |  NIE  ; 
 PAE <=  NGE & NXB & NXC & NXD  |  NHE & NXC & NXD  |  NIE & NXD  |  NJE  ; 
 KZI <=  HZH & hzi & hzk  |  hzh & HZI & hzk  |  hzh & hzi & HZK  |  HZH & HZI & HZK  ;
 kzj <=  HZH & hzi & hzk  |  hzh & HZI & hzk  |  hzh & hzi & HZK  |  hzh & hzi & hzk  ;
 HAA <= FAA ; 
 HBA <= FBA ; 
 HCA <= FCA ; 
 HDA <= FDA ; 
 HZC <=  GZC & gze & gzb  |  gzc & GZE & gzb  |  gzc & gze & GZB  |  GZC & GZE & GZB  ;
 hzd <=  GZC & gze & gzb  |  gzc & GZE & gzb  |  gzc & gze & GZB  |  gzc & gze & gzb  ;
 PFB <= PBB ; 
 PFC <= PBC ; 
 PFD <= PBD ; 
 PFA <= PBA ; 
 MEA <= LEA & ldb |  lea & LDB ; 
 oid <= ifd ; 
 okd <= ifd ; 
 omd <= ifd ; 
 ood <= ifd ; 
 QZJ <= DBA & DBA ; 
 oif <= iiff ; 
 okf <= iiff ; 
 omf <= iiff ; 
 oof <= iiff ; 
 FYC <= EYE & exd |  eye & EXD ; 
 PDF <= RAF & npb |  raf & NPB ; 
 PDG <= RAG & npc |  rag & NPC ; 
 PDH <= RAH & npd |  rah & NPD ; 
 FYE <=  EYS & eyu & eyw  |  eys & EYU & eyw  |  eys & eyu & EYW  |  EYS & EYU & EYW  ;
 fyf <=  EYS & eyu & eyw  |  eys & EYU & eyw  |  eys & eyu & EYW  |  eys & eyu & eyw  ;
 PDK <= RAK & nqc |  rak & NQC ; 
 PDL <= RAL & nqd |  ral & NQD ; 
 PDJ <= RAJ & nqb |  raj & NQB ; 
 PDN <= RAN & nrb |  ran & NRB ; 
 FYG <=  EYY & eyn & eyp  |  eyy & EYN & eyp  |  eyy & eyn & EYP  |  EYY & EYN & EYP  ;
 fyh <=  EYY & eyn & eyp  |  eyy & EYN & eyp  |  eyy & eyn & EYP  |  eyy & eyn & eyp  ;
 PDP <= RAP & nrd |  rap & NRD ; 
 PDO <= RAO & nrc |  rao & NRC ; 
 FYL <=  EXM & eyt & eyv  |  exm & EYT & eyv  |  exm & eyt & EYV  |  EXM & EYT & EYV  ;
 fym <=  EXM & eyt & eyv  |  exm & EYT & eyv  |  exm & eyt & EYV  |  exm & eyt & eyv  ;
 oil <= ige ; 
 okl <= ige ; 
 oml <= ige ; 
 ool <= ige ; 
 FSC <= ERD ; 
 PEB <= RBB & nsb |  rbb & NSB ; 
 MFB <= LEB & LFA ; 
 PEC <= RBC & nsc |  rbc & NSC ; 
 HUA <=  GUA & gtb & guc  |  gua & GTB & guc  |  gua & gtb & GUC  |  GUA & GTB & GUC  ;
 hub <=  GUA & gtb & guc  |  gua & GTB & guc  |  gua & gtb & GUC  |  gua & gtb & guc  ;
 PED <= RBD & nsd |  rbd & NSD ; 
 MQA <= LQA & lob |  lqa & LOB ; 
 PAC <=  NGE & NXB  |  NHE  ; 
 KTA <= HTA & hsb |  hta & HSB ; 
 KZQ <= HZQ & hzn |  hzq & HZN ; 
 QYN <=  CMH & cog & cqf  |  cmh & COG & cqf  |  cmh & cog & CQF  |  CMH & COG & CQF  ;
 qyo <=  CMH & cog & cqf  |  cmh & COG & cqf  |  cmh & cog & CQF  |  cmh & cog & cqf  ;
 PEJ <= RBJ & nub |  rbj & NUB ; 
 MLB <= LLA & LKB ; 
 QYP <=  CSE & cud & cwc  |  cse & CUD & cwc  |  cse & cud & CWC  |  CSE & CUD & CWC  ;
 qyq <=  CSE & cud & cwc  |  cse & CUD & cwc  |  cse & cud & CWC  |  cse & cud & cwc  ;
 PEK <= RBK & nuc |  rbk & NUC ; 
 MRA <= LRA & lqb |  lra & LQB ; 
 QZA <=  CBN & cdm & cfl  |  cbn & CDM & cfl  |  cbn & cdm & CFL  |  CBN & CDM & CFL  ;
 qzb <=  CBN & cdm & cfl  |  cbn & CDM & cfl  |  cbn & cdm & CFL  |  cbn & cdm & cfl  ;
 PEP <= RBP & nvd |  rbp & NVD ; 
 QZC <=  CHK & cjj & cli  |  chk & CJJ & cli  |  chk & cjj & CLI  |  CHK & CJJ & CLI  ;
 qzd <=  CHK & cjj & cli  |  chk & CJJ & cli  |  chk & cjj & CLI  |  chk & cjj & cli  ;
 PEL <= RBL & nud |  rbl & NUD ; 
 NFE <= MUB & MVA ; 
 QZE <=  CNH & cpg & crf  |  cnh & CPG & crf  |  cnh & cpg & CRF  |  CNH & CPG & CRF  ;
 qzf <=  CNH & cpg & crf  |  cnh & CPG & crf  |  cnh & cpg & CRF  |  cnh & cpg & crf  ;
 oim <= igf ; 
 okm <= igf ; 
 omm <= igf ; 
 oom <= igf ; 
 KZR <= HZN & HZQ ; 
 QZG <=  CTE & cvd & cxc  |  cte & CVD & cxc  |  cte & cvd & CXC  |  CTE & CVD & CXC  ;
 qzh <=  CTE & cvd & cxc  |  cte & CVD & cxc  |  cte & cvd & CXC  |  cte & cvd & cxc  ;
 NFK <= MZE & MZI ; 
 KVA <= HVA & hub |  hva & HUB ; 
 QYJ <=  CAN & ccm & cel  |  can & CCM & cel  |  can & ccm & CEL  |  CAN & CCM & CEL  ;
 qyk <=  CAN & ccm & cel  |  can & CCM & cel  |  can & ccm & CEL  |  can & ccm & cel  ;
 PEG <= RBG & ntc |  rbg & NTC ; 
 MUA <=  LUA & ltb & luc  |  lua & LTB & luc  |  lua & ltb & LUC  |  LUA & LTB & LUC  ;
 mub <=  LUA & ltb & luc  |  lua & LTB & luc  |  lua & ltb & LUC  |  lua & ltb & luc  ;
 QYL <=  CGK & cij & cki  |  cgk & CIJ & cki  |  cgk & cij & CKI  |  CGK & CIJ & CKI  ;
 qym <=  CGK & cij & cki  |  cgk & CIJ & cki  |  cgk & cij & CKI  |  cgk & cij & cki  ;
 PEH <= RBH & ntd |  rbh & NTD ; 
 NAA <= MAA ; 
 NAC <= MCA ; 
 QVG <= DDB ; 
 ohf <= ief ; 
 OJA <= IFA ; 
 OLA <= IFA ; 
 ONA <= IFA ; 
 OPA <= IFA ; 
 NAD <= MDA ; 
 NAE <=  MEA  |  MDB  ; 
 FUC <= ETD ; 
 OJB <= IFB ; 
 OLB <= IFB ; 
 ONB <= IFB ; 
 OPB <= IFB ; 
 NAG <=  MGA  |  MFB  ; 
 NAB <= MBA & mbb |  mba & MBB ; 
 NAJ <=  MJA  |  MIB  ; 
 NAI <=  MIA  |  MHB  ; 
 NAK <=  MKA  |  MJB  ; 
 NAL <=  MLA  |  MKB  ; 
 NAM <=  MMA  |  MLB  ; 
 NAN <=  MNA  |  MMB  ; 
 NAO <=  MOA  |  MNB  ; 
 NAP <=  MQA  |  MOB  ; 
 NBJ <=  MZD  |  MZB  ; 
 NBK <=  MZI  |  MZE  ; 
 NBM <=  MZO  |  MZM  ; 
 NBL <=  MZL  |  MZJ  ; 
 NBN <=  MZR  |  MZP  ; 
 NBO <=  MZU  |  MZS  ; 
 NBD <=  MUA  |  MTB  ; 
 FYO <=  EXN & exp & exr  |  exn & EXP & exr  |  exn & exp & EXR  |  EXN & EXP & EXR  ;
 fyp <=  EXN & exp & exr  |  exn & EXP & exr  |  exn & exp & EXR  |  exn & exp & exr  ;
 KZC <= HZC & hzb |  hzc & HZB ; 
 NBF <=  MWA  |  MVB  ; 
 NBH <=  MYA  |  MXB  ; 
 NFN <= MZP & MZR ; 
 KWB <= HWA & HVB ; 
 KYB <= HXB & HYA ; 
 NBI <=  MZA  |  MYB  ; 
 NFD <= MTB & MUA ; 
 KVB <= HUB & HVA ; 
 NBA <=  MRA  |  MQB  ; 
 NFO <= MZS & MZU ; 
 NFJ <= MZB & MZD ; 
 KZD <= HZB & HZC ; 
 QZO <=  CMI & coh & cqg  |  cmi & COH & cqg  |  cmi & coh & CQG  |  CMI & COH & CQG  ;
 qzp <=  CMI & coh & cqg  |  cmi & COH & cqg  |  cmi & coh & CQG  |  cmi & coh & cqg  ;
 FZR <=  EYF & eyh & eyj  |  eyf & EYH & eyj  |  eyf & eyh & EYJ  |  EYF & EYH & EYJ  ;
 fzs <=  EYF & eyh & eyj  |  eyf & EYH & eyj  |  eyf & eyh & EYJ  |  eyf & eyh & eyj  ;
 QZQ <=  CSF & cue & cwd  |  csf & CUE & cwd  |  csf & cue & CWD  |  CSF & CUE & CWD  ;
 qzr <=  CSF & cue & cwd  |  csf & CUE & cwd  |  csf & cue & CWD  |  csf & cue & cwd  ;
 OJC <= IFC ; 
 OLC <= IFC ; 
 ONC <= IFC ; 
 OPC <= IFC ; 
 QZS <=  CYC & dab & dca  |  cyc & DAB & dca  |  cyc & dab & DCA  |  CYC & DAB & DCA  ;
 qzt <=  CYC & dab & dca  |  cyc & DAB & dca  |  cyc & dab & DCA  |  cyc & dab & dca  ;
 QXA <=  CBO & cdn & cfm  |  cbo & CDN & cfm  |  cbo & cdn & CFM  |  CBO & CDN & CFM  ;
 qxb <=  CBO & cdn & cfm  |  cbo & CDN & cfm  |  cbo & cdn & CFM  |  cbo & cdn & cfm  ;
 QXC <=  CHL & cjk & clj  |  chl & CJK & clj  |  chl & cjk & CLJ  |  CHL & CJK & CLJ  ;
 qxd <=  CHL & cjk & clj  |  chl & CJK & clj  |  chl & cjk & CLJ  |  chl & cjk & clj  ;
 QXE <=  CNI & cph & crg  |  cni & CPH & crg  |  cni & cph & CRG  |  CNI & CPH & CRG  ;
 qxf <=  CNI & cph & crg  |  cni & CPH & crg  |  cni & cph & CRG  |  cni & cph & crg  ;
 QZK <=  CAO & ccn & cem  |  cao & CCN & cem  |  cao & ccn & CEM  |  CAO & CCN & CEM  ;
 qzl <=  CAO & ccn & cem  |  cao & CCN & cem  |  cao & ccn & CEM  |  cao & ccn & cem  ;
 NBP <=  MZX  |  MZV  ; 
 NBE <=  MVA  |  MUB  ; 
 QZM <=  CGL & cik & ckj  |  cgl & CIK & ckj  |  cgl & cik & CKJ  |  CGL & CIK & CKJ  ;
 qzn <=  CGL & cik & ckj  |  cgl & CIK & ckj  |  cgl & cik & CKJ  |  cgl & cik & ckj  ;
 NBG <=  MXA  |  MWB  ; 
 MIA <=  LIA & lhb & lic  |  lia & LHB & lic  |  lia & lhb & LIC  |  LIA & LHB & LIC  ;
 mib <=  LIA & lhb & lic  |  lia & LHB & lic  |  lia & lhb & LIC  |  lia & lhb & lic  ;
 OJH <= IGA ; 
 OLH <= IGA ; 
 ONH <= IGA ; 
 OPH <= IGA ; 
 HXA <=  GXA & gxc & gwb  |  gxa & GXC & gwb  |  gxa & gxc & GWB  |  GXA & GXC & GWB  ;
 hxb <=  GXA & gxc & gwb  |  gxa & GXC & gwb  |  gxa & gxc & GWB  |  gxa & gxc & gwb  ;
 NFM <= MZM & MZO ; 
 MZU <=  LZU & lzw & lzs  |  lzu & LZW & lzs  |  lzu & lzw & LZS  |  LZU & LZW & LZS  ;
 mzv <=  LZU & lzw & lzs  |  lzu & LZW & lzs  |  lzu & lzw & LZS  |  lzu & lzw & lzs  ;
 MZA <=  LZA & lzc & lyb  |  lza & LZC & lyb  |  lza & lzc & LYB  |  LZA & LZC & LYB  ;
 mzb <=  LZA & lzc & lyb  |  lza & LZC & lyb  |  lza & lzc & LYB  |  lza & lzc & lyb  ;
 MZL <=  LZL & lzn & lzj  |  lzl & LZN & lzj  |  lzl & lzn & LZJ  |  LZL & LZN & LZJ  ;
 mzm <=  LZL & lzn & lzj  |  lzl & LZN & lzj  |  lzl & lzn & LZJ  |  lzl & lzn & lzj  ;
 MYA <=  LYA & lyc & lxb  |  lya & LYC & lxb  |  lya & lyc & LXB  |  LYA & LYC & LXB  ;
 myb <=  LYA & lyc & lxb  |  lya & LYC & lxb  |  lya & lyc & LXB  |  lya & lyc & lxb  ;
 KZG <= HZG & hzd |  hzg & HZD ; 
 MZI <=  LZI & lzk & lze  |  lzi & LZK & lze  |  lzi & lzk & LZE  |  LZI & LZK & LZE  ;
 mzj <=  LZI & lzk & lze  |  lzi & LZK & lze  |  lzi & lzk & LZE  |  lzi & lzk & lze  ;
 MZO <=  LZO & lzq & lzm  |  lzo & LZQ & lzm  |  lzo & lzq & LZM  |  LZO & LZQ & LZM  ;
 mzp <=  LZO & lzq & lzm  |  lzo & LZQ & lzm  |  lzo & lzq & LZM  |  lzo & lzq & lzm  ;
 MZR <=  LZR & lzt & lzp  |  lzr & LZT & lzp  |  lzr & lzt & LZP  |  LZR & LZT & LZP  ;
 mzs <=  LZR & lzt & lzp  |  lzr & LZT & lzp  |  lzr & lzt & LZP  |  lzr & lzt & lzp  ;
 PBD <= NAD & ngd |  nad & NGD ; 
 KUB <= HUA & HTB ; 
 KTB <= HSB & HTA ; 
 HTB <= GTA & GSB ; 
 MVA <=  LVA & lub & lvc  |  lva & LUB & lvc  |  lva & lub & LVC  |  LVA & LUB & LVC  ;
 mvb <=  LVA & lub & lvc  |  lva & LUB & lvc  |  lva & lub & LVC  |  lva & lub & lvc  ;
 KYA <= HYA & hxb |  hya & HXB ; 
 HVA <=  GVA & gub & gvc  |  gva & GUB & gvc  |  gva & gub & GVC  |  GVA & GUB & GVC  ;
 hvb <=  GVA & gub & gvc  |  gva & GUB & gvc  |  gva & gub & GVC  |  gva & gub & gvc  ;
 MMB <= LMA & LLB ; 
 HWA <=  GWA & gwc & gvb  |  gwa & GWC & gvb  |  gwa & gwc & GVB  |  GWA & GWC & GVB  ;
 hwb <=  GWA & gwc & gvb  |  gwa & GWC & gvb  |  gwa & gwc & GVB  |  gwa & gwc & gvb  ;
 OJI <= IGB ; 
 OLI <= IGB ; 
 ONI <= IGB ; 
 OPI <= IGB ; 
 PBF <= RAF & nhb |  raf & NHB ; 
 PBG <= RAG & nhc |  rag & NHC ; 
 MEB <= LDB & LEA ; 
 MGA <= LGA & lfb |  lga & LFB ; 
 FVC <=  EUD & eve & evf  |  eud & EVE & evf  |  eud & eve & EVF  |  EUD & EVE & EVF  ;
 fvd <=  EUD & eve & evf  |  eud & EVE & evf  |  eud & eve & EVF  |  eud & eve & evf  ;
 OJD <= IFD ; 
 OLD <= IFD ; 
 OND <= IFD ; 
 OPD <= IFD ; 
 MGB <= LFB & LGA ; 
 HZM <=  GZM & gzo & gzj  |  gzm & GZO & gzj  |  gzm & gzo & GZJ  |  GZM & GZO & GZJ  ;
 hzn <=  GZM & gzo & gzj  |  gzm & GZO & gzj  |  gzm & gzo & GZJ  |  gzm & gzo & gzj  ;
 OJE <= IFE ; 
 OLE <= IFE ; 
 ONE <= IFE ; 
 OPE <= IFE ; 
 HZI <=  GZI & gzk & gzh  |  gzi & GZK & gzh  |  gzi & gzk & GZH  |  GZI & GZK & GZH  ;
 hzj <=  GZI & gzk & gzh  |  gzi & GZK & gzh  |  gzi & gzk & GZH  |  gzi & gzk & gzh  ;
 MHA <= LHA & lgb |  lha & LGB ; 
 PBH <= RAH & nhd |  rah & NHD ; 
 FZW <=  EYM & eyo & eyq  |  eym & EYO & eyq  |  eym & eyo & EYQ  |  EYM & EYO & EYQ  ;
 fzx <=  EYM & eyo & eyq  |  eym & EYO & eyq  |  eym & eyo & EYQ  |  eym & eyo & eyq  ;
 FFA <= EFA & efb |  efa & EFB ; 
 HYA <=  GYA & gyc & gxb  |  gya & GYC & gxb  |  gya & gyc & GXB  |  GYA & GYC & GXB  ;
 hyb <=  GYA & gyc & gxb  |  gya & GYC & gxb  |  gya & gyc & GXB  |  gya & gyc & gxb  ;
 FFB <= EFA & EFB ; 
 FYS <= EXL & eyz |  exl & EYZ ; 
 KZA <= HZA & hyb |  hza & HYB ; 
 KZB <= HYB & HZA ; 
 QXK <=  CAP & cco & cen  |  cap & CCO & cen  |  cap & cco & CEN  |  CAP & CCO & CEN  ;
 qxl <=  CAP & cco & cen  |  cap & CCO & cen  |  cap & cco & CEN  |  cap & cco & cen  ;
 QYR <= CYB & daa |  cyb & DAA ; 
 PFK <= PDK & PAC |  PBK & pac ; 
 PFL <= PDL & PAC |  PBL & pac ; 
 PFM <= PDM & PAD |  PBM & pad ; 
 PFN <= PDN & PAD |  PBN & pad ; 
 QXM <=  CGM & cil & ckk  |  cgm & CIL & ckk  |  cgm & cil & CKK  |  CGM & CIL & CKK  ;
 qxn <=  CGM & cil & ckk  |  cgm & CIL & ckk  |  cgm & cil & CKK  |  cgm & cil & ckk  ;
 PBJ <= RAJ & nib |  raj & NIB ; 
 PFO <= PDO & PAD |  PBO & pad ; 
 PFP <= PDP & PAD |  PBP & pad ; 
 PGA <= PEA & PAE |  PCA & pae ; 
 PGB <= PEB & PAE |  PCB & pae ; 
 QXO <=  CMJ & coi & cqh  |  cmj & COI & cqh  |  cmj & coi & CQH  |  CMJ & COI & CQH  ;
 qxp <=  CMJ & coi & cqh  |  cmj & COI & cqh  |  cmj & coi & CQH  |  cmj & coi & cqh  ;
 PGC <= PEC & PAE |  PCC & pae ; 
 PGD <= PED & PAE |  PCD & pae ; 
 PGE <= PEE & PAF |  PCE & paf ; 
 PGF <= PEF & PAF |  PCF & paf ; 
 PGG <= PEG & PAF |  PCG & paf ; 
 PGH <= PEH & PAF |  PCH & paf ; 
 QXQ <=  CSG & cuf & cwe  |  csg & CUF & cwe  |  csg & cuf & CWE  |  CSG & CUF & CWE  ;
 qxr <=  CSG & cuf & cwe  |  csg & CUF & cwe  |  csg & cuf & CWE  |  csg & cuf & cwe  ;
 PBK <= RAK & nic |  rak & NIC ; 
 PGI <=  PCI & pag & pap  |  PEI & PAG  |  PEI & PAP  ; 
 PGK <=  PCK & pag & pap  |  PEK & PAG  |  PEK & PAP  ; 
 QXS <=  CYD & dac & dcb  |  cyd & DAC & dcb  |  cyd & dac & DCB  |  CYD & DAC & DCB  ;
 qxt <=  CYD & dac & dcb  |  cyd & DAC & dcb  |  cyd & dac & DCB  |  cyd & dac & dcb  ;
 PGM <=  PCM & pah & pam  |  PEM & PAH  |  PEM & PAM  ; 
 PGO <=  PCO & pah & pam  |  PEO & PAH  |  PEO & PAM  ; 
 PBL <= RAL & nid |  ral & NID ; 
 QXV <=  CBP & cdo & cfn  |  cbp & CDO & cfn  |  cbp & cdo & CFN  |  CBP & CDO & CFN  ;
 qxw <=  CBP & cdo & cfn  |  cbp & CDO & cfn  |  cbp & cdo & CFN  |  cbp & cdo & cfn  ;
 PBN <= RAN & njb |  ran & NJB ; 
 PBO <= RAO & njc |  rao & NJC ; 
 PBP <= RAP & njd |  rap & NJD ; 
 QXG <=  CTF & cve & cxd  |  ctf & CVE & cxd  |  ctf & cve & CXD  |  CTF & CVE & CXD  ;
 qxh <=  CTF & cve & cxd  |  ctf & CVE & cxd  |  ctf & cve & CXD  |  ctf & cve & cxd  ;
 MHB <= LGB & LHA ; 
 MNB <= LNA & LMB ; 
 QXI <=  CZC & dbb & dda  |  czc & DBB & dda  |  czc & dbb & DDA  |  CZC & DBB & DDA  ;
 qxj <=  CZC & dbb & dda  |  czc & DBB & dda  |  czc & dbb & DDA  |  czc & dbb & dda  ;
 PFE <= PDE & PAB |  PBE & pab ; 
 PFF <= PDF & PAB |  PBF & pab ; 
 PFG <= PDG & PAB |  PBG & pab ; 
 PFH <= PDH & PAB |  PBH & pab ; 
 PFI <= PDI & PAC |  PBI & pac ; 
 PFJ <= PDJ & PAC |  PBJ & pac ; 
 HJB <= FIB ; 
 HPB <= GOB ; 
 HPA <= GPA ; 
 HQA <= GQA ; 
 DZQ <= CYA ; 
 FHB <= EIB ; 
 HQB <= GPB ; 
 FUD <= EUE ; 
 HSA <=  GSA & grb & gsc  |  gsa & GRB & gsc  |  gsa & grb & GSC  |  GSA & GRB & GSC  ;
 hsb <=  GSA & grb & gsc  |  gsa & GRB & gsc  |  gsa & grb & GSC  |  gsa & grb & gsc  ;
 KZH <= HZD & HZG ; 
 PBA <= NAA ; 
 PBB <= NAB ; 
 PBE <= RAE ; 
 PBI <= RAI ; 
 PBM <= RAM ; 
 PCA <= RBA ; 
 PCE <= RBE ; 
 PCI <= RBI ; 
 PCM <= RBM ; 
 PDE <= rae ; 
 PDI <= rai ; 
 PDM <= ram ; 
 PEA <= rba ; 
 PEE <= rbe ; 
 PEI <= rbi ; 
 PEM <= rbm ; 
 PAF <=  NGE & NXB & NXC & NXD & NXE  |  NHE & NXC & NXD & NXE  |  NIE & NXD & NXE  |  NJE & NXE & NXE  |  NKE  ; 
 PCB <= RBB & nkb |  rbb & NKB ; 
 PCC <= RBC & nkc |  rbc & NKC ; 
 PCD <= RBD & nkd |  rbd & NKD ; 
 PCF <= RBF & nlb |  rbf & NLB ; 
 PCG <= RBG & nlc |  rbg & NLC ; 
 PCH <= RBH & nld |  rbh & NLD ; 
 PEO <= RBO & nvc |  rbo & NVC ; 
 PEN <= RBN & nvb |  rbn & NVB ; 
 PAH <=  NIE & NXD & NXE & NXF & NXG  |  NJE & NXE & NXF & NXG  |  NKE & NXF & NXG  |  NLE & NXG & NXG  |  NME  ; 
 NEO <= MNB & MOA ; 
 QAA <= IHA ; 
 QAB <= QAA ; 
 QAC <= QAB ; 
 QAD <= QAC ; 
 QAE <= QAD ; 
 QAF <= QAE ; 
 QAG <= QAF ; 
 QAH <= QAG ; 
 NEE <= MDB & MEA ; 
 OEA <= IEA ; 
 OEB <= IEB ; 
 OEC <= IEC ; 
 OED <= IED ; 
 OEE <= IEE ; 
 OEF <= IEF ; 
 OFA <= IEA ; 
 OFB <= IEB ; 
 OFC <= IEC ; 
 OFD <= IED ; 
 OFE <= IEE ; 
 OFF <= IEF ; 
 FYD <= EYE & EXD ; 
 ohc <= iec ; 
 ohd <= ied ; 
 ohe <= iee ; 
 oga <= iea ; 
 ogb <= ieb ; 
 ogc <= iec ; 
 ogd <= ied ; 
 oge <= iee ; 
 ogf <= ief ; 
 oha <= iea ; 
 ohb <= ieb ; 
 oig <= ifg ; 
 okg <= ifg ; 
 omg <= ifg ; 
 oog <= ifg ; 
 QAI <= QAH ; 
 QAJ <= QAI ; 
 QAK <= QAJ ; 
 QAL <= QAK ; 
 ACE <= AAE ; 
 ACF <= AAE ; 
 ACG <= AAG ; 
 ACH <= AAG ; 
 ACI <= AAI ; 
 ACJ <= AAI ; 
 ACK <= AAK ; 
 ACL <= AAK ; 
 ACM <= AAM ; 
 ACN <= AAM ; 
 ACO <= AAO ; 
 ACP <= AAO ; 
 NEJ <= MIB & MJA ; 
 PCJ <= RBJ & nmb |  rbj & NMB ; 
 PCK <= RBK & nmc |  rbk & NMC ; 
 PCL <= RBL & nmd |  rbl & NMD ; 
 PCN <= RBN & nnb |  rbn & NNB ; 
 PCO <= RBO & nnc |  rbo & NNC ; 
 PCP <= RBP & nnd |  rbp & NND ; 
 PBC <= NAC & neb |  nac & NEB ; 
 QVB <=  CTG & cvf & cxe  |  ctg & CVF & cxe  |  ctg & cvf & CXE  |  CTG & CVF & CXE  ;
 qvc <=  CTG & cvf & cxe  |  ctg & CVF & cxe  |  ctg & cvf & CXE  |  ctg & cvf & cxe  ;
 BAG <= IAG & tee |  BAG & TEE ; 
 BAH <= IAH & tee |  BAH & TEE ; 
 BAO <= IAO & tef |  BAO & TEF ; 
 BAP <= IAP & tef |  BAP & TEF ; 
 BBO <= IBO & teh |  BBO & TEH ; 
 BBP <= IBP & teh |  BBP & TEH ; 
 QVD <=  CZD & dbc & ddb  |  czd & DBC & ddb  |  czd & dbc & DDB  |  CZD & DBC & DDB  ;
 qve <=  CZD & dbc & ddb  |  czd & DBC & ddb  |  czd & dbc & DDB  |  czd & dbc & ddb  ;
 BBG <= IBG & teg |  BBG & TEG ; 
 BBH <= IBH & teg |  BBH & TEG ; 
 HCB <= FCB ; 
 HDB <= FDB ; 
 OJK <= IGD ; 
 OLK <= IGD ; 
 ONK <= IGD ; 
 OPK <= IGD ; 
 OJL <= IGE ; 
 OLL <= IGE ; 
 ONL <= IGE ; 
 OPL <= IGE ; 
 OJF <= IIFF ; 
 OLF <= IIFF ; 
 ONF <= IIFF ; 
 OPF <= IIFF ; 
 HGA <= FGA & ffb |  fga & FFB ; 
 HGB <= FFB & FGA ; 
 NAF <=  MFA  |  MEB  ; 
 HHA <= FHA ; 
 HHB <= FHB ; 
 OJJ <= IGC ; 
 OLJ <= IGC ; 
 ONJ <= IGC ; 
 OPJ <= IGC ; 
 QXX <=  CHM & cjl & clk  |  chm & CJL & clk  |  chm & cjl & CLK  |  CHM & CJL & CLK  ;
 qxy <=  CHM & cjl & clk  |  chm & CJL & clk  |  chm & cjl & CLK  |  chm & cjl & clk  ;
 ACQ <= AAQ ; 
 PGN <=  PCN & pah & pam  |  PEN & PAH  |  PEN & PAM  ; 
 PGP <=  PCP & pah & pam  |  PEP & PAH  |  PEP & PAM  ; 
 QXZ <=  CNJ & cpi & crh  |  cnj & CPI & crh  |  cnj & cpi & CRH  |  CNJ & CPI & CRH  ;
 qva <=  CNJ & cpi & crh  |  cnj & CPI & crh  |  cnj & cpi & CRH  |  cnj & cpi & crh  ;
 TFA <= QAJ ; 
 TFB <= QAJ ; 
 TFC <= QAJ ; 
 TFD <= QAJ ; 
 HZT <=  GZT & gzv & gzr  |  gzt & GZV & gzr  |  gzt & gzv & GZR  |  GZT & GZV & GZR  ;
 hzu <=  GZT & gzv & gzr  |  gzt & GZV & gzr  |  gzt & gzv & GZR  |  gzt & gzv & gzr  ;
 NEG <= MFB & MGA ; 
 FZT <=  EYL & ezt & ezv  |  eyl & EZT & ezv  |  eyl & ezt & EZV  |  EYL & EZT & EZV  ;
 fzu <=  EYL & ezt & ezv  |  eyl & EZT & ezv  |  eyl & ezt & EZV  |  eyl & ezt & ezv  ;
 HZA <=  GZA & gyl & gyb  |  gza & GYL & gyb  |  gza & gyl & GYB  |  GZA & GYL & GYB  ;
 hzb <=  GZA & gyl & gyb  |  gza & GYL & gyb  |  gza & gyl & GYB  |  gza & gyl & gyb  ;
 GZK <= FZL ; 
 PAG <=  NHE & NXC & NXD & NXE & NXF  |  NIE & NXD & NXE & NXF  |  NJE & NXE & NXF  |  NKE & NXF & NXF  |  NLE  ; 
 ADA <= ABA ; 
 ADB <= ABA ; 
 ADC <= ABC ; 
 ADD <= ABC ; 
 ADE <= ABE ; 
 ADF <= ABE ; 
 ADG <= ABG ; 
 ADH <= ABG ; 
 pai <=  nxc  |  nxd  |  nxe  |  nxf  |  nxg  ; 
 ADI <= ABI ; 
 ADJ <= ABI ; 
 ADK <= ABK ; 
 ADL <= ABK ; 
 NEF <= MEB & MFA ; 
 PEF <= RBF & ntb |  rbf & NTB ; 
 ADM <= ABM ; 
 ADN <= ABM ; 
 ADO <= ABO ; 
 ADP <= ABO ; 
 ACA <= AAA ; 
 ACB <= AAA ; 
 ACC <= AAC ; 
 ACD <= AAC ; 
 MAA <= LAA ; 
 MCA <= LCA ; 
 PGJ <=  PCJ & pag & pap  |  PEJ & PAG  |  PEJ & PAP  ; 
 PGL <=  PCL & pag & pap  |  PEL & PAG  |  PEL & PAP  ; 
 OJM <= IGF ; 
 OLM <= IGF ; 
 ONM <= IGF ; 
 OPM <= IGF ; 
 end 
endmodule;

