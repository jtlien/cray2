module ib( IZZ,
 IAA, 
 IAB, 
 IAC, 
 IAD, 
 IAE, 
 IAF, 
 IAG, 
 IAH, 
 IAI, 
 IAJ, 
 IAK, 
 IAL, 
 IAM, 
 IBA, 
 IBB, 
 IBC, 
 IBD, 
 IBE, 
 IBF, 
 IBG, 
 IBH, 
 IBI, 
 IBJ, 
 IBK, 
 IBL, 
 IBM, 
 ICA, 
 ICB, 
 ICC, 
 ICD, 
 ICE, 
 ICF, 
 ICG, 
 ICH, 
 ICI, 
 ICJ, 
 ICK, 
 ICL, 
 ICM, 
 ICN, 
 ICO, 
 ICP, 
 IDA, 
 IDB, 
 IDC, 
 IDD, 
 IDE, 
 IDF, 
 IDG, 
 IDH, 
 IDI, 
 IDJ, 
 IDK, 
 IDL, 
 IDM, 
 IDN, 
 IDO, 
 IDP, 
 IEA, 
 IEB, 
 IEC, 
 IED, 
 IEE, 
 IEF, 
 IEG, 
 IEH, 
 IEI, 
 IEJ, 
 IEK, 
 IEL, 
 IEM, 
 IEN, 
 IEO, 
 IEP, 
 IFA, 
 IFB, 
 IFC, 
 IFD, 
 IFE, 
 IFFF , 
 IFG, 
 IFH, 
 IFI, 
 IGA, 
 IGB, 
 IGC, 
 IHA, 
 IHB, 
 IHC, 
 IJA, 
 IJB, 
 IJC, 
 IJD, 
 IKA, 
 IKB, 
 ILA, 
 ILB, 
 ILC, 
 IMA, 
 IMB, 
 IMC, 
 IMD, 
 IME, 
 IMF, 
 IMG, 
 INA, 
 IOA, 
 IOB, 
 IOC, 
 IOD, 
 IOG, 
 IPA, 
 IPB, 
 IPC, 
 IPD, 
 IPE, 
 IPF, 
 IQA, 
 IQB, 
 IQC, 
 IQD, 
 IQE, 
 IQF, 
 IQG, 
 IQH, 
 IQI, 
 OAA, 
 OAB, 
 OAC, 
 OAD, 
 OAE, 
 OAF, 
 OAG, 
 OAH, 
 OAI, 
 OAJ, 
 OAK, 
 OAL, 
 OAM, 
 OAN, 
 OAO, 
 OAP, 
 OBA, 
 OBB, 
 OBC, 
 OBD, 
 OBE, 
 OBF, 
 OBG, 
 OBH, 
 OBI, 
 OBJ, 
 OBK, 
 OBL, 
 OBM, 
 OBN, 
 OBO, 
 OBP, 
 OEA, 
 OEB, 
 OEC, 
 OED, 
 OEE, 
 OEF, 
 OEG, 
 OEH, 
 OEJ, 
 OEK, 
 OEL, 
 OEM, 
 OEO, 
 OEP, 
 OEQ, 
 OES, 
 OET, 
 OEU, 
 OEV, 
 OEW, 
 OEX, 
 OEY, 
 OFA, 
 OFC, 
 OGA, 
 OGB, 
 OGC, 
 OGD, 
 OGE, 
 OGF, 
 OGG, 
 OGH, 
 OGI, 
 OGJ, 
 OGK, 
 OGL, 
 OGM, 
 OGN, 
 OGO, 
 OGP, 
 OGQ, 
 OGR, 
 OGS, 
 OGT, 
 OGU, 
 OGV, 
 OGW, 
 OGX, 
 OHA, 
 OHB, 
 OHC, 
 OHD, 
 OIA, 
 OIB, 
 OIC, 
 OID, 
 OIE, 
 OJA, 
 OJB, 
 OJC, 
 OJD, 
 OJE, 
 OKA, 
 OKB, 
 OLA, 
 OLB, 
 OLC, 
 OLF, 
 OMA, 
 OMB, 
 OQB, 
 OTA, 
 OTB, 
OTC ); 
    
 input IZZ; 
 input IAA; 
 input IAB; 
 input IAC; 
 input IAD; 
 input IAE; 
 input IAF; 
 input IAG; 
 input IAH; 
 input IAI; 
 input IAJ; 
 input IAK; 
 input IAL; 
 input IAM; 
 input IBA; 
 input IBB; 
 input IBC; 
 input IBD; 
 input IBE; 
 input IBF; 
 input IBG; 
 input IBH; 
 input IBI; 
 input IBJ; 
 input IBK; 
 input IBL; 
 input IBM; 
 input ICA; 
 input ICB; 
 input ICC; 
 input ICD; 
 input ICE; 
 input ICF; 
 input ICG; 
 input ICH; 
 input ICI; 
 input ICJ; 
 input ICK; 
 input ICL; 
 input ICM; 
 input ICN; 
 input ICO; 
 input ICP; 
 input IDA; 
 input IDB; 
 input IDC; 
 input IDD; 
 input IDE; 
 input IDF; 
 input IDG; 
 input IDH; 
 input IDI; 
 input IDJ; 
 input IDK; 
 input IDL; 
 input IDM; 
 input IDN; 
 input IDO; 
 input IDP; 
 input IEA; 
 input IEB; 
 input IEC; 
 input IED; 
 input IEE; 
 input IEF; 
 input IEG; 
 input IEH; 
 input IEI; 
 input IEJ; 
 input IEK; 
 input IEL; 
 input IEM; 
 input IEN; 
 input IEO; 
 input IEP; 
 input IFA; 
 input IFB; 
 input IFC; 
 input IFD; 
 input IFE; 
 input IFFF ; 
 input IFG; 
 input IFH; 
 input IFI; 
 input IGA; 
 input IGB; 
 input IGC; 
 input IHA; 
 input IHB; 
 input IHC; 
 input IJA; 
 input IJB; 
 input IJC; 
 input IJD; 
 input IKA; 
 input IKB; 
 input ILA; 
 input ILB; 
 input ILC; 
 input IMA; 
 input IMB; 
 input IMC; 
 input IMD; 
 input IME; 
 input IMF; 
 input IMG; 
 input INA; 
 input IOA; 
 input IOB; 
 input IOC; 
 input IOD; 
 input IOG; 
 input IPA; 
 input IPB; 
 input IPC; 
 input IPD; 
 input IPE; 
 input IPF; 
 input IQA; 
 input IQB; 
 input IQC; 
 input IQD; 
 input IQE; 
 input IQF; 
 input IQG; 
 input IQH; 
 input IQI; 
 output OAA; 
 output OAB; 
 output OAC; 
 output OAD; 
 output OAE; 
 output OAF; 
 output OAG; 
 output OAH; 
 output OAI; 
 output OAJ; 
 output OAK; 
 output OAL; 
 output OAM; 
 output OAN; 
 output OAO; 
 output OAP; 
 output OBA; 
 output OBB; 
 output OBC; 
 output OBD; 
 output OBE; 
 output OBF; 
 output OBG; 
 output OBH; 
 output OBI; 
 output OBJ; 
 output OBK; 
 output OBL; 
 output OBM; 
 output OBN; 
 output OBO; 
 output OBP; 
 output OEA; 
 output OEB; 
 output OEC; 
 output OED; 
 output OEE; 
 output OEF; 
 output OEG; 
 output OEH; 
 output OEJ; 
 output OEK; 
 output OEL; 
 output OEM; 
 output OEO; 
 output OEP; 
 output OEQ; 
 output OES; 
 output OET; 
 output OEU; 
 output OEV; 
 output OEW; 
 output OEX; 
 output OEY; 
 output OFA; 
 output OFC; 
 output OGA; 
 output OGB; 
 output OGC; 
 output OGD; 
 output OGE; 
 output OGF; 
 output OGG; 
 output OGH; 
 output OGI; 
 output OGJ; 
 output OGK; 
 output OGL; 
 output OGM; 
 output OGN; 
 output OGO; 
 output OGP; 
 output OGQ; 
 output OGR; 
 output OGS; 
 output OGT; 
 output OGU; 
 output OGV; 
 output OGW; 
 output OGX; 
 output OHA; 
 output OHB; 
 output OHC; 
 output OHD; 
 output OIA; 
 output OIB; 
 output OIC; 
 output OID; 
 output OIE; 
 output OJA; 
 output OJB; 
 output OJC; 
 output OJD; 
 output OJE; 
 output OKA; 
 output OKB; 
 output OLA; 
 output OLB; 
 output OLC; 
 output OLF; 
 output OMA; 
 output OMB; 
 output OQB; 
 output OTA; 
 output OTB; 
 output OTC; 
  
  
reg  AAA ;
reg  AAB ;
reg  AAC ;
reg  AAD ;
reg  AAE ;
reg  AAF ;
reg  AAG ;
reg  AAH ;
reg  AAI ;
reg  AAJ ;
reg  AAK ;
reg  AAL ;
reg  AAM ;
reg  AAN ;
reg  AAO ;
reg  AAP ;
reg  ABA ;
reg  ABB ;
reg  ABC ;
reg  ABD ;
reg  ABE ;
reg  ABF ;
reg  ABG ;
reg  ABH ;
reg  ABI ;
reg  ABJ ;
reg  ABK ;
reg  ABL ;
reg  ABM ;
reg  ABN ;
reg  ABO ;
reg  ABP ;
reg  BAG ;
reg  BAH ;
reg  BAI ;
reg  BAJ ;
reg  BAK ;
reg  BAL ;
reg  BAM ;
reg  BAN ;
reg  BAO ;
reg  BAP ;
reg  BBA ;
reg  BBB ;
reg  BBC ;
reg  BBD ;
reg  BBE ;
reg  BBF ;
reg  BBG ;
reg  BBH ;
reg  BBI ;
reg  BBJ ;
reg  BBK ;
reg  BBL ;
reg  BBM ;
reg  BBN ;
reg  BBO ;
reg  BBP ;
reg  BCG ;
reg  BCH ;
reg  BCI ;
reg  BCJ ;
reg  BCK ;
reg  BCL ;
reg  BCM ;
reg  BCN ;
reg  BCO ;
reg  BCP ;
reg  BDA ;
reg  BDB ;
reg  BDC ;
reg  BDD ;
reg  BDE ;
reg  BDF ;
reg  BDG ;
reg  BDH ;
reg  BDI ;
reg  BDJ ;
reg  BDK ;
reg  BDL ;
reg  BDM ;
reg  BDN ;
reg  BDO ;
reg  BDP ;
reg  BEG ;
reg  BEH ;
reg  BEI ;
reg  BEJ ;
reg  BEK ;
reg  BEL ;
reg  BEM ;
reg  BEN ;
reg  BEO ;
reg  BEP ;
reg  BFA ;
reg  BFB ;
reg  BFC ;
reg  BFD ;
reg  BFE ;
reg  BFF ;
reg  BFG ;
reg  BFH ;
reg  BFI ;
reg  BFJ ;
reg  BFK ;
reg  BFL ;
reg  BFM ;
reg  BFN ;
reg  BFO ;
reg  BFP ;
reg  CAA ;
reg  CAB ;
reg  CAC ;
reg  DAA ;
reg  DAB ;
reg  DAC ;
reg  DAD ;
reg  DAE ;
reg  DAF ;
reg  DAG ;
reg  DAH ;
reg  DAI ;
reg  DAJ ;
reg  DAK ;
reg  DAL ;
reg  DAM ;
reg  DAN ;
reg  DAO ;
reg  DAP ;
reg  DBA ;
reg  DBB ;
reg  DBC ;
reg  DBD ;
reg  DBE ;
reg  DBF ;
reg  DBG ;
reg  DBH ;
reg  DBI ;
reg  DBJ ;
reg  DBK ;
reg  DBL ;
reg  DBM ;
reg  DBN ;
reg  DBO ;
reg  DBP ;
reg  eaa ;
reg  eab ;
reg  eac ;
reg  ead ;
reg  eae ;
reg  eaf ;
reg  eag ;
reg  eah ;
reg  eai ;
reg  eaj ;
reg  eak ;
reg  eal ;
reg  eam ;
reg  ean ;
reg  eao ;
reg  eap ;
reg  ebj ;
reg  ebk ;
reg  ebl ;
reg  ebp ;
reg  eci ;
reg  ecj ;
reg  eck ;
reg  ecl ;
reg  ecm ;
reg  ecn ;
reg  eco ;
reg  ecp ;
reg  EDA ;
reg  EDB ;
reg  EDC ;
reg  EDD ;
reg  EDE ;
reg  EDF ;
reg  EDG ;
reg  EDH ;
reg  EDI ;
reg  EDJ ;
reg  EDK ;
reg  EDL ;
reg  EDM ;
reg  EDN ;
reg  EDO ;
reg  EDP ;
reg  gaa ;
reg  gab ;
reg  gac ;
reg  gad ;
reg  gae ;
reg  gaf ;
reg  gag ;
reg  gah ;
reg  gai ;
reg  gal ;
reg  gam ;
reg  gan ;
reg  gao ;
reg  gap ;
reg  gba ;
reg  gbc ;
reg  gbd ;
reg  gbe ;
reg  gbf ;
reg  gbg ;
reg  gbh ;
reg  gbi ;
reg  gbj ;
reg  gbk ;
reg  gbm ;
reg  gbn ;
reg  gbo ;
reg  gbp ;
reg  gca ;
reg  gcb ;
reg  gcc ;
reg  gcd ;
reg  gch ;
reg  gci ;
reg  gcj ;
reg  gck ;
reg  gcl ;
reg  gcm ;
reg  gcn ;
reg  haa ;
reg  hab ;
reg  hac ;
reg  had ;
reg  hae ;
reg  haf ;
reg  hag ;
reg  hah ;
reg  hba ;
reg  hbb ;
reg  hbc ;
reg  hbd ;
reg  hbe ;
reg  hbf ;
reg  hbg ;
reg  hbh ;
reg  hca ;
reg  hcb ;
reg  hcc ;
reg  hcd ;
reg  hce ;
reg  hcf ;
reg  hcg ;
reg  hch ;
reg  hda ;
reg  hdb ;
reg  hdc ;
reg  hdd ;
reg  hde ;
reg  hdf ;
reg  hdg ;
reg  hdh ;
reg  hea ;
reg  heb ;
reg  hec ;
reg  hed ;
reg  hee ;
reg  hef ;
reg  heg ;
reg  heh ;
reg  hfa ;
reg  hfb ;
reg  hfc ;
reg  hfd ;
reg  hfh ;
reg  KAA ;
reg  KAB ;
reg  KAC ;
reg  KAD ;
reg  KAE ;
reg  KAF ;
reg  LAA ;
reg  LAB ;
reg  LAC ;
reg  LAD ;
reg  LAE ;
reg  LAF ;
reg  LBA ;
reg  LBB ;
reg  LBC ;
reg  LBD ;
reg  LBE ;
reg  LBF ;
reg  MAA ;
reg  MAB ;
reg  MAC ;
reg  NAA ;
reg  NAB ;
reg  NAC ;
reg  NAD ;
reg  NBA ;
reg  NBB ;
reg  NBC ;
reg  OAA ;
reg  OAB ;
reg  OAC ;
reg  OAD ;
reg  OAE ;
reg  OAF ;
reg  OAG ;
reg  OAH ;
reg  OAI ;
reg  OAJ ;
reg  OAK ;
reg  OAL ;
reg  OAM ;
reg  OAN ;
reg  OAO ;
reg  OAP ;
reg  OBA ;
reg  OBB ;
reg  OBC ;
reg  OBD ;
reg  OBE ;
reg  OBF ;
reg  OBG ;
reg  OBH ;
reg  OBI ;
reg  OBJ ;
reg  OBK ;
reg  OBL ;
reg  OBM ;
reg  OBN ;
reg  OBO ;
reg  OBP ;
reg  oca ;
reg  ocb ;
reg  occ ;
reg  ocd ;
reg  oce ;
reg  ocf ;
reg  ocg ;
reg  och ;
reg  oci ;
reg  ocj ;
reg  ock ;
reg  ocl ;
reg  ocm ;
reg  ocn ;
reg  oco ;
reg  ocp ;
reg  oda ;
reg  odb ;
reg  odc ;
reg  odd ;
reg  ode ;
reg  odf ;
reg  odg ;
reg  odh ;
reg  odi ;
reg  odj ;
reg  odk ;
reg  odl ;
reg  odm ;
reg  odn ;
reg  odo ;
reg  odp ;
reg  OEA ;
reg  OEB ;
reg  OEC ;
reg  OED ;
reg  OEE ;
reg  OEF ;
reg  OEG ;
reg  OEH ;
reg  oei ;
reg  OEJ ;
reg  OEK ;
reg  OEL ;
reg  OEM ;
reg  OEN ;
reg  OEO ;
reg  OEP ;
reg  OEQ ;
reg  oer ;
reg  OES ;
reg  OET ;
reg  OEU ;
reg  OEV ;
reg  OEW ;
reg  OEX ;
reg  OEY ;
reg  OFA ;
reg  ofb ;
reg  OFC ;
reg  OGA ;
reg  OGB ;
reg  OGC ;
reg  OGD ;
reg  OGE ;
reg  OGF ;
reg  OGG ;
reg  OGH ;
reg  OGI ;
reg  OGJ ;
reg  OGK ;
reg  OGL ;
reg  OGM ;
reg  OGN ;
reg  OGO ;
reg  OGP ;
reg  OGQ ;
reg  OGR ;
reg  OGS ;
reg  OGT ;
reg  OGU ;
reg  OGV ;
reg  OGW ;
reg  OGX ;
reg  OHA ;
reg  OHB ;
reg  OHC ;
reg  OHD ;
reg  OIA ;
reg  OIB ;
reg  OIC ;
reg  OID ;
reg  OIE ;
reg  OJA ;
reg  OJB ;
reg  OJC ;
reg  OJD ;
reg  OJE ;
reg  OKA ;
reg  OKB ;
reg  OLA ;
reg  OLB ;
reg  OLC ;
reg  old ;
reg  OLF ;
reg  OMA ;
reg  OMB ;
reg  oqa ;
reg  OQB ;
reg  ora ;
reg  orb ;
reg  orc ;
reg  ord ;
reg  ore ;
reg  orf ;
reg  OTA ;
reg  OTB ;
reg  OTC ;
reg  otd ;
reg  ote ;
reg  otf ;
reg  PAA ;
reg  PAB ;
reg  PAC ;
reg  PAD ;
reg  PAE ;
reg  PAF ;
reg  PAG ;
reg  PAH ;
reg  PAI ;
reg  PAJ ;
reg  PAK ;
reg  PAL ;
reg  PAM ;
reg  PAN ;
reg  PAO ;
reg  PAP ;
reg  PBA ;
reg  PBB ;
reg  PBC ;
reg  PBD ;
reg  PBE ;
reg  PBF ;
reg  PBG ;
reg  PBH ;
reg  PBI ;
reg  PBJ ;
reg  PBK ;
reg  PBL ;
reg  PBM ;
reg  PBN ;
reg  PBO ;
reg  PBP ;
reg  PCA ;
reg  PCB ;
reg  PCC ;
reg  PCD ;
reg  PCE ;
reg  PCF ;
reg  PCG ;
reg  PCH ;
reg  PCI ;
reg  PCJ ;
reg  PCK ;
reg  PCL ;
reg  PCM ;
reg  PCN ;
reg  PCO ;
reg  PCP ;
reg  PDA ;
reg  PDB ;
reg  PDC ;
reg  PDD ;
reg  PDE ;
reg  PDF ;
reg  PDG ;
reg  PDH ;
reg  PDI ;
reg  PDJ ;
reg  PDK ;
reg  PDL ;
reg  PDM ;
reg  PDN ;
reg  PDO ;
reg  PDP ;
reg  PEA ;
reg  PEB ;
reg  PEC ;
reg  PED ;
reg  PEE ;
reg  PEF ;
reg  PEG ;
reg  PEH ;
reg  PEI ;
reg  PEJ ;
reg  PEK ;
reg  PEL ;
reg  PEM ;
reg  PEN ;
reg  PEO ;
reg  PEP ;
reg  PFA ;
reg  PFB ;
reg  PFC ;
reg  PFD ;
reg  PFE ;
reg  PFF ;
reg  PFG ;
reg  PFH ;
reg  PFI ;
reg  PFJ ;
reg  PFK ;
reg  PFL ;
reg  PFM ;
reg  PFN ;
reg  PFO ;
reg  PFP ;
reg  QAA ;
reg  QAB ;
reg  QAC ;
reg  QAD ;
reg  QBA ;
reg  QCA ;
reg  QCC ;
reg  QEA ;
reg  QEB ;
reg  QFA ;
reg  QFB ;
reg  qfc ;
reg  QGA ;
reg  QGB ;
reg  QGC ;
reg  QGD ;
reg  QGE ;
reg  QHA ;
reg  QHC ;
reg  QHD ;
reg  QHE ;
reg  QHF ;
reg  qia ;
reg  qib ;
reg  qic ;
reg  qid ;
reg  QKA ;
reg  QKB ;
reg  QKC ;
reg  QKD ;
reg  QKE ;
reg  QKF ;
reg  QKG ;
reg  QKH ;
reg  QKI ;
reg  QKJ ;
reg  QKK ;
reg  QKL ;
reg  QKM ;
reg  QKN ;
reg  QLA ;
reg  QLB ;
reg  QLC ;
reg  QLD ;
reg  QLE ;
reg  QLF ;
reg  QLG ;
reg  QLI ;
reg  QLJ ;
reg  QLK ;
reg  QLL ;
reg  QLM ;
reg  QLN ;
reg  QLO ;
reg  QLP ;
reg  QLQ ;
reg  QLR ;
reg  QLS ;
reg  qma ;
reg  qmb ;
reg  qmc ;
reg  qme ;
reg  qmf ;
reg  qmg ;
reg  qmi ;
reg  qmj ;
reg  QMK ;
reg  qna ;
reg  qnb ;
reg  qnc ;
reg  QND ;
reg  qne ;
reg  qnf ;
reg  qng ;
reg  qni ;
reg  qnj ;
reg  qnm ;
reg  qnn ;
reg  qnq ;
reg  qnr ;
reg  qnu ;
reg  qnv ;
reg  qoa ;
reg  qpa ;
reg  qpb ;
reg  qpc ;
reg  qpd ;
reg  QQA ;
reg  QQB ;
reg  QQC ;
reg  QQD ;
reg  QQE ;
reg  QQF ;
reg  QQG ;
reg  QQH ;
reg  QQI ;
reg  QQJ ;
reg  QQK ;
reg  QQL ;
reg  QQM ;
reg  QQN ;
reg  QQW ;
reg  qqx ;
reg  QRA ;
reg  QRB ;
reg  QRC ;
reg  QRD ;
reg  QRE ;
reg  QRF ;
reg  QSA ;
reg  QSB ;
reg  QSC ;
reg  QSD ;
reg  QSE ;
reg  QSF ;
reg  QSG ;
reg  QSH ;
reg  qsi ;
reg  QTA ;
reg  QTB ;
reg  QTC ;
reg  QTD ;
reg  QTE ;
reg  QTF ;
reg  QTG ;
reg  QTH ;
reg  QTI ;
reg  QTJ ;
reg  QTM ;
reg  QTN ;
reg  qtp ;
reg  qtq ;
reg  qtr ;
reg  QTW ;
reg  QTX ;
reg  QUA ;
reg  QUB ;
reg  QUC ;
reg  QUD ;
reg  QUE ;
reg  QUF ;
reg  qva ;
reg  qvb ;
reg  qvc ;
reg  qvd ;
reg  qve ;
reg  qvf ;
reg  qvg ;
reg  qvh ;
reg  qvi ;
reg  qvj ;
reg  QWA ;
reg  QWB ;
reg  QWC ;
reg  qwd ;
reg  qwe ;
reg  qwf ;
reg  qwg ;
reg  qwh ;
reg  qwi ;
reg  QWJ ;
reg  QXA ;
reg  QXB ;
reg  QXC ;
reg  QXD ;
reg  QXE ;
reg  QXF ;
reg  QYA ;
reg  QYB ;
reg  QYC ;
reg  QYD ;
reg  qza ;
reg  qzb ;
reg  QZD ;
reg  QZE ;
reg  QZF ;
reg  RAA ;
reg  RAB ;
reg  RAC ;
reg  RAD ;
reg  RAE ;
reg  RAF ;
reg  RAG ;
reg  rba ;
reg  RBB ;
reg  RBC ;
reg  RBD ;
reg  RBE ;
reg  RBF ;
reg  RBG ;
reg  REB ;
reg  REC ;
reg  RFA ;
reg  RFB ;
reg  RGA ;
reg  RGB ;
reg  RGC ;
reg  RGD ;
reg  RHA ;
reg  RHB ;
reg  RHC ;
reg  RHD ;
reg  RHE ;
reg  RHF ;
reg  RHG ;
reg  RHH ;
reg  RHI ;
reg  RHJ ;
reg  RIA ;
reg  RIB ;
reg  RIC ;
reg  RID ;
reg  RIE ;
reg  RIF ;
reg  RIX ;
reg  RJA ;
reg  RJB ;
reg  RJC ;
reg  RJD ;
reg  RJE ;
reg  RJF ;
reg  RJG ;
reg  RJH ;
reg  RJI ;
reg  RJK ;
reg  RJL ;
reg  RKA ;
reg  RKB ;
reg  RKC ;
reg  RKD ;
reg  RLA ;
reg  RLB ;
reg  RLC ;
reg  RLD ;
reg  RMA ;
reg  RMB ;
reg  RMC ;
reg  RMD ;
reg  RME ;
reg  RMF ;
reg  RMG ;
reg  RMH ;
reg  RMI ;
reg  RMJ ;
reg  RMK ;
reg  RML ;
reg  RMM ;
reg  RMN ;
reg  RMO ;
reg  RMP ;
reg  RMQ ;
reg  RMR ;
reg  RMS ;
reg  RMT ;
reg  RMU ;
reg  RNA ;
reg  RNB ;
reg  RNC ;
reg  RND ;
reg  RNK ;
reg  RNL ;
reg  RNM ;
reg  RNN ;
reg  RNO ;
reg  RNP ;
reg  rqa ;
reg  RQB ;
reg  rqc ;
reg  RRA ;
reg  RRB ;
reg  RRC ;
reg  RRD ;
reg  RRE ;
reg  RRF ;
reg  RRG ;
reg  RRH ;
reg  RSA ;
reg  RSB ;
reg  RSC ;
wire  aaa ;
wire  aab ;
wire  aac ;
wire  aad ;
wire  aae ;
wire  aaf ;
wire  aag ;
wire  aah ;
wire  aai ;
wire  aaj ;
wire  aak ;
wire  aal ;
wire  aam ;
wire  aan ;
wire  aao ;
wire  aap ;
wire  aba ;
wire  abb ;
wire  abc ;
wire  abd ;
wire  abe ;
wire  abf ;
wire  abg ;
wire  abh ;
wire  abi ;
wire  abj ;
wire  abk ;
wire  abl ;
wire  abm ;
wire  abn ;
wire  abo ;
wire  abp ;
wire  bag ;
wire  bah ;
wire  bai ;
wire  baj ;
wire  bak ;
wire  bal ;
wire  bam ;
wire  ban ;
wire  bao ;
wire  bap ;
wire  bba ;
wire  bbb ;
wire  bbc ;
wire  bbd ;
wire  bbe ;
wire  bbf ;
wire  bbg ;
wire  bbh ;
wire  bbi ;
wire  bbj ;
wire  bbk ;
wire  bbl ;
wire  bbm ;
wire  bbn ;
wire  bbo ;
wire  bbp ;
wire  bcg ;
wire  bch ;
wire  bci ;
wire  bcj ;
wire  bck ;
wire  bcl ;
wire  bcm ;
wire  bcn ;
wire  bco ;
wire  bcp ;
wire  bda ;
wire  bdb ;
wire  bdc ;
wire  bdd ;
wire  bde ;
wire  bdf ;
wire  bdg ;
wire  bdh ;
wire  bdi ;
wire  bdj ;
wire  bdk ;
wire  bdl ;
wire  bdm ;
wire  bdn ;
wire  bdo ;
wire  bdp ;
wire  beg ;
wire  beh ;
wire  bei ;
wire  bej ;
wire  bek ;
wire  bel ;
wire  bem ;
wire  ben ;
wire  beo ;
wire  bep ;
wire  bfa ;
wire  bfb ;
wire  bfc ;
wire  bfd ;
wire  bfe ;
wire  bff ;
wire  bfg ;
wire  bfh ;
wire  bfi ;
wire  bfj ;
wire  bfk ;
wire  bfl ;
wire  bfm ;
wire  bfn ;
wire  bfo ;
wire  bfp ;
wire  caa ;
wire  cab ;
wire  cac ;
wire  daa ;
wire  dab ;
wire  dac ;
wire  dad ;
wire  dae ;
wire  daf ;
wire  dag ;
wire  dah ;
wire  dai ;
wire  daj ;
wire  dak ;
wire  dal ;
wire  dam ;
wire  dan ;
wire  dao ;
wire  dap ;
wire  dba ;
wire  dbb ;
wire  dbc ;
wire  dbd ;
wire  dbe ;
wire  dbf ;
wire  dbg ;
wire  dbh ;
wire  dbi ;
wire  dbj ;
wire  dbk ;
wire  dbl ;
wire  dbm ;
wire  dbn ;
wire  dbo ;
wire  dbp ;
wire  EAA ;
wire  EAB ;
wire  EAC ;
wire  EAD ;
wire  EAE ;
wire  EAF ;
wire  EAG ;
wire  EAH ;
wire  EAI ;
wire  EAJ ;
wire  EAK ;
wire  EAL ;
wire  EAM ;
wire  EAN ;
wire  EAO ;
wire  EAP ;
wire  EBJ ;
wire  EBK ;
wire  EBL ;
wire  EBP ;
wire  ECI ;
wire  ECJ ;
wire  ECK ;
wire  ECL ;
wire  ECM ;
wire  ECN ;
wire  ECO ;
wire  ECP ;
wire  eda ;
wire  edb ;
wire  edc ;
wire  edd ;
wire  ede ;
wire  edf ;
wire  edg ;
wire  edh ;
wire  edi ;
wire  edj ;
wire  edk ;
wire  edl ;
wire  edm ;
wire  edn ;
wire  edo ;
wire  edp ;
wire  faa ;
wire  FAA ;
wire  fab ;
wire  FAB ;
wire  fac ;
wire  FAC ;
wire  fad ;
wire  FAD ;
wire  fae ;
wire  FAE ;
wire  faf ;
wire  FAF ;
wire  fag ;
wire  FAG ;
wire  fah ;
wire  FAH ;
wire  fai ;
wire  FAI ;
wire  faj ;
wire  FAJ ;
wire  fak ;
wire  FAK ;
wire  fal ;
wire  FAL ;
wire  fap ;
wire  FAP ;
wire  fba ;
wire  FBA ;
wire  fbb ;
wire  FBB ;
wire  fbc ;
wire  FBC ;
wire  fbd ;
wire  FBD ;
wire  fbe ;
wire  FBE ;
wire  fbg ;
wire  FBG ;
wire  fbh ;
wire  FBH ;
wire  GAA ;
wire  GAB ;
wire  GAC ;
wire  GAD ;
wire  GAE ;
wire  GAF ;
wire  GAG ;
wire  GAH ;
wire  GAI ;
wire  GAL ;
wire  GAM ;
wire  GAN ;
wire  GAO ;
wire  GAP ;
wire  GBA ;
wire  GBC ;
wire  GBD ;
wire  GBE ;
wire  GBF ;
wire  GBG ;
wire  GBH ;
wire  GBI ;
wire  GBJ ;
wire  GBK ;
wire  GBM ;
wire  GBN ;
wire  GBO ;
wire  GBP ;
wire  GCA ;
wire  GCB ;
wire  GCC ;
wire  GCD ;
wire  GCH ;
wire  GCI ;
wire  GCJ ;
wire  GCK ;
wire  GCL ;
wire  GCM ;
wire  GCN ;
wire  HAA ;
wire  HAB ;
wire  HAC ;
wire  HAD ;
wire  HAE ;
wire  HAF ;
wire  HAG ;
wire  HAH ;
wire  HBA ;
wire  HBB ;
wire  HBC ;
wire  HBD ;
wire  HBE ;
wire  HBF ;
wire  HBG ;
wire  HBH ;
wire  HCA ;
wire  HCB ;
wire  HCC ;
wire  HCD ;
wire  HCE ;
wire  HCF ;
wire  HCG ;
wire  HCH ;
wire  HDA ;
wire  HDB ;
wire  HDC ;
wire  HDD ;
wire  HDE ;
wire  HDF ;
wire  HDG ;
wire  HDH ;
wire  HEA ;
wire  HEB ;
wire  HEC ;
wire  HED ;
wire  HEE ;
wire  HEF ;
wire  HEG ;
wire  HEH ;
wire  HFA ;
wire  HFB ;
wire  HFC ;
wire  HFD ;
wire  HFH ;
wire  iaa ;
wire  iab ;
wire  iac ;
wire  iad ;
wire  iae ;
wire  iaf ;
wire  iag ;
wire  iah ;
wire  iai ;
wire  iaj ;
wire  iak ;
wire  ial ;
wire  iam ;
wire  iba ;
wire  ibb ;
wire  ibc ;
wire  ibd ;
wire  ibe ;
wire  ibf ;
wire  ibg ;
wire  ibh ;
wire  ibi ;
wire  ibj ;
wire  ibk ;
wire  ibl ;
wire  ibm ;
wire  ica ;
wire  icb ;
wire  icc ;
wire  icd ;
wire  ice ;
wire  icf ;
wire  icg ;
wire  ich ;
wire  ici ;
wire  icj ;
wire  ick ;
wire  icl ;
wire  icm ;
wire  icn ;
wire  ico ;
wire  icp ;
wire  ida ;
wire  idb ;
wire  idc ;
wire  idd ;
wire  ide ;
wire  idf ;
wire  idg ;
wire  idh ;
wire  idi ;
wire  idj ;
wire  idk ;
wire  idl ;
wire  idm ;
wire  idn ;
wire  ido ;
wire  idp ;
wire  iea ;
wire  ieb ;
wire  iec ;
wire  ied ;
wire  iee ;
wire  ief ;
wire  ieg ;
wire  ieh ;
wire  iei ;
wire  iej ;
wire  iek ;
wire  iel ;
wire  iem ;
wire  ien ;
wire  ieo ;
wire  iep ;
wire  ifa ;
wire  ifb ;
wire  ifc ;
wire  ifd ;
wire  ife ;
wire  ifff  ;
wire  ifg ;
wire  ifh ;
wire  ifi ;
wire  iga ;
wire  igb ;
wire  igc ;
wire  iha ;
wire  ihb ;
wire  ihc ;
wire  ija ;
wire  ijb ;
wire  ijc ;
wire  ijd ;
wire  ika ;
wire  ikb ;
wire  ila ;
wire  ilb ;
wire  ilc ;
wire  ima ;
wire  imb ;
wire  imc ;
wire  imd ;
wire  ime ;
wire  imf ;
wire  img ;
wire  ina ;
wire  ioa ;
wire  iob ;
wire  ioc ;
wire  iod ;
wire  iog ;
wire  ipa ;
wire  ipb ;
wire  ipc ;
wire  ipd ;
wire  ipe ;
wire  ipf ;
wire  iqa ;
wire  iqb ;
wire  iqc ;
wire  iqd ;
wire  iqe ;
wire  iqf ;
wire  iqg ;
wire  iqh ;
wire  iqi ;
wire  jad ;
wire  JAD ;
wire  jae ;
wire  JAE ;
wire  jaf ;
wire  JAF ;
wire  jai ;
wire  JAI ;
wire  jaj ;
wire  JAJ ;
wire  jak ;
wire  JAK ;
wire  jal ;
wire  JAL ;
wire  jam ;
wire  JAM ;
wire  jan ;
wire  JAN ;
wire  jao ;
wire  JAO ;
wire  jap ;
wire  JAP ;
wire  jaq ;
wire  JAQ ;
wire  jar ;
wire  JAR ;
wire  jba ;
wire  JBA ;
wire  jbb ;
wire  JBB ;
wire  jbc ;
wire  JBC ;
wire  jbd ;
wire  JBD ;
wire  jbe ;
wire  JBE ;
wire  jca ;
wire  JCA ;
wire  jcb ;
wire  JCB ;
wire  jcc ;
wire  JCC ;
wire  jcd ;
wire  JCD ;
wire  jce ;
wire  JCE ;
wire  jcf ;
wire  JCF ;
wire  jcg ;
wire  JCG ;
wire  jch ;
wire  JCH ;
wire  jci ;
wire  JCI ;
wire  jcj ;
wire  JCJ ;
wire  jck ;
wire  JCK ;
wire  jcl ;
wire  JCL ;
wire  jcm ;
wire  JCM ;
wire  jcn ;
wire  JCN ;
wire  jco ;
wire  JCO ;
wire  jcp ;
wire  JCP ;
wire  jcq ;
wire  JCQ ;
wire  jcr ;
wire  JCR ;
wire  jcs ;
wire  JCS ;
wire  jct ;
wire  JCT ;
wire  jda ;
wire  JDA ;
wire  jdb ;
wire  JDB ;
wire  jdc ;
wire  JDC ;
wire  jdd ;
wire  JDD ;
wire  jde ;
wire  JDE ;
wire  jdf ;
wire  JDF ;
wire  jdg ;
wire  JDG ;
wire  jdh ;
wire  JDH ;
wire  jdi ;
wire  JDI ;
wire  jdj ;
wire  JDJ ;
wire  jdk ;
wire  JDK ;
wire  jdl ;
wire  JDL ;
wire  jdm ;
wire  JDM ;
wire  jdn ;
wire  JDN ;
wire  jdo ;
wire  JDO ;
wire  jdp ;
wire  JDP ;
wire  jea ;
wire  JEA ;
wire  jeb ;
wire  JEB ;
wire  jec ;
wire  JEC ;
wire  jed ;
wire  JED ;
wire  jee ;
wire  JEE ;
wire  jef ;
wire  JEF ;
wire  jeg ;
wire  JEG ;
wire  jeh ;
wire  JEH ;
wire  jei ;
wire  JEI ;
wire  jej ;
wire  JEJ ;
wire  jek ;
wire  JEK ;
wire  jel ;
wire  JEL ;
wire  jem ;
wire  JEM ;
wire  jen ;
wire  JEN ;
wire  jeo ;
wire  JEO ;
wire  jep ;
wire  JEP ;
wire  jfa ;
wire  JFA ;
wire  jfb ;
wire  JFB ;
wire  jfc ;
wire  JFC ;
wire  jfd ;
wire  JFD ;
wire  jfe ;
wire  JFE ;
wire  jff ;
wire  JFF ;
wire  jfg ;
wire  JFG ;
wire  jfh ;
wire  JFH ;
wire  jfi ;
wire  JFI ;
wire  jfj ;
wire  JFJ ;
wire  jga ;
wire  JGA ;
wire  jgb ;
wire  JGB ;
wire  jgc ;
wire  JGC ;
wire  jgd ;
wire  JGD ;
wire  jge ;
wire  JGE ;
wire  jgf ;
wire  JGF ;
wire  jgg ;
wire  JGG ;
wire  jgh ;
wire  JGH ;
wire  jgi ;
wire  JGI ;
wire  jgj ;
wire  JGJ ;
wire  jgk ;
wire  JGK ;
wire  jgl ;
wire  JGL ;
wire  jgm ;
wire  JGM ;
wire  jgn ;
wire  JGN ;
wire  jgo ;
wire  JGO ;
wire  jgp ;
wire  JGP ;
wire  jha ;
wire  JHA ;
wire  jhb ;
wire  JHB ;
wire  jhc ;
wire  JHC ;
wire  jhd ;
wire  JHD ;
wire  jhe ;
wire  JHE ;
wire  jhf ;
wire  JHF ;
wire  jhg ;
wire  JHG ;
wire  jhh ;
wire  JHH ;
wire  jhi ;
wire  JHI ;
wire  jhj ;
wire  JHJ ;
wire  jhk ;
wire  JHK ;
wire  jhl ;
wire  JHL ;
wire  jhm ;
wire  JHM ;
wire  jhn ;
wire  JHN ;
wire  jho ;
wire  JHO ;
wire  jhp ;
wire  JHP ;
wire  jic ;
wire  JIC ;
wire  jid ;
wire  JID ;
wire  jja ;
wire  JJA ;
wire  jjb ;
wire  JJB ;
wire  jjc ;
wire  JJC ;
wire  jjd ;
wire  JJD ;
wire  jje ;
wire  JJE ;
wire  jjf ;
wire  JJF ;
wire  jjg ;
wire  JJG ;
wire  jjh ;
wire  JJH ;
wire  jji ;
wire  JJI ;
wire  jjj ;
wire  JJJ ;
wire  jjk ;
wire  JJK ;
wire  jjl ;
wire  JJL ;
wire  jjm ;
wire  JJM ;
wire  jjn ;
wire  JJN ;
wire  jjp ;
wire  JJP ;
wire  jka ;
wire  JKA ;
wire  jkb ;
wire  JKB ;
wire  jkc ;
wire  JKC ;
wire  jkd ;
wire  JKD ;
wire  jke ;
wire  JKE ;
wire  jla ;
wire  JLA ;
wire  jlb ;
wire  JLB ;
wire  jlc ;
wire  JLC ;
wire  jld ;
wire  JLD ;
wire  jle ;
wire  JLE ;
wire  jlf ;
wire  JLF ;
wire  jlg ;
wire  JLG ;
wire  jma ;
wire  JMA ;
wire  jmb ;
wire  JMB ;
wire  jna ;
wire  JNA ;
wire  jnb ;
wire  JNB ;
wire  jnc ;
wire  JNC ;
wire  jnd ;
wire  JND ;
wire  jne ;
wire  JNE ;
wire  jpa ;
wire  JPA ;
wire  jqa ;
wire  JQA ;
wire  jqb ;
wire  JQB ;
wire  jqc ;
wire  JQC ;
wire  jqd ;
wire  JQD ;
wire  jqe ;
wire  JQE ;
wire  jqf ;
wire  JQF ;
wire  jra ;
wire  JRA ;
wire  jrb ;
wire  JRB ;
wire  jrc ;
wire  JRC ;
wire  jrd ;
wire  JRD ;
wire  jre ;
wire  JRE ;
wire  jsa ;
wire  JSA ;
wire  jsb ;
wire  JSB ;
wire  jsc ;
wire  JSC ;
wire  jsd ;
wire  JSD ;
wire  jtb ;
wire  JTB ;
wire  jxa ;
wire  JXA ;
wire  jxb ;
wire  JXB ;
wire  kaa ;
wire  kab ;
wire  kac ;
wire  kad ;
wire  kae ;
wire  kaf ;
wire  laa ;
wire  lab ;
wire  lac ;
wire  lad ;
wire  lae ;
wire  laf ;
wire  lba ;
wire  lbb ;
wire  lbc ;
wire  lbd ;
wire  lbe ;
wire  lbf ;
wire  maa ;
wire  mab ;
wire  mac ;
wire  naa ;
wire  nab ;
wire  nac ;
wire  nad ;
wire  nba ;
wire  nbb ;
wire  nbc ;
wire  oaa ;
wire  oab ;
wire  oac ;
wire  oad ;
wire  oae ;
wire  oaf ;
wire  oag ;
wire  oah ;
wire  oai ;
wire  oaj ;
wire  oak ;
wire  oal ;
wire  oam ;
wire  oan ;
wire  oao ;
wire  oap ;
wire  oba ;
wire  obb ;
wire  obc ;
wire  obd ;
wire  obe ;
wire  obf ;
wire  obg ;
wire  obh ;
wire  obi ;
wire  obj ;
wire  obk ;
wire  obl ;
wire  obm ;
wire  obn ;
wire  obo ;
wire  obp ;
wire  OCA ;
wire  OCB ;
wire  OCC ;
wire  OCD ;
wire  OCE ;
wire  OCF ;
wire  OCG ;
wire  OCH ;
wire  OCI ;
wire  OCJ ;
wire  OCK ;
wire  OCL ;
wire  OCM ;
wire  OCN ;
wire  OCO ;
wire  OCP ;
wire  ODA ;
wire  ODB ;
wire  ODC ;
wire  ODD ;
wire  ODE ;
wire  ODF ;
wire  ODG ;
wire  ODH ;
wire  ODI ;
wire  ODJ ;
wire  ODK ;
wire  ODL ;
wire  ODM ;
wire  ODN ;
wire  ODO ;
wire  ODP ;
wire  oea ;
wire  oeb ;
wire  oec ;
wire  oed ;
wire  oee ;
wire  oef ;
wire  oeg ;
wire  oeh ;
wire  OEI ;
wire  oej ;
wire  oek ;
wire  oel ;
wire  oem ;
wire  oen ;
wire  oeo ;
wire  oep ;
wire  oeq ;
wire  OER ;
wire  oes ;
wire  oet ;
wire  oeu ;
wire  oev ;
wire  oew ;
wire  oex ;
wire  oey ;
wire  ofa ;
wire  OFB ;
wire  ofc ;
wire  oga ;
wire  ogb ;
wire  ogc ;
wire  ogd ;
wire  oge ;
wire  ogf ;
wire  ogg ;
wire  ogh ;
wire  ogi ;
wire  ogj ;
wire  ogk ;
wire  ogl ;
wire  ogm ;
wire  ogn ;
wire  ogo ;
wire  ogp ;
wire  ogq ;
wire  ogr ;
wire  ogs ;
wire  ogt ;
wire  ogu ;
wire  ogv ;
wire  ogw ;
wire  ogx ;
wire  oha ;
wire  ohb ;
wire  ohc ;
wire  ohd ;
wire  oia ;
wire  oib ;
wire  oic ;
wire  oid ;
wire  oie ;
wire  oja ;
wire  ojb ;
wire  ojc ;
wire  ojd ;
wire  oje ;
wire  oka ;
wire  okb ;
wire  ola ;
wire  olb ;
wire  olc ;
wire  OLD ;
wire  olf ;
wire  oma ;
wire  omb ;
wire  OQA ;
wire  oqb ;
wire  ORA ;
wire  ORB ;
wire  ORC ;
wire  ORD ;
wire  ORE ;
wire  ORF ;
wire  ota ;
wire  otb ;
wire  otc ;
wire  OTD ;
wire  OTE ;
wire  OTF ;
wire  paa ;
wire  pab ;
wire  pac ;
wire  pad ;
wire  pae ;
wire  paf ;
wire  pag ;
wire  pah ;
wire  pai ;
wire  paj ;
wire  pak ;
wire  pal ;
wire  pam ;
wire  pan ;
wire  pao ;
wire  pap ;
wire  pba ;
wire  pbb ;
wire  pbc ;
wire  pbd ;
wire  pbe ;
wire  pbf ;
wire  pbg ;
wire  pbh ;
wire  pbi ;
wire  pbj ;
wire  pbk ;
wire  pbl ;
wire  pbm ;
wire  pbn ;
wire  pbo ;
wire  pbp ;
wire  pca ;
wire  pcb ;
wire  pcc ;
wire  pcd ;
wire  pce ;
wire  pcf ;
wire  pcg ;
wire  pch ;
wire  pci ;
wire  pcj ;
wire  pck ;
wire  pcl ;
wire  pcm ;
wire  pcn ;
wire  pco ;
wire  pcp ;
wire  pda ;
wire  pdb ;
wire  pdc ;
wire  pdd ;
wire  pde ;
wire  pdf ;
wire  pdg ;
wire  pdh ;
wire  pdi ;
wire  pdj ;
wire  pdk ;
wire  pdl ;
wire  pdm ;
wire  pdn ;
wire  pdo ;
wire  pdp ;
wire  pea ;
wire  peb ;
wire  pec ;
wire  ped ;
wire  pee ;
wire  pef ;
wire  peg ;
wire  peh ;
wire  pei ;
wire  pej ;
wire  pek ;
wire  pel ;
wire  pem ;
wire  pen ;
wire  peo ;
wire  pep ;
wire  pfa ;
wire  pfb ;
wire  pfc ;
wire  pfd ;
wire  pfe ;
wire  pff ;
wire  pfg ;
wire  pfh ;
wire  pfi ;
wire  pfj ;
wire  pfk ;
wire  pfl ;
wire  pfm ;
wire  pfn ;
wire  pfo ;
wire  pfp ;
wire  qaa ;
wire  qab ;
wire  qac ;
wire  qad ;
wire  qba ;
wire  qca ;
wire  qcc ;
wire  qea ;
wire  qeb ;
wire  qfa ;
wire  qfb ;
wire  QFC ;
wire  qga ;
wire  qgb ;
wire  qgc ;
wire  qgd ;
wire  qge ;
wire  qha ;
wire  qhc ;
wire  qhd ;
wire  qhe ;
wire  qhf ;
wire  QIA ;
wire  QIB ;
wire  QIC ;
wire  QID ;
wire  qka ;
wire  qkb ;
wire  qkc ;
wire  qkd ;
wire  qke ;
wire  qkf ;
wire  qkg ;
wire  qkh ;
wire  qki ;
wire  qkj ;
wire  qkk ;
wire  qkl ;
wire  qkm ;
wire  qkn ;
wire  qla ;
wire  qlb ;
wire  qlc ;
wire  qld ;
wire  qle ;
wire  qlf ;
wire  qlg ;
wire  qli ;
wire  qlj ;
wire  qlk ;
wire  qll ;
wire  qlm ;
wire  qln ;
wire  qlo ;
wire  qlp ;
wire  qlq ;
wire  qlr ;
wire  qls ;
wire  QMA ;
wire  QMB ;
wire  QMC ;
wire  QME ;
wire  QMF ;
wire  QMG ;
wire  QMI ;
wire  QMJ ;
wire  qmk ;
wire  QNA ;
wire  QNB ;
wire  QNC ;
wire  qnd ;
wire  QNE ;
wire  QNF ;
wire  QNG ;
wire  QNI ;
wire  QNJ ;
wire  QNM ;
wire  QNN ;
wire  QNQ ;
wire  QNR ;
wire  QNU ;
wire  QNV ;
wire  QOA ;
wire  QPA ;
wire  QPB ;
wire  QPC ;
wire  QPD ;
wire  qqa ;
wire  qqb ;
wire  qqc ;
wire  qqd ;
wire  qqe ;
wire  qqf ;
wire  qqg ;
wire  qqh ;
wire  qqi ;
wire  qqj ;
wire  qqk ;
wire  qql ;
wire  qqm ;
wire  qqn ;
wire  qqw ;
wire  QQX ;
wire  qra ;
wire  qrb ;
wire  qrc ;
wire  qrd ;
wire  qre ;
wire  qrf ;
wire  qsa ;
wire  qsb ;
wire  qsc ;
wire  qsd ;
wire  qse ;
wire  qsf ;
wire  qsg ;
wire  qsh ;
wire  QSI ;
wire  qta ;
wire  qtb ;
wire  qtc ;
wire  qtd ;
wire  qte ;
wire  qtf ;
wire  qtg ;
wire  qth ;
wire  qti ;
wire  qtj ;
wire  qtm ;
wire  qtn ;
wire  QTP ;
wire  QTQ ;
wire  QTR ;
wire  qtw ;
wire  qtx ;
wire  qua ;
wire  qub ;
wire  quc ;
wire  qud ;
wire  que ;
wire  quf ;
wire  QVA ;
wire  QVB ;
wire  QVC ;
wire  QVD ;
wire  QVE ;
wire  QVF ;
wire  QVG ;
wire  QVH ;
wire  QVI ;
wire  QVJ ;
wire  qwa ;
wire  qwb ;
wire  qwc ;
wire  QWD ;
wire  QWE ;
wire  QWF ;
wire  QWG ;
wire  QWH ;
wire  QWI ;
wire  qwj ;
wire  qxa ;
wire  qxb ;
wire  qxc ;
wire  qxd ;
wire  qxe ;
wire  qxf ;
wire  qya ;
wire  qyb ;
wire  qyc ;
wire  qyd ;
wire  QZA ;
wire  QZB ;
wire  qzd ;
wire  qze ;
wire  qzf ;
wire  raa ;
wire  rab ;
wire  rac ;
wire  rad ;
wire  rae ;
wire  raf ;
wire  rag ;
wire  RBA ;
wire  rbb ;
wire  rbc ;
wire  rbd ;
wire  rbe ;
wire  rbf ;
wire  rbg ;
wire  reb ;
wire  rec ;
wire  rfa ;
wire  rfb ;
wire  rga ;
wire  rgb ;
wire  rgc ;
wire  rgd ;
wire  rha ;
wire  rhb ;
wire  rhc ;
wire  rhd ;
wire  rhe ;
wire  rhf ;
wire  rhg ;
wire  rhh ;
wire  rhi ;
wire  rhj ;
wire  ria ;
wire  rib ;
wire  ric ;
wire  rid ;
wire  rie ;
wire  rif ;
wire  rix ;
wire  rja ;
wire  rjb ;
wire  rjc ;
wire  rjd ;
wire  rje ;
wire  rjf ;
wire  rjg ;
wire  rjh ;
wire  rji ;
wire  rjk ;
wire  rjl ;
wire  rka ;
wire  rkb ;
wire  rkc ;
wire  rkd ;
wire  rla ;
wire  rlb ;
wire  rlc ;
wire  rld ;
wire  rma ;
wire  rmb ;
wire  rmc ;
wire  rmd ;
wire  rme ;
wire  rmf ;
wire  rmg ;
wire  rmh ;
wire  rmi ;
wire  rmj ;
wire  rmk ;
wire  rml ;
wire  rmm ;
wire  rmn ;
wire  rmo ;
wire  rmp ;
wire  rmq ;
wire  rmr ;
wire  rms ;
wire  rmt ;
wire  rmu ;
wire  rna ;
wire  rnb ;
wire  rnc ;
wire  rnd ;
wire  rnk ;
wire  rnl ;
wire  rnm ;
wire  rnn ;
wire  rno ;
wire  rnp ;
wire  RQA ;
wire  rqb ;
wire  RQC ;
wire  rra ;
wire  rrb ;
wire  rrc ;
wire  rrd ;
wire  rre ;
wire  rrf ;
wire  rrg ;
wire  rrh ;
wire  rsa ;
wire  rsb ;
wire  rsc ;
wire  taa ;
wire  TAA ;
wire  tab ;
wire  TAB ;
wire  tac ;
wire  TAC ;
wire  tad ;
wire  TAD ;
wire  tae ;
wire  TAE ;
wire  taf ;
wire  TAF ;
wire  tag ;
wire  TAG ;
wire  tah ;
wire  TAH ;
wire  tba ;
wire  TBA ;
wire  tbb ;
wire  TBB ;
wire  tbc ;
wire  TBC ;
wire  tbd ;
wire  TBD ;
wire  tbe ;
wire  TBE ;
wire  tbf ;
wire  TBF ;
wire  tbg ;
wire  TBG ;
wire  tbh ;
wire  TBH ;
wire  tca ;
wire  TCA ;
wire  tcb ;
wire  TCB ;
wire  tcc ;
wire  TCC ;
wire  tcd ;
wire  TCD ;
wire  tce ;
wire  TCE ;
wire  tcf ;
wire  TCF ;
wire  tcg ;
wire  TCG ;
wire  tch ;
wire  TCH ;
wire  tda ;
wire  TDA ;
wire  tdb ;
wire  TDB ;
wire  tdc ;
wire  TDC ;
wire  tdd ;
wire  TDD ;
wire  tde ;
wire  TDE ;
wire  tdf ;
wire  TDF ;
wire  tdg ;
wire  TDG ;
wire  tdh ;
wire  TDH ;
wire  tea ;
wire  TEA ;
wire  teb ;
wire  TEB ;
wire  tec ;
wire  TEC ;
wire  ted ;
wire  TED ;
wire  tee ;
wire  TEE ;
wire  tef ;
wire  TEF ;
wire  tfa ;
wire  TFA ;
wire  tfb ;
wire  TFB ;
wire  tfc ;
wire  TFC ;
wire  tfd ;
wire  TFD ;
wire  tga ;
wire  TGA ;
wire  tgb ;
wire  TGB ;
wire  tgc ;
wire  TGC ;
wire  tgd ;
wire  TGD ;
wire  tge ;
wire  TGE ;
wire  tgf ;
wire  TGF ;
wire  tha ;
wire  THA ;
wire  tla ;
wire  TLA ;
wire  tlb ;
wire  TLB ;
wire  tlc ;
wire  TLC ;
wire  tld ;
wire  TLD ;
wire  tma ;
wire  TMA ;
wire  tmb ;
wire  TMB ;
wire  tmc ;
wire  TMC ;
wire  tmd ;
wire  TMD ;
wire  tpa ;
wire  TPA ;
wire  tpb ;
wire  TPB ;
wire  tpc ;
wire  TPC ;
wire  tpd ;
wire  TPD ;
wire  tpe ;
wire  TPE ;
wire  waa ;
wire  WAA ;
wire  wab ;
wire  WAB ;
wire  wac ;
wire  WAC ;
wire  wad ;
wire  WAD ;
wire  wae ;
wire  WAE ;
wire  waf ;
wire  WAF ;
wire  wag ;
wire  WAG ;
wire  wah ;
wire  WAH ;
wire  wai ;
wire  WAI ;
wire  waj ;
wire  WAJ ;
wire  wak ;
wire  WAK ;
wire  wal ;
wire  WAL ;
wire  wam ;
wire  WAM ;
wire  wan ;
wire  WAN ;
wire  wao ;
wire  WAO ;
wire  wap ;
wire  WAP ;
wire  wba ;
wire  WBA ;
wire  wbb ;
wire  WBB ;
wire  wbc ;
wire  WBC ;
wire  wbd ;
wire  WBD ;
wire  wbe ;
wire  WBE ;
wire  wbf ;
wire  WBF ;
wire  wbg ;
wire  WBG ;
wire  wbh ;
wire  WBH ;
wire  wbi ;
wire  WBI ;
wire  wbj ;
wire  WBJ ;
wire  wbk ;
wire  WBK ;
wire  wbl ;
wire  WBL ;
wire  wbm ;
wire  WBM ;
wire  wbn ;
wire  WBN ;
wire  wbo ;
wire  WBO ;
wire  wbp ;
wire  WBP ;
wire  wca ;
wire  WCA ;
wire  wcb ;
wire  WCB ;
wire  wcc ;
wire  WCC ;
wire  wcd ;
wire  WCD ;
wire  wce ;
wire  WCE ;
wire  wcf ;
wire  WCF ;
wire  wcg ;
wire  WCG ;
wire  wch ;
wire  WCH ;
wire  wci ;
wire  WCI ;
wire  wcj ;
wire  WCJ ;
wire  wck ;
wire  WCK ;
wire  wcl ;
wire  WCL ;
wire  wcm ;
wire  WCM ;
wire  wcn ;
wire  WCN ;
wire  wco ;
wire  WCO ;
wire  wcp ;
wire  WCP ;
wire  wda ;
wire  WDA ;
wire  wdb ;
wire  WDB ;
wire  wdc ;
wire  WDC ;
wire  wdd ;
wire  WDD ;
wire  wde ;
wire  WDE ;
wire  wdf ;
wire  WDF ;
wire  wdg ;
wire  WDG ;
wire  wdh ;
wire  WDH ;
wire  wdi ;
wire  WDI ;
wire  wdj ;
wire  WDJ ;
wire  wdk ;
wire  WDK ;
wire  wdl ;
wire  WDL ;
wire  wdm ;
wire  WDM ;
wire  wdn ;
wire  WDN ;
wire  wdo ;
wire  WDO ;
wire  wdp ;
wire  WDP ;
wire  ZZI ;
wire  ZZO ;
assign ZZI = 1'b1;
assign ZZO = 1'b0;
assign paa = ~PAA;  //complement 
assign pca = ~PCA;  //complement 
assign pea = ~PEA;  //complement 
assign JGA =  QVA  ; 
assign jga = ~JGA;  //complement  
assign JGI =  QVD  ; 
assign jgi = ~JGI;  //complement 
assign JPA =  QVA & paa  |  qva & PAA  ; 
assign jpa = ~JPA; //complement 
assign JDI =  QWD  ; 
assign jdi = ~JDI;  //complement  
assign pai = ~PAI;  //complement 
assign pci = ~PCI;  //complement 
assign pei = ~PEI;  //complement 
assign QVA = ~qva;  //complement 
assign QVJ = ~qvj;  //complement 
assign bai = ~BAI;  //complement 
assign bci = ~BCI;  //complement 
assign bei = ~BEI;  //complement 
assign pba = ~PBA;  //complement 
assign pda = ~PDA;  //complement 
assign pfa = ~PFA;  //complement 
assign JFA =  PEB & PEC & PED  ; 
assign jfa = ~JFA;  //complement  
assign JFC =  PEI & PEJ & PEK & PEL  ; 
assign jfc = ~JFC;  //complement 
assign bba = ~BBA;  //complement 
assign bda = ~BDA;  //complement 
assign bfa = ~BFA;  //complement 
assign JDB =  BEI & BEJ & BEK & BEL  ; 
assign jdb = ~JDB;  //complement  
assign JDD =  BFA & BFB & BFC & BFD  ; 
assign jdd = ~JDD;  //complement 
assign pbi = ~PBI;  //complement 
assign pdi = ~PDI;  //complement 
assign pfi = ~PFI;  //complement 
assign JHA =  QVF  ; 
assign jha = ~JHA;  //complement  
assign JHI =  QVG & QVI  ; 
assign jhi = ~JHI;  //complement 
assign bbi = ~BBI;  //complement 
assign bdi = ~BDI;  //complement 
assign bfi = ~BFI;  //complement 
assign JEA =  QWF  ; 
assign jea = ~JEA;  //complement  
assign JEI =  QWH  ; 
assign jei = ~JEI;  //complement 
assign HBA = ~hba;  //complement 
assign HCA = ~hca;  //complement 
assign HDA = ~hda;  //complement 
assign HEA = ~hea;  //complement 
assign HBB = ~hbb;  //complement 
assign HCB = ~hcb;  //complement 
assign HDB = ~hdb;  //complement 
assign HEB = ~heb;  //complement 
assign HBC = ~hbc;  //complement 
assign HCC = ~hcc;  //complement 
assign HDC = ~hdc;  //complement 
assign HEC = ~hec;  //complement 
assign HBD = ~hbd;  //complement 
assign HCD = ~hcd;  //complement 
assign HDD = ~hdd;  //complement 
assign HED = ~hed;  //complement 
assign HBE = ~hbe;  //complement 
assign HCE = ~hce;  //complement 
assign HDE = ~hde;  //complement 
assign HEE = ~hee;  //complement 
assign HBF = ~hbf;  //complement 
assign HCF = ~hcf;  //complement 
assign HDF = ~hdf;  //complement 
assign HEF = ~hef;  //complement 
assign HBG = ~hbg;  //complement 
assign HCG = ~hcg;  //complement 
assign HDG = ~hdg;  //complement 
assign HEG = ~heg;  //complement 
assign HBH = ~hbh;  //complement 
assign HCH = ~hch;  //complement 
assign HDH = ~hdh;  //complement 
assign HEH = ~heh;  //complement 
assign HFA = ~hfa;  //complement 
assign HFB = ~hfb;  //complement 
assign HFC = ~hfc;  //complement 
assign HFD = ~hfd;  //complement 
assign HFH = ~hfh;  //complement 
assign jaq = qtm & hdf ; 
assign JAQ = ~jaq ; //complement 
assign jar = qtm & hef ; 
assign JAR = ~jar ;  //complement 
assign GAA = ~gaa;  //complement 
assign GAI = ~gai;  //complement 
assign FAA =  ebp & eao & ean & eam  ; 
assign faa = ~FAA;  //complement  
assign FAI =  eal & eak & eaj  ; 
assign fai = ~FAI;  //complement 
assign jfj =  gbc & gbd & gbe & gbf & gbg & gae  ; 
assign JFJ = ~jfj;  //complement  
assign jfi =  gbn & gbi & gbj  ; 
assign JFI = ~jfi;  //complement 
assign GBA = ~gba;  //complement 
assign GBI = ~gbi;  //complement 
assign FBA =  ebl & ebk  ; 
assign fba = ~FBA;  //complement  
assign QPA = ~qpa;  //complement 
assign QPB = ~qpb;  //complement 
assign GCA = ~gca;  //complement 
assign GCI = ~gci;  //complement 
assign HAE = ~hae;  //complement 
assign HAF = ~haf;  //complement 
assign HAA = ~haa;  //complement 
assign HAB = ~hab;  //complement 
assign HAC = ~hac;  //complement 
assign HAD = ~had;  //complement 
assign qxe = ~QXE;  //complement 
assign qxf = ~QXF;  //complement 
assign naa = ~NAA;  //complement 
assign nba = ~NBA;  //complement 
assign qtw = ~QTW;  //complement 
assign qtx = ~QTX;  //complement 
assign JBE =  HAF & hac & had  ; 
assign jbe = ~JBE;  //complement 
assign qtf = ~QTF;  //complement 
assign qtg = ~QTG;  //complement 
assign qth = ~QTH;  //complement 
assign qti = ~QTI;  //complement 
assign JAD =  HED & HEE  ; 
assign jad = ~JAD;  //complement 
assign JAE =  HEA & HEF  ; 
assign jae = ~JAE;  //complement 
assign JAF =  HEB & HEF  ; 
assign jaf = ~JAF;  //complement 
assign JCT =  QTP  ; 
assign jct = ~JCT;  //complement 
assign JAI = HEG & HEA ; 
assign jai = ~JAI ; //complement 
assign JAJ = HEG & HEB ; 
assign jaj = ~JAJ ;  //complement 
assign JAK = HEG & HEC ; 
assign jak = ~JAK ;  //complement 
assign JAL = HEG & HED; 
assign jal = ~JAL; 
assign qnd = ~QND;  //complement 
assign QOA = ~qoa;  //complement 
assign JAM = HFH & HFA ; 
assign jam = ~JAM ; //complement 
assign JAN = HFH & HFB ; 
assign jan = ~JAN ;  //complement 
assign JAO = HFH & HFC ; 
assign jao = ~JAO ;  //complement 
assign JAP = HFH & HFD; 
assign jap = ~JAP; 
assign lba = ~LBA;  //complement 
assign JLA =  QLE  ; 
assign jla = ~JLA;  //complement  
assign EAA = ~eaa;  //complement 
assign WAA =  AAA & QXA  ; 
assign waa = ~WAA;  //complement 
assign WAI =  BAI & qxa  |  AAI & QXA  ; 
assign wai = ~WAI;  //complement 
assign aaa = ~AAA;  //complement 
assign oaa = ~OAA;  //complement 
assign oai = ~OAI;  //complement 
assign EAI = ~eai;  //complement 
assign ECI = ~eci;  //complement 
assign daa = ~DAA;  //complement 
assign dai = ~DAI;  //complement 
assign eda = ~EDA;  //complement 
assign edi = ~EDI;  //complement 
assign aai = ~AAI;  //complement 
assign ogc = ~OGC;  //complement 
assign wca = aaa; 
assign WCA = ~wca; //complement 
assign wci = aai; 
assign WCI = ~wci;  //complement 
assign wda = aba; 
assign WDA = ~wda;  //complement 
assign wdi = abi; 
assign WDI = ~wdi;  //complement 
assign taa = rjd; 
assign TAA = ~taa; //complement 
assign tab = rjd; 
assign TAB = ~tab;  //complement 
assign tac = rjd; 
assign TAC = ~tac;  //complement 
assign tad = rjd; 
assign TAD = ~tad;  //complement 
assign dba = ~DBA;  //complement 
assign dbi = ~DBI;  //complement 
assign aba = ~ABA;  //complement 
assign ogk = ~OGK;  //complement 
assign otb = ~OTB;  //complement 
assign ORA = ~ora;  //complement 
assign JSC =  QQI & NBA & NBB  ; 
assign jsc = ~JSC;  //complement 
assign JSA =  QQI  ; 
assign jsa = ~JSA;  //complement 
assign JSB =  QQI & NBA  ; 
assign jsb = ~JSB;  //complement 
assign WBA =  BBA & qxb  |  ABA & QXB  ; 
assign wba = ~WBA;  //complement 
assign WBI =  BBI & qxb  |  ABI & QXB  ; 
assign wbi = ~WBI;  //complement 
assign ogs = ~OGS;  //complement 
assign abi = ~ABI;  //complement 
assign oba = ~OBA;  //complement 
assign obi = ~OBI;  //complement 
assign qtb = ~QTB;  //complement 
assign qtc = ~QTC;  //complement 
assign qtd = ~QTD;  //complement 
assign qte = ~QTE;  //complement 
assign qta = ~QTA;  //complement 
assign tma = qtn; 
assign TMA = ~tma; //complement 
assign tmb = qtn; 
assign TMB = ~tmb;  //complement 
assign tmc = qtn; 
assign TMC = ~tmc;  //complement 
assign tmd = qtn; 
assign TMD = ~tmd;  //complement 
assign OCA = ~oca;  //complement 
assign OCI = ~oci;  //complement 
assign ODA = ~oda;  //complement 
assign ODI = ~odi;  //complement 
assign JNA =  MAA & QNG  |  NAA & RQC  ; 
assign jna = ~JNA;  //complement 
assign qgc = ~QGC;  //complement 
assign qge = ~QGE;  //complement 
assign qtm = ~QTM;  //complement 
assign qtn = ~QTN;  //complement 
assign qgd = ~QGD;  //complement 
assign QTP = ~qtp;  //complement 
assign JMA =  QOA  ; 
assign jma = ~JMA;  //complement 
assign JMB =  QOA & KAA  ; 
assign jmb = ~JMB;  //complement 
assign JND =  QNG  ; 
assign jnd = ~JND;  //complement 
assign qtj = ~QTJ;  //complement 
assign qzd = ~QZD;  //complement 
assign qya = ~QYA;  //complement 
assign qyb = ~QYB;  //complement 
assign qyc = ~QYC;  //complement 
assign qyd = ~QYD;  //complement 
assign oea = ~OEA;  //complement 
assign kaa = ~KAA;  //complement 
assign qze = ~QZE;  //complement 
assign laa = ~LAA;  //complement 
assign pab = ~PAB;  //complement 
assign pcb = ~PCB;  //complement 
assign peb = ~PEB;  //complement 
assign JGB =  QVB  ; 
assign jgb = ~JGB;  //complement  
assign JGJ =  QVD & PCI  ; 
assign jgj = ~JGJ;  //complement 
assign JDJ =  QWD & BCI  ; 
assign jdj = ~JDJ;  //complement  
assign paj = ~PAJ;  //complement 
assign pcj = ~PCJ;  //complement 
assign pej = ~PEJ;  //complement 
assign QVH = ~qvh;  //complement 
assign QVI = ~qvi;  //complement 
assign baj = ~BAJ;  //complement 
assign bcj = ~BCJ;  //complement 
assign bej = ~BEJ;  //complement 
assign qwb = ~QWB;  //complement 
assign qwc = ~QWC;  //complement 
assign QWI = ~qwi;  //complement 
assign pbb = ~PBB;  //complement 
assign pdb = ~PDB;  //complement 
assign pfb = ~PFB;  //complement 
assign JFE =  PFA & PFB & PFC & PFD  ; 
assign jfe = ~JFE;  //complement  
assign JFG =  PFI & PFJ & PFK & PFL  ; 
assign jfg = ~JFG;  //complement 
assign bbb = ~BBB;  //complement 
assign bdb = ~BDB;  //complement 
assign bfb = ~BFB;  //complement 
assign JDF =  BFI & BFJ & BFK & BFL  ; 
assign jdf = ~JDF;  //complement  
assign pbj = ~PBJ;  //complement 
assign pdj = ~PDJ;  //complement 
assign pfj = ~PFJ;  //complement 
assign JHB =  QVF & PDA  ; 
assign jhb = ~JHB;  //complement  
assign JHJ =  QVG & QVI & PDI  ; 
assign jhj = ~JHJ;  //complement 
assign bbj = ~BBJ;  //complement 
assign bdj = ~BDJ;  //complement 
assign bfj = ~BFJ;  //complement 
assign JEB =  QWF & BDA  ; 
assign jeb = ~JEB;  //complement  
assign JEJ =  QWH & BDI  ; 
assign jej = ~JEJ;  //complement 
assign rha = ~RHA;  //complement 
assign rhb = ~RHB;  //complement 
assign rhc = ~RHC;  //complement 
assign rhd = ~RHD;  //complement 
assign rhe = ~RHE;  //complement 
assign rhf = ~RHF;  //complement 
assign rhg = ~RHG;  //complement 
assign rhh = ~RHH;  //complement 
assign rhi = ~RHI;  //complement 
assign rhj = ~RHJ;  //complement 
assign ria = ~RIA;  //complement 
assign rib = ~RIB;  //complement 
assign ric = ~RIC;  //complement 
assign rid = ~RID;  //complement 
assign rie = ~RIE;  //complement 
assign rif = ~RIF;  //complement 
assign jic =  qha & rha & rhb & rhc & rhd & rhe  ; 
assign JIC = ~jic;  //complement  
assign jid =  rhf & rhg & rhh & rhi & rhj & qhc  ; 
assign JID = ~jid;  //complement  
assign jrb =  ria & rib & ric & rid & rie & rif  ; 
assign JRB = ~jrb;  //complement  
assign GAB = ~gab;  //complement 
assign FAB =  ebp & eao & ean & EAM  ; 
assign fab = ~FAB;  //complement  
assign FAJ =  eal & eak & EAJ  ; 
assign faj = ~FAJ;  //complement 
assign GBJ = ~gbj;  //complement 
assign FBB =  ebl & EBK  ; 
assign fbb = ~FBB;  //complement  
assign QPC = ~qpc;  //complement 
assign QPD = ~qpd;  //complement 
assign GCB = ~gcb;  //complement 
assign GCJ = ~gcj;  //complement 
assign HAG = ~hag;  //complement 
assign HAH = ~hah;  //complement 
assign nab = ~NAB;  //complement 
assign nbb = ~NBB;  //complement 
assign qha = ~QHA;  //complement 
assign qkf = ~QKF;  //complement 
assign qkg = ~QKG;  //complement 
assign qkh = ~QKH;  //complement 
assign qki = ~QKI;  //complement 
assign qkk = ~QKK;  //complement 
assign JBB =  qkf & QKG  |  QKF & QKH  |  QKI  |  RJI  ; 
assign jbb = ~JBB;  //complement 
assign qkl = ~QKL;  //complement 
assign qkm = ~QKM;  //complement 
assign qkn = ~QKN;  //complement 
assign lbb = ~LBB;  //complement 
assign JLB =  QLE & lba  ; 
assign jlb = ~JLB;  //complement  
assign EAB = ~eab;  //complement 
assign WAB =  AAB & QXA  ; 
assign wab = ~WAB;  //complement 
assign WAJ =  BAJ & qxa  |  AAJ & QXA  ; 
assign waj = ~WAJ;  //complement 
assign aab = ~AAB;  //complement 
assign oab = ~OAB;  //complement 
assign oaj = ~OAJ;  //complement 
assign EAJ = ~eaj;  //complement 
assign EBJ = ~ebj;  //complement 
assign ECJ = ~ecj;  //complement 
assign dab = ~DAB;  //complement 
assign daj = ~DAJ;  //complement 
assign edb = ~EDB;  //complement 
assign edj = ~EDJ;  //complement 
assign aaj = ~AAJ;  //complement 
assign ogd = ~OGD;  //complement 
assign wcb = aab; 
assign WCB = ~wcb; //complement 
assign wcj = aaj; 
assign WCJ = ~wcj;  //complement 
assign wdb = abb; 
assign WDB = ~wdb;  //complement 
assign wdj = abj; 
assign WDJ = ~wdj;  //complement 
assign TBA = QZA; 
assign tba = ~TBA; //complement 
assign TBB = QZA; 
assign tbb = ~TBB;  //complement 
assign tbc = qza; 
assign TBC = ~tbc;  //complement 
assign tbd = qza; 
assign TBD = ~tbd;  //complement 
assign dbb = ~DBB;  //complement 
assign dbj = ~DBJ;  //complement 
assign abb = ~ABB;  //complement 
assign ogl = ~OGL;  //complement 
assign ORB = ~orb;  //complement 
assign JSD =  QQI & NBA & NBB & NBC  ; 
assign jsd = ~JSD;  //complement  
assign WBB =  BBB & qxb  |  ABB & QXB  ; 
assign wbb = ~WBB;  //complement 
assign WBJ =  BBJ & qxb  |  ABJ & QXB  ; 
assign wbj = ~WBJ;  //complement 
assign ogt = ~OGT;  //complement 
assign abj = ~ABJ;  //complement 
assign obb = ~OBB;  //complement 
assign obj = ~OBJ;  //complement 
assign qkj = ~QKJ;  //complement 
assign QZA = ~qza;  //complement 
assign QZB = ~qzb;  //complement 
assign TBE = QZB; 
assign tbe = ~TBE; //complement 
assign TBF = QZB; 
assign tbf = ~TBF;  //complement 
assign TBG = QZB; 
assign tbg = ~TBG;  //complement 
assign TBH = QZB; 
assign tbh = ~TBH;  //complement 
assign OCB = ~ocb;  //complement 
assign OCJ = ~ocj;  //complement 
assign ODB = ~odb;  //complement 
assign ODJ = ~odj;  //complement 
assign JNB =  MAB & QNG  |  NAB & RQC  ; 
assign jnb = ~JNB;  //complement 
assign JNE =  QNG  |  RQC  ; 
assign jne = ~JNE;  //complement 
assign oja = ~OJA;  //complement 
assign rfa = ~RFA;  //complement 
assign jba =  qga & qgb  ; 
assign JBA = ~jba;  //complement 
assign qga = ~QGA;  //complement 
assign ojb = ~OJB;  //complement 
assign rfb = ~RFB;  //complement 
assign JBC = RGA & ~cab & ~caa  |  RGB & ~cab & caa  |  RGC & cab & ~caa  |  RGD & cab & caa; 
assign jbc = ~JBC;  //complement 
assign JBD = RGA & ~cab & ~caa  |         RGB & ~cab & caa  |  RGC & cab & ~caa  |  RGD & cab & caa ; 
assign jbd = ~JBD;  //complement 
assign caa = ~CAA;  //complement 
assign cab = ~CAB;  //complement 
assign cac = ~CAC;  //complement 
assign oeb = ~OEB;  //complement 
assign kab = ~KAB;  //complement 
assign rga = ~RGA;  //complement 
assign rgb = ~RGB;  //complement 
assign rgc = ~RGC;  //complement 
assign rgd = ~RGD;  //complement 
assign lab = ~LAB;  //complement 
assign pac = ~PAC;  //complement 
assign pcc = ~PCC;  //complement 
assign pec = ~PEC;  //complement 
assign JGC =  QVB & PCB  ; 
assign jgc = ~JGC;  //complement  
assign JGK =  QVD & PCI & PCJ  ; 
assign jgk = ~JGK;  //complement 
assign TFA = QWA; 
assign tfa = ~TFA; //complement 
assign TFB = QWA; 
assign tfb = ~TFB;  //complement 
assign TPA = QWJ; 
assign tpa = ~TPA;  //complement 
assign TPB = QWJ; 
assign tpb = ~TPB;  //complement 
assign JDK =  QWD & BCI & BCJ  ; 
assign jdk = ~JDK;  //complement  
assign TPE =  QWJ  ; 
assign tpe = ~TPE;  //complement 
assign pak = ~PAK;  //complement 
assign pck = ~PCK;  //complement 
assign pek = ~PEK;  //complement 
assign qub = ~QUB;  //complement 
assign quc = ~QUC;  //complement 
assign que = ~QUE;  //complement 
assign bak = ~BAK;  //complement 
assign bck = ~BCK;  //complement 
assign bek = ~BEK;  //complement 
assign qwa = ~QWA;  //complement 
assign qwj = ~QWJ;  //complement 
assign pbc = ~PBC;  //complement 
assign pdc = ~PDC;  //complement 
assign pfc = ~PFC;  //complement 
assign qua = ~QUA;  //complement 
assign bbc = ~BBC;  //complement 
assign bdc = ~BDC;  //complement 
assign bfc = ~BFC;  //complement 
assign pbk = ~PBK;  //complement 
assign pdk = ~PDK;  //complement 
assign pfk = ~PFK;  //complement 
assign JHC =  QVF & PDA & PDB  ; 
assign jhc = ~JHC;  //complement  
assign JHK =  QVG & QVI & PDI & PDJ  ; 
assign jhk = ~JHK;  //complement 
assign bbk = ~BBK;  //complement 
assign bdk = ~BDK;  //complement 
assign bfk = ~BFK;  //complement 
assign JEC =  QWF & BDA & BDB  ; 
assign jec = ~JEC;  //complement  
assign JEK =  QWH & BDI & BDJ  ; 
assign jek = ~JEK;  //complement 
assign rma = ~RMA;  //complement 
assign rmc = ~RMC;  //complement 
assign rmd = ~RMD;  //complement 
assign rnm = ~RNM;  //complement 
assign rnn = ~RNN;  //complement 
assign rno = ~RNO;  //complement 
assign rnp = ~RNP;  //complement 
assign rmk = ~RMK;  //complement 
assign rmg = ~RMG;  //complement 
assign rmh = ~RMH;  //complement 
assign rmi = ~RMI;  //complement 
assign rmj = ~RMJ;  //complement 
assign rmn = ~RMN;  //complement 
assign rml = ~RML;  //complement 
assign rmm = ~RMM;  //complement 
assign rmo = ~RMO;  //complement 
assign rmp = ~RMP;  //complement 
assign rmf = ~RMF;  //complement 
assign rmr = ~RMR;  //complement 
assign rmq = ~RMQ;  //complement 
assign rms = ~RMS;  //complement 
assign rmt = ~RMT;  //complement 
assign rmu = ~RMU;  //complement 
assign GAC = ~gac;  //complement 
assign FAC =  ebp & eao & ean  ; 
assign fac = ~FAC;  //complement  
assign FAK =  eal & EAK & eaj  ; 
assign fak = ~FAK;  //complement 
assign GBC = ~gbc;  //complement 
assign GBK = ~gbk;  //complement 
assign FBC =  EBL & ebk  ; 
assign fbc = ~FBC;  //complement  
assign qkb = ~QKB;  //complement 
assign GCC = ~gcc;  //complement 
assign GCK = ~gck;  //complement 
assign QNI = ~qni;  //complement 
assign QNM = ~qnm;  //complement 
assign jrc =  rna & rnb & rnc & rnd  ; 
assign JRC = ~jrc;  //complement  
assign qka = ~QKA;  //complement 
assign rnl = ~RNL;  //complement 
assign QNJ = ~qnj;  //complement 
assign QNN = ~qnn;  //complement 
assign nac = ~NAC;  //complement 
assign nbc = ~NBC;  //complement 
assign rnb = ~RNB;  //complement 
assign rnc = ~RNC;  //complement 
assign rnd = ~RND;  //complement 
assign rna = ~RNA;  //complement 
assign rnk = ~RNK;  //complement 
assign rme = ~RME;  //complement 
assign rmb = ~RMB;  //complement 
assign JCN =  RAG & QKJ  ; 
assign jcn = ~JCN;  //complement 
assign JJA =  RBG  ; 
assign jja = ~JJA;  //complement 
assign lbc = ~LBC;  //complement 
assign JLC =  QLE & lba & lbb  ; 
assign jlc = ~JLC;  //complement  
assign EAC = ~eac;  //complement 
assign WAC =  AAC & QXA  ; 
assign wac = ~WAC;  //complement 
assign WAK =  BAK & qxa  |  AAK & QXA  ; 
assign wak = ~WAK;  //complement 
assign aac = ~AAC;  //complement 
assign oha = ~OHA;  //complement 
assign oac = ~OAC;  //complement 
assign oak = ~OAK;  //complement 
assign EAK = ~eak;  //complement 
assign EBK = ~ebk;  //complement 
assign ECK = ~eck;  //complement 
assign dac = ~DAC;  //complement 
assign dak = ~DAK;  //complement 
assign edc = ~EDC;  //complement 
assign edk = ~EDK;  //complement 
assign aak = ~AAK;  //complement 
assign oge = ~OGE;  //complement 
assign wcc = aac; 
assign WCC = ~wcc; //complement 
assign wck = aak; 
assign WCK = ~wck;  //complement 
assign wdc = abc; 
assign WDC = ~wdc;  //complement 
assign wdk = abk; 
assign WDK = ~wdk;  //complement 
assign tca = qxe; 
assign TCA = ~tca; //complement 
assign tcb = qxe; 
assign TCB = ~tcb;  //complement 
assign tcc = qxe; 
assign TCC = ~tcc;  //complement 
assign tcd = qxe; 
assign TCD = ~tcd;  //complement 
assign dbc = ~DBC;  //complement 
assign dbk = ~DBK;  //complement 
assign qzf = ~QZF;  //complement 
assign abc = ~ABC;  //complement 
assign ogm = ~OGM;  //complement 
assign ORC = ~orc;  //complement 
assign maa = ~MAA;  //complement 
assign WBC =  BBC & qxb  |  ABC & QXB  ; 
assign wbc = ~WBC;  //complement 
assign WBK =  BBK & qxb  |  ABK & QXB  ; 
assign wbk = ~WBK;  //complement 
assign abk = ~ABK;  //complement 
assign ogu = ~OGU;  //complement 
assign obc = ~OBC;  //complement 
assign obk = ~OBK;  //complement 
assign qfa = ~QFA;  //complement 
assign OCC = ~occ;  //complement 
assign OCK = ~ock;  //complement 
assign ODC = ~odc;  //complement 
assign ODK = ~odk;  //complement 
assign JNC =  MAC & QNG  ; 
assign jnc = ~JNC;  //complement 
assign qgb = ~QGB;  //complement 
assign qkc = ~QKC;  //complement 
assign qkd = ~QKD;  //complement 
assign qke = ~QKE;  //complement 
assign oka = ~OKA;  //complement 
assign oec = ~OEC;  //complement 
assign kac = ~KAC;  //complement 
assign okb = ~OKB;  //complement 
assign lac = ~LAC;  //complement 
assign pad = ~PAD;  //complement 
assign pcd = ~PCD;  //complement 
assign ped = ~PED;  //complement 
assign JGD =  QVB & PCB & PCC  ; 
assign jgd = ~JGD;  //complement  
assign JGL =  QVD & PCI & PCJ & PCK  ; 
assign jgl = ~JGL;  //complement 
assign JDL =  QWD & BCI & BCJ & BCK  ; 
assign jdl = ~JDL;  //complement  
assign pal = ~PAL;  //complement 
assign pcl = ~PCL;  //complement 
assign pel = ~PEL;  //complement 
assign QVB = ~qvb;  //complement 
assign bal = ~BAL;  //complement 
assign bcl = ~BCL;  //complement 
assign bel = ~BEL;  //complement 
assign QWD = ~qwd;  //complement 
assign pbd = ~PBD;  //complement 
assign pdd = ~PDD;  //complement 
assign pfd = ~PFD;  //complement 
assign qud = ~QUD;  //complement 
assign bbd = ~BBD;  //complement 
assign bdd = ~BDD;  //complement 
assign bfd = ~BFD;  //complement 
assign pbl = ~PBL;  //complement 
assign pdl = ~PDL;  //complement 
assign pfl = ~PFL;  //complement 
assign JHL =  QVG & QVI & PDI & PDJ & PDK  ; 
assign jhl = ~JHL;  //complement  
assign JHD =  QVF & PDA & PDB & PDC  ; 
assign jhd = ~JHD;  //complement 
assign bbl = ~BBL;  //complement 
assign bdl = ~BDL;  //complement 
assign bfl = ~BFL;  //complement 
assign JED =  QWF & BDA & BDB & BDC  ; 
assign jed = ~JED;  //complement  
assign JEL =  QWH & BDI & BDJ & BDK  ; 
assign jel = ~JEL;  //complement 
assign jka =  qlf & rka & rkb & rkc & rkd  ; 
assign JKA = ~jka;  //complement  
assign JKB =  QLL & QLM  ; 
assign jkb = ~JKB;  //complement 
assign rkb = ~RKB;  //complement 
assign rkc = ~RKC;  //complement 
assign rkd = ~RKD;  //complement 
assign rlb = ~RLB;  //complement 
assign rlc = ~RLC;  //complement 
assign rld = ~RLD;  //complement 
assign qle = ~QLE;  //complement 
assign qld = ~QLD;  //complement 
assign qlk = ~QLK;  //complement 
assign qln = ~QLN;  //complement 
assign qlo = ~QLO;  //complement 
assign qla = ~QLA;  //complement 
assign qlb = ~QLB;  //complement 
assign qlc = ~QLC;  //complement 
assign qll = ~QLL;  //complement 
assign jqa =  qln & qqm & qqk  ; 
assign JQA = ~jqa;  //complement 
assign JQB =  qql & qlp & qqw  ; 
assign jqb = ~JQB;  //complement 
assign jjg =  qln & qqw  ; 
assign JJG = ~jjg;  //complement 
assign qlg = ~QLG;  //complement 
assign qli = ~QLI;  //complement 
assign GAD = ~gad;  //complement 
assign GAL = ~gal;  //complement 
assign FAD =  ebp & eao & ean & eam  ; 
assign fad = ~FAD;  //complement  
assign FAL =  eal & EAK & EAJ  ; 
assign fal = ~FAL;  //complement 
assign GBD = ~gbd;  //complement 
assign FBD =  EBL & EBK  ; 
assign fbd = ~FBD;  //complement  
assign GCD = ~gcd;  //complement 
assign GCL = ~gcl;  //complement 
assign QNQ = ~qnq;  //complement 
assign QNU = ~qnu;  //complement 
assign rka = ~RKA;  //complement 
assign qlj = ~QLJ;  //complement 
assign QNR = ~qnr;  //complement 
assign QNV = ~qnv;  //complement 
assign nad = ~NAD;  //complement 
assign rla = ~RLA;  //complement 
assign qea = ~QEA;  //complement 
assign qeb = ~QEB;  //complement 
assign qlm = ~QLM;  //complement 
assign JJB =  RBG & qcc  |  RJK  ; 
assign jjb = ~JJB;  //complement 
assign qrb = ~QRB;  //complement 
assign qrc = ~QRC;  //complement 
assign qrd = ~QRD;  //complement 
assign qre = ~QRE;  //complement 
assign qlp = ~QLP;  //complement 
assign qlq = ~QLQ;  //complement 
assign jrd =  qia & qib & qic  ; 
assign JRD = ~jrd;  //complement 
assign JCO =  RAG & QKJ  ; 
assign jco = ~JCO;  //complement 
assign jjk =  rlc  ; 
assign JJK = ~jjk;  //complement 
assign jre =  qlq & qsi  ; 
assign JRE = ~jre;  //complement 
assign qlf = ~QLF;  //complement 
assign lbd = ~LBD;  //complement 
assign JLD =  QLE & lba & lbb & lbc  ; 
assign jld = ~JLD;  //complement  
assign EAD = ~ead;  //complement 
assign WAD =  AAD & QXA  ; 
assign wad = ~WAD;  //complement 
assign WAL =  BAL & qxa  |  AAL & QXA  ; 
assign wal = ~WAL;  //complement 
assign aad = ~AAD;  //complement 
assign ohb = ~OHB;  //complement 
assign oad = ~OAD;  //complement 
assign oal = ~OAL;  //complement 
assign EAL = ~eal;  //complement 
assign EBL = ~ebl;  //complement 
assign ECL = ~ecl;  //complement 
assign dad = ~DAD;  //complement 
assign dal = ~DAL;  //complement 
assign edd = ~EDD;  //complement 
assign edl = ~EDL;  //complement 
assign aal = ~AAL;  //complement 
assign ogf = ~OGF;  //complement 
assign wcd = aad; 
assign WCD = ~wcd; //complement 
assign wcl = aal; 
assign WCL = ~wcl;  //complement 
assign wdd = abd; 
assign WDD = ~wdd;  //complement 
assign wdl = abl; 
assign WDL = ~wdl;  //complement 
assign tda = QXF; 
assign TDA = ~tda; //complement 
assign tdb = QXF; 
assign TDB = ~tdb;  //complement 
assign tdc = QXF; 
assign TDC = ~tdc;  //complement 
assign tdd = QXF; 
assign TDD = ~tdd;  //complement 
assign dbd = ~DBD;  //complement 
assign dbl = ~DBL;  //complement 
assign abd = ~ABD;  //complement 
assign ogn = ~OGN;  //complement 
assign ORD = ~ord;  //complement 
assign mab = ~MAB;  //complement 
assign WBD =  BBD & qxb  |  ABD & QXB  ; 
assign wbd = ~WBD;  //complement 
assign WBL =  BBL & qxb  |  ABL & QXB  ; 
assign wbl = ~WBL;  //complement 
assign abl = ~ABL;  //complement 
assign ogv = ~OGV;  //complement 
assign obd = ~OBD;  //complement 
assign obl = ~OBL;  //complement 
assign tea = qea; 
assign TEA = ~tea; //complement 
assign teb = qea; 
assign TEB = ~teb;  //complement 
assign tec = qeb; 
assign TEC = ~tec;  //complement 
assign ted = qeb; 
assign TED = ~ted;  //complement 
assign qlr = ~QLR;  //complement 
assign qls = ~QLS;  //complement 
assign olf = ~OLF;  //complement 
assign qfb = ~QFB;  //complement 
assign OCD = ~ocd;  //complement 
assign OCL = ~ocl;  //complement 
assign ODD = ~odd;  //complement 
assign ODL = ~odl;  //complement 
assign qca = ~QCA;  //complement 
assign qcc = ~QCC;  //complement 
assign qrf = ~QRF;  //complement 
assign rix = ~RIX;  //complement 
assign qra = ~QRA;  //complement 
assign ojc = ~OJC;  //complement 
assign oma = ~OMA;  //complement 
assign omb = ~OMB;  //complement 
assign jkc =  qlg & qli  ; 
assign JKC = ~jkc;  //complement  
assign jra =  qia & qib & qic & qid  ; 
assign JRA = ~jra;  //complement 
assign otc = ~OTC;  //complement 
assign QIB = ~qib;  //complement 
assign QIC = ~qic;  //complement 
assign QID = ~qid;  //complement 
assign QIA = ~qia;  //complement 
assign oed = ~OED;  //complement 
assign OEI = ~oei;  //complement 
assign kad = ~KAD;  //complement 
assign oje = ~OJE;  //complement 
assign reb = ~REB;  //complement 
assign ojd = ~OJD;  //complement 
assign lad = ~LAD;  //complement 
assign pae = ~PAE;  //complement 
assign pce = ~PCE;  //complement 
assign pee = ~PEE;  //complement 
assign JGE =  QVC  ; 
assign jge = ~JGE;  //complement  
assign JGM =  QVE  ; 
assign jgm = ~JGM;  //complement 
assign JDM =  QWE  ; 
assign jdm = ~JDM;  //complement  
assign pam = ~PAM;  //complement 
assign pcm = ~PCM;  //complement 
assign pem = ~PEM;  //complement 
assign QVC = ~qvc;  //complement 
assign bam = ~BAM;  //complement 
assign bcm = ~BCM;  //complement 
assign bem = ~BEM;  //complement 
assign QWE = ~qwe;  //complement 
assign pbe = ~PBE;  //complement 
assign pde = ~PDE;  //complement 
assign pfe = ~PFE;  //complement 
assign quf = ~QUF;  //complement 
assign bbe = ~BBE;  //complement 
assign bde = ~BDE;  //complement 
assign bfe = ~BFE;  //complement 
assign pbm = ~PBM;  //complement 
assign pdm = ~PDM;  //complement 
assign pfm = ~PFM;  //complement 
assign JHE =  QVF & QVH  ; 
assign jhe = ~JHE;  //complement  
assign JHM =  QVG & QVJ  ; 
assign jhm = ~JHM;  //complement 
assign bbm = ~BBM;  //complement 
assign bdm = ~BDM;  //complement 
assign bfm = ~BFM;  //complement 
assign JEE =  QWG  ; 
assign jee = ~JEE;  //complement  
assign JEM =  QWH & QWI  ; 
assign jem = ~JEM;  //complement 
assign GAE = ~gae;  //complement 
assign GAM = ~gam;  //complement 
assign FAE =  eap & EAO & ean & eam  ; 
assign fae = ~FAE;  //complement  
assign GBE = ~gbe;  //complement 
assign GBM = ~gbm;  //complement 
assign FBE =  EBL  ; 
assign fbe = ~FBE;  //complement  
assign GCM = ~gcm;  //complement 
assign QMA = ~qma;  //complement 
assign QME = ~qme;  //complement 
assign tld =  qma & qne  ; 
assign TLD = ~tld;  //complement 
assign QMB = ~qmb;  //complement 
assign QMC = ~qmc;  //complement 
assign QMF = ~qmf;  //complement 
assign QMG = ~qmg;  //complement 
assign rjk = ~RJK;  //complement 
assign rja = ~RJA;  //complement 
assign rje = ~RJE;  //complement 
assign rjb = ~RJB;  //complement 
assign rjc = ~RJC;  //complement 
assign rjd = ~RJD;  //complement 
assign rjl = ~RJL;  //complement 
assign raa = ~RAA;  //complement 
assign raf = ~RAF;  //complement 
assign rag = ~RAG;  //complement 
assign JCM =  RAG & qkg  ; 
assign jcm = ~JCM;  //complement 
assign JCP =  RAG & QKJ  ; 
assign jcp = ~JCP;  //complement 
assign JJC =  RBG  ; 
assign jjc = ~JJC;  //complement 
assign lbe = ~LBE;  //complement 
assign JLE =  QLE & lba & lbb & lbc & lbd  ; 
assign jle = ~JLE;  //complement  
assign EAE = ~eae;  //complement 
assign WAE =  AAE & QXA  ; 
assign wae = ~WAE;  //complement 
assign WAM =  BAM & qxa  |  AAM & QXA  ; 
assign wam = ~WAM;  //complement 
assign aae = ~AAE;  //complement 
assign ohc = ~OHC;  //complement 
assign oae = ~OAE;  //complement 
assign oam = ~OAM;  //complement 
assign EAM = ~eam;  //complement 
assign ECM = ~ecm;  //complement 
assign dae = ~DAE;  //complement 
assign dam = ~DAM;  //complement 
assign ede = ~EDE;  //complement 
assign edm = ~EDM;  //complement 
assign GBF = ~gbf;  //complement 
assign GBN = ~gbn;  //complement 
assign wce = aae; 
assign WCE = ~wce; //complement 
assign wcm = aam; 
assign WCM = ~wcm;  //complement 
assign wde = abe; 
assign WDE = ~wde;  //complement 
assign wdm = abm; 
assign WDM = ~wdm;  //complement 
assign qxa = ~QXA;  //complement 
assign qxb = ~QXB;  //complement 
assign dbe = ~DBE;  //complement 
assign dbm = ~DBM;  //complement 
assign abe = ~ABE;  //complement 
assign ogo = ~OGO;  //complement 
assign ORE = ~ore;  //complement 
assign mac = ~MAC;  //complement 
assign WBE =  BBE & qxb  |  ABE & QXB  ; 
assign wbe = ~WBE;  //complement 
assign WBM =  BBM & qxb  |  ABM & QXB  ; 
assign wbm = ~WBM;  //complement 
assign abm = ~ABM;  //complement 
assign ogw = ~OGW;  //complement 
assign obe = ~OBE;  //complement 
assign obm = ~OBM;  //complement 
assign rjf = ~RJF;  //complement 
assign rjg = ~RJG;  //complement 
assign rjh = ~RJH;  //complement 
assign rji = ~RJI;  //complement 
assign jcd =  rja & rjb & rjc & raa & rab  ; 
assign JCD = ~jcd;  //complement  
assign oia = ~OIA;  //complement 
assign rec = ~REC;  //complement 
assign OCE = ~oce;  //complement 
assign OCM = ~ocm;  //complement 
assign ODE = ~ode;  //complement 
assign ODM = ~odm;  //complement 
assign rab = ~RAB;  //complement 
assign rac = ~RAC;  //complement 
assign rad = ~RAD;  //complement 
assign rae = ~RAE;  //complement 
assign jca =  raa & rab & rac & rad & rae & raf  ; 
assign JCA = ~jca;  //complement  
assign jce =  raa & rja  ; 
assign JCE = ~jce;  //complement 
assign oic = ~OIC;  //complement 
assign oib = ~OIB;  //complement 
assign oid = ~OID;  //complement 
assign jcc =  rag & rbg  ; 
assign JCC = ~jcc;  //complement 
assign JCR =  RQB  ; 
assign jcr = ~JCR;  //complement 
assign oee = ~OEE;  //complement 
assign oie = ~OIE;  //complement 
assign olc = ~OLC;  //complement 
assign ota = ~OTA;  //complement 
assign kae = ~KAE;  //complement 
assign OTD = ~otd;  //complement 
assign lae = ~LAE;  //complement 
assign paf = ~PAF;  //complement 
assign pcf = ~PCF;  //complement 
assign pef = ~PEF;  //complement 
assign JGF =  QVC & PCE  ; 
assign jgf = ~JGF;  //complement  
assign JGN =  QVE & PCM  ; 
assign jgn = ~JGN;  //complement 
assign JDN =  QWE & BCM  ; 
assign jdn = ~JDN;  //complement  
assign pan = ~PAN;  //complement 
assign pcn = ~PCN;  //complement 
assign pen = ~PEN;  //complement 
assign QVD = ~qvd;  //complement 
assign ban = ~BAN;  //complement 
assign bcn = ~BCN;  //complement 
assign ben = ~BEN;  //complement 
assign QWF = ~qwf;  //complement 
assign pbf = ~PBF;  //complement 
assign pdf = ~PDF;  //complement 
assign pff = ~PFF;  //complement 
assign tpc = qwj; 
assign TPC = ~tpc; //complement 
assign tpd = qwj; 
assign TPD = ~tpd;  //complement 
assign bbf = ~BBF;  //complement 
assign bdf = ~BDF;  //complement 
assign bff = ~BFF;  //complement 
assign tfc = qwa; 
assign TFC = ~tfc; //complement 
assign tfd = qwa; 
assign TFD = ~tfd;  //complement 
assign pbn = ~PBN;  //complement 
assign pdn = ~PDN;  //complement 
assign pfn = ~PFN;  //complement 
assign JHF =  QVF & QVH & PDE  ; 
assign jhf = ~JHF;  //complement  
assign JHN =  QVG & QVJ & PDM  ; 
assign jhn = ~JHN;  //complement 
assign bbn = ~BBN;  //complement 
assign bdn = ~BDN;  //complement 
assign bfn = ~BFN;  //complement 
assign JEF =  QWG & BDE  ; 
assign jef = ~JEF;  //complement  
assign JEN =  QWH & QWI & BDM  ; 
assign jen = ~JEN;  //complement 
assign qql = ~QQL;  //complement 
assign RQA = ~rqa;  //complement 
assign qqm = ~QQM;  //complement 
assign qqi = ~QQI;  //complement 
assign JQC =  qql & qlp  ; 
assign jqc = ~JQC;  //complement 
assign JJL =  QQL  ; 
assign jjl = ~JJL;  //complement 
assign jjm =  qln  ; 
assign JJM = ~jjm;  //complement 
assign qqn = ~QQN;  //complement 
assign rqb = ~RQB;  //complement 
assign RQC = ~rqc;  //complement 
assign GAN = ~gan;  //complement 
assign GAF = ~gaf;  //complement 
assign FAF =  eap & EAO & ean & EAM  ; 
assign faf = ~FAF;  //complement  
assign aam = ~AAM;  //complement 
assign ogg = ~OGG;  //complement 
assign GCN = ~gcn;  //complement 
assign qmk = ~QMK;  //complement 
assign QMI = ~qmi;  //complement 
assign TCE = QXE; 
assign tce = ~TCE; //complement 
assign TCF = QXE; 
assign tcf = ~TCF;  //complement 
assign TCG = QXE; 
assign tcg = ~TCG;  //complement 
assign TCH = QXE; 
assign tch = ~TCH;  //complement 
assign JJN =  QQL  ; 
assign jjn = ~JJN;  //complement  
assign jfh =  gbm & gbn  ; 
assign JFH = ~jfh;  //complement 
assign QMJ = ~qmj;  //complement 
assign QQX = ~qqx;  //complement 
assign JJP =  QQL & QQC  ; 
assign jjp = ~JJP;  //complement 
assign JQE =  QQA & qqb  ; 
assign jqe = ~JQE;  //complement 
assign jcb =  rba & rbb & rbc & rbd & rbe & rbf  ; 
assign JCB = ~jcb;  //complement  
assign JJH =  QQC  ; 
assign jjh = ~JJH;  //complement 
assign qqh = ~QQH;  //complement 
assign JCS = RQC; 
assign jcs = ~JCS; //complement 
assign JJE = QQE; 
assign jje = ~JJE;  //complement 
assign JJF = QQE; 
assign jjf = ~JJF;  //complement 
assign JQD = QQA; 
assign jqd = ~JQD;  //complement 
assign jcf =  reb & qqa & qqc & qka & qta & qtx  ; 
assign JCF = ~jcf;  //complement  
assign JTB =  qqa & qlq & qtw & qqb  ; 
assign jtb = ~JTB;  //complement 
assign qqj = ~QQJ;  //complement 
assign qqd = ~QQD;  //complement 
assign qqe = ~QQE;  //complement 
assign qqf = ~QQF;  //complement 
assign qqg = ~QQG;  //complement 
assign JCG =  RAG & qkj  ; 
assign jcg = ~JCG;  //complement 
assign JCQ =  RAG & QKJ  ; 
assign jcq = ~JCQ;  //complement 
assign JJD =  RBG  ; 
assign jjd = ~JJD;  //complement 
assign qqk = ~QQK;  //complement 
assign lbf = ~LBF;  //complement 
assign JLF =  QLE & lba & lbb & lbc & lbd & lbe  ; 
assign jlf = ~JLF;  //complement  
assign EAF = ~eaf;  //complement 
assign WAF =  AAF & QXC  ; 
assign waf = ~WAF;  //complement 
assign WAN =  BAN & qxc  |  AAN & QXC  ; 
assign wan = ~WAN;  //complement 
assign aaf = ~AAF;  //complement 
assign ohd = ~OHD;  //complement 
assign oaf = ~OAF;  //complement 
assign oan = ~OAN;  //complement 
assign EAN = ~ean;  //complement 
assign ECN = ~ecn;  //complement 
assign daf = ~DAF;  //complement 
assign dan = ~DAN;  //complement 
assign edf = ~EDF;  //complement 
assign edn = ~EDN;  //complement 
assign aan = ~AAN;  //complement 
assign ogh = ~OGH;  //complement 
assign wcf = aaf; 
assign WCF = ~wcf; //complement 
assign wcn = aan; 
assign WCN = ~wcn;  //complement 
assign wdf = abf; 
assign WDF = ~wdf;  //complement 
assign wdn = abn; 
assign WDN = ~wdn;  //complement 
assign qxc = ~QXC;  //complement 
assign qxd = ~QXD;  //complement 
assign dbf = ~DBF;  //complement 
assign dbn = ~DBN;  //complement 
assign abf = ~ABF;  //complement 
assign ogp = ~OGP;  //complement 
assign ORF = ~orf;  //complement 
assign JJI = QQC; 
assign jji = ~JJI; //complement 
assign JJJ = QQC; 
assign jjj = ~JJJ;  //complement 
assign TEE = QQX; 
assign tee = ~TEE;  //complement 
assign TEF = QQX; 
assign tef = ~TEF;  //complement 
assign WBF =  BBF & qxd  |  ABF & QXD  ; 
assign wbf = ~WBF;  //complement 
assign WBN =  BBN & qxd  |  ABN & QXD  ; 
assign wbn = ~WBN;  //complement 
assign abn = ~ABN;  //complement 
assign ogx = ~OGX;  //complement 
assign obf = ~OBF;  //complement 
assign obn = ~OBN;  //complement 
assign rbf = ~RBF;  //complement 
assign rbg = ~RBG;  //complement 
assign rbb = ~RBB;  //complement 
assign rbc = ~RBC;  //complement 
assign rbd = ~RBD;  //complement 
assign rbe = ~RBE;  //complement 
assign RBA = ~rba;  //complement 
assign OCF = ~ocf;  //complement 
assign OCN = ~ocn;  //complement 
assign ODF = ~odf;  //complement 
assign ODN = ~odn;  //complement 
assign qqc = ~QQC;  //complement 
assign qhe = ~QHE;  //complement 
assign qhf = ~QHF;  //complement 
assign QTQ = ~qtq;  //complement 
assign QTR = ~qtr;  //complement 
assign qhc = ~QHC;  //complement 
assign oej = ~OEJ;  //complement 
assign qhd = ~QHD;  //complement 
assign qqa = ~QQA;  //complement 
assign qqb = ~QQB;  //complement 
assign qqw = ~QQW;  //complement 
assign oem = ~OEM;  //complement 
assign oef = ~OEF;  //complement 
assign OTE = ~ote;  //complement 
assign kaf = ~KAF;  //complement 
assign oep = ~OEP;  //complement 
assign laf = ~LAF;  //complement 
assign pag = ~PAG;  //complement 
assign pcg = ~PCG;  //complement 
assign peg = ~PEG;  //complement 
assign JGG =  QVC & PCE & PCF  ; 
assign jgg = ~JGG;  //complement  
assign JGO =  QVE & PCM & PCN  ; 
assign jgo = ~JGO;  //complement 
assign bag = ~BAG;  //complement 
assign bcg = ~BCG;  //complement 
assign beg = ~BEG;  //complement 
assign JDG =  QWC  ; 
assign jdg = ~JDG;  //complement  
assign JDO =  QWE & BCM & BCN  ; 
assign jdo = ~JDO;  //complement 
assign pao = ~PAO;  //complement 
assign pco = ~PCO;  //complement 
assign peo = ~PEO;  //complement 
assign QVE = ~qve;  //complement 
assign bao = ~BAO;  //complement 
assign bco = ~BCO;  //complement 
assign beo = ~BEO;  //complement 
assign QWG = ~qwg;  //complement 
assign pbg = ~PBG;  //complement 
assign pdg = ~PDG;  //complement 
assign pfg = ~PFG;  //complement 
assign JFB =  PEE & PEF & PEG & PEH  ; 
assign jfb = ~JFB;  //complement  
assign JFD =  PEM & PEN & PEO & PEP  ; 
assign jfd = ~JFD;  //complement 
assign bbg = ~BBG;  //complement 
assign bdg = ~BDG;  //complement 
assign bfg = ~BFG;  //complement 
assign JDA =  BEG & BEH & QWB  ; 
assign jda = ~JDA;  //complement  
assign pbo = ~PBO;  //complement 
assign pdo = ~PDO;  //complement 
assign pfo = ~PFO;  //complement 
assign JHG =  QVF & QVH & PDE & PDF  ; 
assign jhg = ~JHG;  //complement  
assign JHO =  QVG & QVJ & PDM & PDN  ; 
assign jho = ~JHO;  //complement 
assign bbo = ~BBO;  //complement 
assign bdo = ~BDO;  //complement 
assign bfo = ~BFO;  //complement 
assign JEG =  QWG & BDE & BDF  ; 
assign jeg = ~JEG;  //complement  
assign JEO =  QWH & QWI & BDM & BDN  ; 
assign jeo = ~JEO;  //complement 
assign GAG = ~gag;  //complement 
assign GAO = ~gao;  //complement 
assign FAG =  eap & EAO & EAN & eam  ; 
assign fag = ~FAG;  //complement  
assign GBG = ~gbg;  //complement 
assign GBO = ~gbo;  //complement 
assign FBG =  EBJ  ; 
assign fbg = ~FBG;  //complement  
assign QNA = ~qna;  //complement 
assign QNE = ~qne;  //complement 
assign JCI =  GAN & gal  ; 
assign jci = ~JCI;  //complement  
assign jcj =  gbm & gbo  ; 
assign JCJ = ~jcj;  //complement 
assign QNB = ~qnb;  //complement 
assign QNC = ~qnc;  //complement 
assign QNF = ~qnf;  //complement 
assign QNG = ~qng;  //complement 
assign jch =  qqa & qqb & qqn & qta & qtx  ; 
assign JCH = ~jch;  //complement  
assign jke =  qnj & qnr & qnv  ; 
assign JKE = ~jke;  //complement 
assign tha =  rqb  ; 
assign THA = ~tha;  //complement 
assign JLG =  LBA & lbb & lbc & lbd & lbe & lbf  ; 
assign jlg = ~JLG;  //complement  
assign EAG = ~eag;  //complement 
assign WAG =  BAG & qxc  |  AAG & QXC  ; 
assign wag = ~WAG;  //complement 
assign WAO =  BAO & qxc  |  AAO & QXC  ; 
assign wao = ~WAO;  //complement 
assign aag = ~AAG;  //complement 
assign oga = ~OGA;  //complement 
assign oag = ~OAG;  //complement 
assign oao = ~OAO;  //complement 
assign EAO = ~eao;  //complement 
assign ECO = ~eco;  //complement 
assign dag = ~DAG;  //complement 
assign dao = ~DAO;  //complement 
assign edg = ~EDG;  //complement 
assign edo = ~EDO;  //complement 
assign aao = ~AAO;  //complement 
assign ogi = ~OGI;  //complement 
assign wcg = aag; 
assign WCG = ~wcg; //complement 
assign wco = aao; 
assign WCO = ~wco;  //complement 
assign wdg = abg; 
assign WDG = ~wdg;  //complement 
assign wdo = abo; 
assign WDO = ~wdo;  //complement 
assign tde = QXF; 
assign TDE = ~tde; //complement 
assign tdf = QXF; 
assign TDF = ~tdf;  //complement 
assign tdg = QXF; 
assign TDG = ~tdg;  //complement 
assign tdh = QXF; 
assign TDH = ~tdh;  //complement 
assign dbg = ~DBG;  //complement 
assign dbo = ~DBO;  //complement 
assign abg = ~ABG;  //complement 
assign ogq = ~OGQ;  //complement 
assign QSI = ~qsi;  //complement 
assign TAE = RJL; 
assign tae = ~TAE; //complement 
assign TAF = RJL; 
assign taf = ~TAF;  //complement 
assign TAG = RJL; 
assign tag = ~TAG;  //complement 
assign TAH = RJL; 
assign tah = ~TAH;  //complement 
assign WBG =  BBG & qxd  |  ABG & QXD  ; 
assign wbg = ~WBG;  //complement 
assign WBO =  BBO & qxd  |  ABO & QXD  ; 
assign wbo = ~WBO;  //complement 
assign abo = ~ABO;  //complement 
assign obg = ~OBG;  //complement 
assign obo = ~OBO;  //complement 
assign JQF =  QQB & qtp  ; 
assign jqf = ~JQF;  //complement 
assign OLD = ~old;  //complement 
assign OCG = ~ocg;  //complement 
assign OCO = ~oco;  //complement 
assign ODG = ~odg;  //complement 
assign ODO = ~odo;  //complement 
assign JXA =  QLN & QSD  ; 
assign jxa = ~JXA;  //complement 
assign oes = ~OES;  //complement 
assign ofc = ~OFC;  //complement 
assign olb = ~OLB;  //complement 
assign oqb = ~OQB;  //complement 
assign OTF = ~otf;  //complement 
assign oet = ~OET;  //complement 
assign oeh = ~OEH;  //complement 
assign oeq = ~OEQ;  //complement 
assign OER = ~oer;  //complement 
assign ofa = ~OFA;  //complement 
assign ola = ~OLA;  //complement 
assign OFB = ~ofb;  //complement 
assign OQA = ~oqa;  //complement 
assign pah = ~PAH;  //complement 
assign pch = ~PCH;  //complement 
assign peh = ~PEH;  //complement 
assign JGH =  QVC & PCE & PCF & PCG  ; 
assign jgh = ~JGH;  //complement  
assign JGP =  QVE & PCM & PCN & PCO  ; 
assign jgp = ~JGP;  //complement 
assign bah = ~BAH;  //complement 
assign bch = ~BCH;  //complement 
assign beh = ~BEH;  //complement 
assign JDH =  QWC & BCG  ; 
assign jdh = ~JDH;  //complement  
assign JDP =  QWE & BCM & BCN & BCO  ; 
assign jdp = ~JDP;  //complement 
assign pap = ~PAP;  //complement 
assign pcp = ~PCP;  //complement 
assign pep = ~PEP;  //complement 
assign QVF = ~qvf;  //complement 
assign QVG = ~qvg;  //complement 
assign bap = ~BAP;  //complement 
assign bcp = ~BCP;  //complement 
assign bep = ~BEP;  //complement 
assign QWH = ~qwh;  //complement 
assign pbh = ~PBH;  //complement 
assign pdh = ~PDH;  //complement 
assign pfh = ~PFH;  //complement 
assign JHH =  QVF & QVH & PDE & PDF & PDG  ; 
assign jhh = ~JHH;  //complement  
assign JFF =  PFE & PFF & PFG & PFH  ; 
assign jff = ~JFF;  //complement 
assign bbh = ~BBH;  //complement 
assign bdh = ~BDH;  //complement 
assign bfh = ~BFH;  //complement 
assign JDC =  BEM & BEN & BEO & BEP  ; 
assign jdc = ~JDC;  //complement  
assign JDE =  BFE & BFF & BFG & BFH  ; 
assign jde = ~JDE;  //complement 
assign pbp = ~PBP;  //complement 
assign pdp = ~PDP;  //complement 
assign pfp = ~PFP;  //complement 
assign JHP =  QVG & QVJ & PDM & PDN & PDO  ; 
assign jhp = ~JHP;  //complement  
assign bbp = ~BBP;  //complement 
assign bdp = ~BDP;  //complement 
assign bfp = ~BFP;  //complement 
assign JEH =  QWG & BDE & BDF & BDG  ; 
assign jeh = ~JEH;  //complement  
assign GAH = ~gah;  //complement 
assign GAP = ~gap;  //complement 
assign FAH =  eap & EAO & EAN & EAM  ; 
assign fah = ~FAH;  //complement  
assign FAP =  EAL & EAK & EAJ  ; 
assign fap = ~FAP;  //complement 
assign GBH = ~gbh;  //complement 
assign GBP = ~gbp;  //complement 
assign FBH =  EBK  ; 
assign fbh = ~FBH;  //complement  
assign GCH = ~gch;  //complement 
assign tga = qba; 
assign TGA = ~tga; //complement 
assign tgb = qba; 
assign TGB = ~tgb;  //complement 
assign tgc = qba; 
assign TGC = ~tgc;  //complement 
assign tgd = qba; 
assign TGD = ~tgd;  //complement 
assign JEP =  QWH & QWI & BDM & BDN & BDO  ; 
assign jep = ~JEP;  //complement  
assign jck =  gbm & gbn & gbp  ; 
assign JCK = ~jck;  //complement  
assign jcl =  gbm & gbn & gbo & gbp  ; 
assign JCL = ~jcl;  //complement 
assign JXB =  QSC & qlq & qqa  ; 
assign jxb = ~JXB;  //complement 
assign qsc = ~QSC;  //complement 
assign qsd = ~QSD;  //complement 
assign rsa = ~RSA;  //complement 
assign rsb = ~RSB;  //complement 
assign rsc = ~RSC;  //complement 
assign qse = ~QSE;  //complement 
assign qsf = ~QSF;  //complement 
assign qsg = ~QSG;  //complement 
assign tla =  qma & rsb & rqc  ; 
assign TLA = ~tla;  //complement 
assign tlb =  rsa  ; 
assign TLB = ~tlb;  //complement 
assign tlc =  qmc & qnc & rsc & rqc  ; 
assign TLC = ~tlc;  //complement  
assign EAH = ~eah;  //complement 
assign WAH =  BAH & qxc  |  AAH & QXC  ; 
assign wah = ~WAH;  //complement 
assign WAP =  BAP & qxc  |  AAP & QXC  ; 
assign wap = ~WAP;  //complement 
assign aah = ~AAH;  //complement 
assign ogb = ~OGB;  //complement 
assign oah = ~OAH;  //complement 
assign oap = ~OAP;  //complement 
assign EAP = ~eap;  //complement 
assign EBP = ~ebp;  //complement 
assign ECP = ~ecp;  //complement 
assign dah = ~DAH;  //complement 
assign dap = ~DAP;  //complement 
assign edh = ~EDH;  //complement 
assign edp = ~EDP;  //complement 
assign aap = ~AAP;  //complement 
assign ogj = ~OGJ;  //complement 
assign wch = aah; 
assign WCH = ~wch; //complement 
assign wcp = aap; 
assign WCP = ~wcp;  //complement 
assign wdh = abh; 
assign WDH = ~wdh;  //complement 
assign wdp = abp; 
assign WDP = ~wdp;  //complement 
assign TGE = QBA; 
assign tge = ~TGE; //complement 
assign TGF = QBA; 
assign tgf = ~TGF;  //complement 
assign dbh = ~DBH;  //complement 
assign dbp = ~DBP;  //complement 
assign qba = ~QBA;  //complement 
assign abh = ~ABH;  //complement 
assign ogr = ~OGR;  //complement 
assign jkd =  qmj & qnm & qnq & qnj  ; 
assign JKD = ~jkd;  //complement  
assign WBH =  BBH & qxd  |  ABH & QXD  ; 
assign wbh = ~WBH;  //complement 
assign WBP =  BBP & qxd  |  ABP & QXD  ; 
assign wbp = ~WBP;  //complement 
assign abp = ~ABP;  //complement 
assign obh = ~OBH;  //complement 
assign obp = ~OBP;  //complement 
assign qsb = ~QSB;  //complement 
assign qsa = ~QSA;  //complement 
assign qaa = ~QAA;  //complement 
assign qab = ~QAB;  //complement 
assign qac = ~QAC;  //complement 
assign qad = ~QAD;  //complement 
assign OCH = ~och;  //complement 
assign OCP = ~ocp;  //complement 
assign ODH = ~odh;  //complement 
assign ODP = ~odp;  //complement 
assign rre = ~RRE;  //complement 
assign rrf = ~RRF;  //complement 
assign rrg = ~RRG;  //complement 
assign rrh = ~RRH;  //complement 
assign rra = ~RRA;  //complement 
assign rrb = ~RRB;  //complement 
assign rrc = ~RRC;  //complement 
assign rrd = ~RRD;  //complement 
assign oeg = ~OEG;  //complement 
assign QFC = ~qfc;  //complement 
assign qsh = ~QSH;  //complement 
assign oel = ~OEL;  //complement 
assign oev = ~OEV;  //complement 
assign oen = ~OEN;  //complement 
assign oeo = ~OEO;  //complement 
assign oex = ~OEX;  //complement 
assign oey = ~OEY;  //complement 
assign oek = ~OEK;  //complement 
assign oeu = ~OEU;  //complement 
assign oew = ~OEW;  //complement 
assign iaa = ~IAA; //complement 
assign iab = ~IAB; //complement 
assign iac = ~IAC; //complement 
assign iad = ~IAD; //complement 
assign iae = ~IAE; //complement 
assign iaf = ~IAF; //complement 
assign iag = ~IAG; //complement 
assign iah = ~IAH; //complement 
assign iai = ~IAI; //complement 
assign iaj = ~IAJ; //complement 
assign iak = ~IAK; //complement 
assign ial = ~IAL; //complement 
assign iam = ~IAM; //complement 
assign iba = ~IBA; //complement 
assign ibb = ~IBB; //complement 
assign ibc = ~IBC; //complement 
assign ibd = ~IBD; //complement 
assign ibe = ~IBE; //complement 
assign ibf = ~IBF; //complement 
assign ibg = ~IBG; //complement 
assign ibh = ~IBH; //complement 
assign ibi = ~IBI; //complement 
assign ibj = ~IBJ; //complement 
assign ibk = ~IBK; //complement 
assign ibl = ~IBL; //complement 
assign ibm = ~IBM; //complement 
assign ica = ~ICA; //complement 
assign icb = ~ICB; //complement 
assign icc = ~ICC; //complement 
assign icd = ~ICD; //complement 
assign ice = ~ICE; //complement 
assign icf = ~ICF; //complement 
assign icg = ~ICG; //complement 
assign ich = ~ICH; //complement 
assign ici = ~ICI; //complement 
assign icj = ~ICJ; //complement 
assign ick = ~ICK; //complement 
assign icl = ~ICL; //complement 
assign icm = ~ICM; //complement 
assign icn = ~ICN; //complement 
assign ico = ~ICO; //complement 
assign icp = ~ICP; //complement 
assign ida = ~IDA; //complement 
assign idb = ~IDB; //complement 
assign idc = ~IDC; //complement 
assign idd = ~IDD; //complement 
assign ide = ~IDE; //complement 
assign idf = ~IDF; //complement 
assign idg = ~IDG; //complement 
assign idh = ~IDH; //complement 
assign idi = ~IDI; //complement 
assign idj = ~IDJ; //complement 
assign idk = ~IDK; //complement 
assign idl = ~IDL; //complement 
assign idm = ~IDM; //complement 
assign idn = ~IDN; //complement 
assign ido = ~IDO; //complement 
assign idp = ~IDP; //complement 
assign iea = ~IEA; //complement 
assign ieb = ~IEB; //complement 
assign iec = ~IEC; //complement 
assign ied = ~IED; //complement 
assign iee = ~IEE; //complement 
assign ief = ~IEF; //complement 
assign ieg = ~IEG; //complement 
assign ieh = ~IEH; //complement 
assign iei = ~IEI; //complement 
assign iej = ~IEJ; //complement 
assign iek = ~IEK; //complement 
assign iel = ~IEL; //complement 
assign iem = ~IEM; //complement 
assign ien = ~IEN; //complement 
assign ieo = ~IEO; //complement 
assign iep = ~IEP; //complement 
assign ifa = ~IFA; //complement 
assign ifb = ~IFB; //complement 
assign ifc = ~IFC; //complement 
assign ifd = ~IFD; //complement 
assign ife = ~IFE; //complement 
assign ifff  = ~IFFF ; //complement 
assign ifg = ~IFG; //complement 
assign ifh = ~IFH; //complement 
assign ifi = ~IFI; //complement 
assign iga = ~IGA; //complement 
assign igb = ~IGB; //complement 
assign igc = ~IGC; //complement 
assign iha = ~IHA; //complement 
assign ihb = ~IHB; //complement 
assign ihc = ~IHC; //complement 
assign ija = ~IJA; //complement 
assign ijb = ~IJB; //complement 
assign ijc = ~IJC; //complement 
assign ijd = ~IJD; //complement 
assign ika = ~IKA; //complement 
assign ikb = ~IKB; //complement 
assign ila = ~ILA; //complement 
assign ilb = ~ILB; //complement 
assign ilc = ~ILC; //complement 
assign ima = ~IMA; //complement 
assign imb = ~IMB; //complement 
assign imc = ~IMC; //complement 
assign imd = ~IMD; //complement 
assign ime = ~IME; //complement 
assign imf = ~IMF; //complement 
assign img = ~IMG; //complement 
assign ina = ~INA; //complement 
assign ioa = ~IOA; //complement 
assign iob = ~IOB; //complement 
assign ioc = ~IOC; //complement 
assign iod = ~IOD; //complement 
assign iog = ~IOG; //complement 
assign ipa = ~IPA; //complement 
assign ipb = ~IPB; //complement 
assign ipc = ~IPC; //complement 
assign ipd = ~IPD; //complement 
assign ipe = ~IPE; //complement 
assign ipf = ~IPF; //complement 
assign iqa = ~IQA; //complement 
assign iqb = ~IQB; //complement 
assign iqc = ~IQC; //complement 
assign iqd = ~IQD; //complement 
assign iqe = ~IQE; //complement 
assign iqf = ~IQF; //complement 
assign iqg = ~IQG; //complement 
assign iqh = ~IQH; //complement 
assign iqi = ~IQI; //complement 
always@(posedge IZZ )
   begin 
 PAA <=  PAA & jga & tpe  |  paa & JGA  |  AAA & TPE  ; 
 PCA <=  PAA & jga & tpe  |  paa & JGA  |  AAA & TPE  ; 
 PEA <=  PAA & jga & tpe  |  paa & JGA  |  AAA & TPE  ; 
 PAI <=  PAI & jgi & tpb  |  pai & JGI  |  AAI & TPB  ; 
 PCI <=  PAI & jgi & tpb  |  pai & JGI  |  AAI & TPB  ; 
 PEI <=  PAI & jgi & tpb  |  pai & JGI  |  AAI & TPB  ; 
 qva <=  qua  ; 
 qvj <=  jfe  |  jff  |  jfg  ; 
 BAI <=  BAI & jdi & tfb  |  bai & JDI  |  AAI & TFB  ; 
 BCI <=  BAI & jdi & tfb  |  bai & JDI  |  AAI & TFB  ; 
 BEI <=  BAI & jdi & tfb  |  bai & JDI  |  AAI & TFB  ; 
 PBA <=  PBA & jha & tpc  |  pba & JHA  |  ABA & TPC  ; 
 PDA <=  PBA & jha & tpc  |  pba & JHA  |  ABA & TPC  ; 
 PFA <=  PBA & jha & tpc  |  pba & JHA  |  ABA & TPC  ; 
 BBA <=  BBA & jea & tfc  |  bba & JEA  |  ABA & TFC  ; 
 BDA <=  BBA & jea & tfc  |  bba & JEA  |  ABA & TFC  ; 
 BFA <=  BBA & jea & tfc  |  bba & JEA  |  ABA & TFC  ; 
 PBI <=  PBI & jhi & tpd  |  pbi & JHA  |  ABI & TPD  ; 
 PDI <=  PBI & jhi & tpd  |  pbi & JHA  |  ABI & TPD  ; 
 PFI <=  PBI & jhi & tpd  |  pbi & JHA  |  ABI & TPD  ; 
 BBI <=  BBI & jei & tfd  |  bbi & JEI  |  ABI & TFD  ; 
 BDI <=  BBI & jei & tfd  |  bbi & JEI  |  ABI & TFD  ; 
 BFI <=  BBI & jei & tfd  |  bbi & JEI  |  ABI & TFD  ; 
 hba <= haa ; 
 hca <= hba ; 
 hda <= hca ; 
 hea <= hda ; 
 hbb <= hab ; 
 hcb <= hbb ; 
 hdb <= hcb ; 
 heb <= hdb ; 
 hbc <= hac ; 
 hcc <= hbc ; 
 hdc <= hcc ; 
 hec <= hdc ; 
 hbd <= had ; 
 hcd <= hbd ; 
 hdd <= hcd ; 
 hed <= hdd ; 
 hbe <= hae ; 
 hce <= hbe ; 
 hde <= hce ; 
 hee <= hde ; 
 hbf <= haf ; 
 hcf <= hbf ; 
 hdf <= hcf ; 
 hef <= hdf ; 
 hbg <= hag ; 
 hcg <= hbg ; 
 hdg <= hcg ; 
 heg <= hdg ; 
 hbh <= hah ; 
 hch <= hbh ; 
 hdh <= hch ; 
 heh <= hdh ; 
 hfa <= hea ; 
 hfb <= heb ; 
 hfc <= hec ; 
 hfd <= hed ; 
 hfh <= heh ; 
 gaa <=  fbg & TGA  |  gaa & tga  ; 
 gai <=  eai & TGA  |  gai & tga  ; 
 gba <=  faa & TGC  |  fak & TGD  |  gba & tgc  ; 
 gbi <=  fae & TGC  |  fbc & TGD  |  gbi & tgc  ; 
 qpa <=  qab  ; 
 qpb <=  qab  |  jfi  ; 
 gca <=  fag & TGE  |  fba & TGF  |  gca & tge  ; 
 gci <=  eaa & TGE  |  ZZO & TGF  |  gci & tge  ; 
 hae <=  gam  |  gad  ; 
 haf <=  gan  |  gad  ; 
 haa <=  GAB  |  GAA  ; 
 hab <=  GAB  |  gaa  ; 
 hac <=  gab  |  GAA  ; 
 had <=  gab  |  gaa  ; 
 QXE <=  GAC & QAA  ; 
 QXF <=  GAC & QAA  |  RJC  |  QYA  ; 
 NAA <=  NAA & jsa & tha  |  naa & JSA  |  WCC & THA  ; 
 NBA <=  NAA & jsa & tha  |  naa & JSA  |  WCC & THA  ; 
 QTW <=  JIC  |  JID  ; 
 QTX <=  QTX & rji  |  QTJ & JTB  |  QTN  ; 
 QTF <= QTE ; 
 QTG <= QTF ; 
 QTH <= QTG ; 
 QTI <= QTH ; 
 QND <=  QNC  ; 
 qoa <=  rld  |  QND  ; 
 LBA <=  LBA & jla & tla  |  lba & JLA  |  LAA & TLA  ; 
 eaa <=  iea  ; 
 AAA <=  IAA & TAA  |  DAA & TBA  |  IEA & TCA  |  WAA & TDA  |  TMA  ; 
 OAA <=  DAA & TEA  |  EAA & TEC  |  NAA & TEE  ; 
 OAI <=  DAI & TEA  |  ECI & TEC  |  WCK & TEE  ; 
 eai <=  iei  ; 
 eci <=  iei  ; 
 DAA <= ICA ; 
 DAI <= ICI ; 
 EDA <= EAA ; 
 EDI <= EAI ; 
 AAI <=  IAI & TAB  |  DAI & TBB  |  IEI & TCB  |  WAI & TDA  |  TMB  ; 
 OGC <=  IAI & TAB  |  DAI & TBB  |  IEI & TCB  |  WAI & TDA  |  TMB  ; 
 DBA <= IDA ; 
 DBI <= IDI ; 
 ABA <=  IBA & TAC  |  DBA & TBC  |  EAA & TCC  |  WBA & TDC  |  TMC  ; 
 OGK <=  IBA & TAC  |  DBA & TBC  |  EAA & TCC  |  WBA & TDC  |  TMC  ; 
 OTB <= QTW ; 
 ora <= gci ; 
 OGS <=  IBI & TAD  |  DBI & TBD  |  ECI & TCD  |  WBI & TDD  |  TMD  ; 
 ABI <=  IBI & TAD  |  DBI & TBD  |  ECI & TCD  |  WBI & TDD  |  TMD  ; 
 OBA <=  DBA & TEB  |  EDA & TED  |  WDC & TEF  ; 
 OBI <=  DBI & TEB  |  EDI & TED  |  WDK & TEF  ; 
 QTB <= QTA ; 
 QTC <= QTB ; 
 QTD <= QTC ; 
 QTE <= QTD ; 
 QTA <=  QTA & qtx  |  QAA & GCH  |  IMB  ; 
 oca <= pca ; 
 oci <= pci ; 
 oda <= pda ; 
 odi <= pdi ; 
 QGC <= IFI ; 
 QGE <= IGC ; 
 QTM <= IMA ; 
 QTN <= QTM ; 
 QGD <=  IGA  |  IGB  ; 
 qtp <=  QTM  |  qtn  ; 
 QTJ <= QTI ; 
 QZD <= QYD ; 
 QYA <= IMC ; 
 QYB <= IMD ; 
 QYC <= IME ; 
 QYD <= IMF ; 
 OEA <= KAA ; 
 KAA <=  KAA & tlc & jma  |  kaa & JMA  |  JNA  ; 
 QZE <=  QZE & qzd  |  QYA  ; 
 LAA <=  IPA & tlb & jcr  |  IQA & TLB  ; 
 PAB <=  PAB & jgb & tpe  |  pab & JGB  |  AAB & TPE  ; 
 PCB <=  PAB & jgb & tpe  |  pab & JGB  |  AAB & TPE  ; 
 PEB <=  PAB & jgb & tpe  |  pab & JGB  |  AAB & TPE  ; 
 PAJ <=  PAJ & jgj & tpb  |  paj & JGJ  |  AAJ & TPB  ; 
 PCJ <=  PAJ & jgj & tpb  |  paj & JGJ  |  AAJ & TPB  ; 
 PEJ <=  PAJ & jgj & tpb  |  paj & JGJ  |  AAJ & TPB  ; 
 qvh <=  jfe  ; 
 qvi <=  jfe  |  jff  ; 
 BAJ <=  BAJ & jdj & tfb  |  baj & JDJ  |  AAJ & TFB  ; 
 BCJ <=  BAJ & jdj & tfb  |  baj & JDJ  |  AAJ & TFB  ; 
 BEJ <=  BAJ & jdj & tfb  |  baj & JDJ  |  AAJ & TFB  ; 
 QWB <= QWA ; 
 QWC <= QWB ; 
 qwi <= jdf ; 
 PBB <=  PBB & jhb & tpc  |  pbb & JHB  |  ABB & TPC  ; 
 PDB <=  PBB & jhb & tpc  |  pbb & JHB  |  ABB & TPC  ; 
 PFB <=  PBB & jhb & tpc  |  pbb & JHB  |  ABB & TPC  ; 
 BBB <=  BBB & jeb & tfc  |  bbb & JEB  |  ABB & TFC  ; 
 BDB <=  BBB & jeb & tfc  |  bbb & JEB  |  ABB & TFC  ; 
 BFB <=  BBB & jeb & tfc  |  bbb & JEB  |  ABB & TFC  ; 
 PBJ <=  PBJ & jhj & tpd  |  pbj & JHB  |  ABJ & TPD  ; 
 PDJ <=  PBJ & jhj & tpd  |  pbj & JHB  |  ABJ & TPD  ; 
 PFJ <=  PBJ & jhj & tpd  |  pbj & JHB  |  ABJ & TPD  ; 
 BBJ <=  BBJ & jej & tfd  |  bbj & JEJ  |  ABJ & TFD  ; 
 BDJ <=  BBJ & jej & tfd  |  bbj & JEJ  |  ABJ & TFD  ; 
 BFJ <=  BBJ & jej & tfd  |  bbj & JEJ  |  ABJ & TFD  ; 
 RHA <= QHA ; 
 RHB <= RHA ; 
 RHC <= RHB ; 
 RHD <= RHC ; 
 RHE <= RHD ; 
 RHF <= RHE ; 
 RHG <= RHF ; 
 RHH <= RHG ; 
 RHI <= RHH ; 
 RHJ <= RHI ; 
 RIA <=  QHA & QIC  ; 
 RIB <=  RHA & QIC  |  RIA & qic  ; 
 RIC <=  RHB & QIC  |  RIB & qic  ; 
 RID <=  RHC & QIC  |  RIC & qic  ; 
 RIE <=  RHD & QIC  |  RID & qic  ; 
 RIF <=  RHE & QIC  |  RIE & qic  ; 
 gab <=  fbh & TGA  |  gab & tga  ; 
 gbj <=  faf & TGC  |  fbc & TGD  |  gbj & tgc  ; 
 qpc <=  qab  |  jfj  ; 
 qpd <=  qab  |  gbk  ; 
 gcb <=  fag & TGE  |  fbb & TGF  |  gcb & tge  ; 
 gcj <=  eab & TGE  |  ZZO & TGF  |  gcj & tge  ; 
 hag <=  gao  |  gad  ; 
 hah <=  gap  |  gad  ; 
 NAB <=  NAB & jsb & tha  |  nab & JSB  |  WCD & THA  ; 
 NBB <=  NAB & jsb & tha  |  nab & JSB  |  WCD & THA  ; 
 QHA <=  RHJ & QRC  |  QLD & qlk  |  GAF & QAA  |  JJH & qrc  ; 
 QKF <=  QKF & hbf  |  QKC & QKD  ; 
 QKG <= JAE ; 
 QKH <= JAF ; 
 QKI <=  qgd & JAI  |  QGD & JAJ  |  qge & JAK  |  QGE & JAL  |  JAD  ; 
 QKK <=  QKA & jic & jid  |  QKK & qkn  ; 
 QKL <= QKK ; 
 QKM <= QKL ; 
 QKN <= QKM ; 
 LBB <=  LBB & jlb & tla  |  lbb & JLB  |  LAB & TLA  ; 
 eab <=  ieb  ; 
 AAB <=  IAB & TAA  |  DAB & TBA  |  IEB & TCA  |  WAB & TDA  |  TMA  ; 
 OAB <=  DAB & TEA  |  EAB & TEC  |  NAB & TEE  ; 
 OAJ <=  DAJ & TEA  |  ECJ & TEC  |  WCL & TEE  ; 
 eaj <=  iej  ; 
 ebj <=  iej  ; 
 ecj <=  iej  ; 
 DAB <= ICB ; 
 DAJ <= ICJ ; 
 EDB <= EAB ; 
 EDJ <= EAJ ; 
 AAJ <=  IAJ & TAB  |  DAJ & TBB  |  IEJ & TCB  |  WAJ & TDA  |  TMB  ; 
 OGD <=  IAJ & TAB  |  DAJ & TBB  |  IEJ & TCB  |  WAJ & TDA  |  TMB  ; 
 DBB <= IDB ; 
 DBJ <= IDJ ; 
 ABB <=  IBB & TAC  |  DBB & TBC  |  EAB & TCC  |  WBB & TDC  |  TMC  ; 
 OGL <=  IBB & TAC  |  DBB & TBC  |  EAB & TCC  |  WBB & TDC  |  TMC  ; 
 orb <= gcj ; 
 OGT <=  IBJ & TAD  |  DBJ & TBD  |  ECJ & TCD  |  WBJ & TDD  |  TMD  ; 
 ABJ <=  IBJ & TAD  |  DBJ & TBD  |  ECJ & TCD  |  WBJ & TDD  |  TMD  ; 
 OBB <=  DBB & TEB  |  EDB & TED  |  WDD & TEF  ; 
 OBJ <=  DBJ & TEB  |  EDJ & TED  |  WDL & TEF  ; 
 QKJ <=  jbe & JAM  |  JBA & JAN  |  qgc & JAO  |  QGC & JAP  |  JBB  ; 
 qza <= qya ; 
 qzb <= qya ; 
 ocb <= pcb ; 
 ocj <= pcj ; 
 odb <= pdb ; 
 odj <= pdj ; 
 OJA <=  RFA & reb  |  WCA & REB  ; 
 RFA <=  RFA & reb  |  WCA & REB  ; 
 QGA <=  ifa  |  ifb  |  ifc  |  ifd  ; 
 OJB <=  RFB & reb  |  WCB & REB  ; 
 RFB <=  RFB & reb  |  WCB & REB  ; 
 CAA <= ILA ; 
 CAB <= ILB ; 
 CAC <= ILC ; 
 OEB <= KAB ; 
 KAB <=  KAB & tlc & jmb  |  kab & JMB  |  JNB  ; 
 RGA <= INA ; 
 RGB <= RGA ; 
 RGC <= RGB ; 
 RGD <= RGC ; 
 LAB <=  IPB & tlb & jcr  |  IQB & TLB  ; 
 PAC <=  PAC & jgc & tpe  |  pac & JGC  |  AAC & TPE  ; 
 PCC <=  PAC & jgc & tpe  |  pac & JGC  |  AAC & TPE  ; 
 PEC <=  PAC & jgc & tpe  |  pac & JGC  |  AAC & TPE  ; 
 PAK <=  PAK & jgk & tpb  |  pak & JGK  |  AAK & TPB  ; 
 PCK <=  PAK & jgk & tpb  |  pak & JGK  |  AAK & TPB  ; 
 PEK <=  PAK & jgk & tpb  |  pak & JGK  |  AAK & TPB  ; 
 QUB <= QPD ; 
 QUC <= QUB ; 
 QUE <= QUD ; 
 BAK <=  BAK & jdk & tfb  |  bak & JDK  |  AAK & TFB  ; 
 BCK <=  BAK & jdk & tfb  |  bak & JDK  |  AAK & TFB  ; 
 BEK <=  BAK & jdk & tfb  |  bak & JDK  |  AAK & TFB  ; 
 QWA <=  JCN  |  JJA  ; 
 QWJ <=  JCN  |  QZF  ; 
 PBC <=  PBC & jhc & tpc  |  pbc & JHC  |  ABC & TPC  ; 
 PDC <=  PBC & jhc & tpc  |  pbc & JHC  |  ABC & TPC  ; 
 PFC <=  PBC & jhc & tpc  |  pbc & JHC  |  ABC & TPC  ; 
 QUA <=  QPA & qpb  ; 
 BBC <=  BBC & jec & tfc  |  bbc & JEC  |  ABC & TFC  ; 
 BDC <=  BBC & jec & tfc  |  bbc & JEC  |  ABC & TFC  ; 
 BFC <=  BBC & jec & tfc  |  bbc & JEC  |  ABC & TFC  ; 
 PBK <=  PBK & jhk & tpd  |  pbk & JHC  |  ABK & TPD  ; 
 PDK <=  PBK & jhk & tpd  |  pbk & JHC  |  ABK & TPD  ; 
 PFK <=  PBK & jhk & tpd  |  pbk & JHC  |  ABK & TPD  ; 
 BBK <=  BBK & jek & tfd  |  bbk & JEK  |  ABK & TFD  ; 
 BDK <=  BBK & jek & tfd  |  bbk & JEK  |  ABK & TFD  ; 
 BFK <=  BBK & jek & tfd  |  bbk & JEK  |  ABK & TFD  ; 
 RMA <= JKB ; 
 RMC <= RMB ; 
 RMD <= RMC ; 
 RNM <= RNL ; 
 RNN <= RNM ; 
 RNO <= RNN ; 
 RNP <= RNO ; 
 RMK <=  RMJ & qhd  |  RMU  ; 
 RMG <= RMF ; 
 RMH <= RMG ; 
 RMI <= RMH ; 
 RMJ <= RMI ; 
 RMN <=  RMQ & QRA  ; 
 RML <= RMK ; 
 RMM <= RML ; 
 RMO <= RMN ; 
 RMP <= RMO ; 
 RMF <=  RME & QRA  |  RNP  ; 
 RMR <=  RMQ & QRA  ; 
 RMQ <= RMP ; 
 RMS <= RMR ; 
 RMT <= RMS ; 
 RMU <= RMT ; 
 gac <=  fac & TGA  |  gac & tga  ; 
 gbc <=  faa & TGC  |  fal & TGD  |  gbc & tgc  ; 
 gbk <=  faf & TGC  |  fal & TGD  |  gbk & tgc  ; 
 QKB <=  JCI & QAC  |  QKB & jaq  ; 
 gcc <=  fag & TGE  |  fbc & TGF  |  gcc & tge  ; 
 gck <=  eac & TGE  |  ZZO & TGF  |  gck & tge  ; 
 qni <=  qac  |  gca  ; 
 qnm <=  qac  |  gcb  ; 
 QKA <=  QKA & qkk  |  GAL & QAC  ; 
 RNL <= RNK ; 
 qnj <= qni ; 
 qnn <= qnm ; 
 NAC <=  NAC & jsc & tha  |  nac & JSC  |  WCE & THA  ; 
 NBC <=  NAC & jsc & tha  |  nac & JSC  |  WCE & THA  ; 
 RNB <= RNA ; 
 RNC <= RNB ; 
 RND <= RNC ; 
 RNA <=  JKB & QHD  |  RME  ; 
 RNK <=  RMJ & QHD  ; 
 RME <=  RKA & jic & jid  |  RMD  ; 
 RMB <=  RMQ & qra  |  RMA  ; 
 LBC <=  LBC & jlc & tla  |  lbc & JLC  |  LAC & TLA  ; 
 eac <=  iec  ; 
 AAC <=  IAC & TAA  |  DAC & TBA  |  IEC & TCA  |  WAC & TDA  |  TMA  ; 
 OHA <=  IAC & TAA  |  DAC & TBA  |  IEC & TCA  |  WAC & TDA  |  TMA  ; 
 OAC <=  DAC & TEA  |  EAC & TEC  |  NAC & TEE  ; 
 OAK <=  DAK & TEA  |  ECK & TEC  |  WCM & TEE  ; 
 eak <=  iek  ; 
 ebk <=  iek  ; 
 eck <=  iek  ; 
 DAC <= ICC ; 
 DAK <= ICK ; 
 EDC <= EAC ; 
 EDK <= EAK ; 
 AAK <=  IAK & TAB  |  DAK & TBB  |  IEK & TCB  |  WAK & TDA  |  TMB  ; 
 OGE <=  IAK & TAB  |  DAK & TBB  |  IEK & TCB  |  WAK & TDA  |  TMB  ; 
 DBC <= IDC ; 
 DBK <= IDK ; 
 QZF <= QZE ; 
 ABC <=  IBC & TAC  |  DBC & TBC  |  EAC & TCC  |  WBC & TDC  |  TMC  ; 
 OGM <=  IBC & TAC  |  DBC & TBC  |  EAC & TCC  |  WBC & TDC  |  TMC  ; 
 orc <= gck ; 
 MAA <=  MAA & tld  |  GAG & TLD  ; 
 ABK <=  IBK & TAD  |  DBK & TBD  |  ECK & TCD  |  WBK & TDD  |  TMD  ; 
 OGU <=  IBK & TAD  |  DBK & TBD  |  ECK & TCD  |  WBK & TDD  |  TMD  ; 
 OBC <=  DBC & TEB  |  EDC & TED  |  WDE & TEF  ; 
 OBK <=  DBK & TEB  |  EDK & TED  |  WDM & TEF  ; 
 QFA <= IMG ; 
 occ <= pcc ; 
 ock <= pck ; 
 odc <= pdc ; 
 odk <= pdk ; 
 QGB <=  ife  |  ifff   |  ifg  |  ifh  ; 
 QKC <=  QKC & jar  |  JBE  ; 
 QKD <=  IKA & JBC  |  IKB & JBD  ; 
 QKE <=  QKB & JBC  |  QKB & JBD  ; 
 OKA <=  IKA & jbc  |  IKA & qkk  |  JBC & QKB  ; 
 OEC <= KAC ; 
 KAC <=  KAC & tlc  |  MAA & QMG  |  JNC  ; 
 OKB <=  IKB & jbd  |  IKB & qkk  |  JBD & QKB  ; 
 LAC <=  IPC & tlb & jcr  |  IQC & TLB  ; 
 PAD <=  PAD & jgd & tpa  |  pad & JGD  |  AAD & TPA  ; 
 PCD <=  PAD & jgd & tpa  |  pad & JGD  |  AAD & TPA  ; 
 PED <=  PAD & jgd & tpa  |  pad & JGD  |  AAD & TPA  ; 
 PAL <=  PAL & jgl & tpb  |  pal & JGL  |  AAL & TPB  ; 
 PCL <=  PAL & jgl & tpb  |  pal & JGL  |  AAL & TPB  ; 
 PEL <=  PAL & jgl & tpb  |  pal & JGL  |  AAL & TPB  ; 
 qvb <=  quf  ; 
 BAL <=  BAL & jdl & tfb  |  bal & JDL  |  AAL & TFB  ; 
 BCL <=  BAL & jdl & tfb  |  bal & JDL  |  AAL & TFB  ; 
 BEL <=  BAL & jdl & tfb  |  bal & JDL  |  AAL & TFB  ; 
 qwd <=  jda  ; 
 PBD <=  PBD & jhd & tpc  |  pbd & JHD  |  ABD & TPC  ; 
 PDD <=  PBD & jhd & tpc  |  pbd & JHD  |  ABD & TPC  ; 
 PFD <=  PBD & jhd & tpc  |  pbd & JHD  |  ABD & TPC  ; 
 QUD <=  QUC  |  QPC  ; 
 BBD <=  BBD & jed & tfc  |  bbd & JED  |  ABD & TFC  ; 
 BDD <=  BBD & jed & tfc  |  bbd & JED  |  ABD & TFC  ; 
 BFD <=  BBD & jed & tfc  |  bbd & JED  |  ABD & TFC  ; 
 PBL <=  PBL & jhl & tpd  |  pbl & JHD  |  ABL & TPD  ; 
 PDL <=  PBL & jhl & tpd  |  pbl & JHD  |  ABL & TPD  ; 
 PFL <=  PBL & jhl & tpd  |  pbl & JHD  |  ABL & TPD  ; 
 BBL <=  BBL & jel & tfd  |  bbl & JEL  |  ABL & TFD  ; 
 BDL <=  BBL & jel & tfd  |  bbl & JEL  |  ABL & TFD  ; 
 BFL <=  BBL & jel & tfd  |  bbl & JEL  |  ABL & TFD  ; 
 RKB <= RKA ; 
 RKC <= RKB ; 
 RKD <= RKC ; 
 RLB <= RLA ; 
 RLC <= RLB ; 
 RLD <= RLC ; 
 QLE <=  JKA & qrb  |  QLC  |  JJE & RLB  ; 
 QLD <=  JKA & qrb & qlo  |  QLC  ; 
 QLK <=  QLK & jjg  |  QLD & JLG  ; 
 QLN <=  RML & rha  |  QLF & QLK  |  QTP  ; 
 QLO <=  RML & rha  |  QLF & QLK  |  QTP  ; 
 QLA <= JBC ; 
 QLB <= QLA ; 
 QLC <= QLB ; 
 QLL <=  QLL & qlm  |  RKD & rmg  ; 
 QLG <=  QLG & jjg  |  RKA  ; 
 QLI <=  QLI & jjg  |  QLJ  ; 
 gad <=  fad & TGA  |  gad & tga  ; 
 gal <=  fad & TGA  |  gal & tga  |  fap & TGB  ; 
 gbd <=  faa & TGC  |  fbc & TGD  |  gbd & tgc  ; 
 gcd <=  fag & TGE  |  fbd & TGF  |  gcd & tge  ; 
 gcl <=  ead & TGE  |  ZZO & TGF  |  gcl & tge  ; 
 qnq <=  qac  |  gcb  ; 
 qnu <=  qac  |  gcd  ; 
 RKA <=  GBO & QAB  ; 
 QLJ <=  GBP & QAB  ; 
 qnr <= qnq ; 
 qnv <= qnu ; 
 NAD <=  NAD & jsd & tha  |  nad & JSD  |  WCF & THA  ; 
 RLA <=  QLD & qlk  |  GAF & QAB  |  JJH & qrc  ; 
 QEA <=  QYB  |  QYC  ; 
 QEB <=  QNQ  |  QNU  ; 
 QLM <=  QLL & jic & jid  ; 
 QRB <= QRA ; 
 QRC <= QRB ; 
 QRD <= QRC ; 
 QRE <= QRD ; 
 QLP <=  QLP & jqa  |  JCL & QAB  |  JXB  |  JQB & JQD  ; 
 QLQ <=  QLP & jqa  |  JCL & QAB  |  JXB  |  JQB & JQD  ; 
 QLF <=  QLF & jjg  |  JCK & QAB  |  RSA  ; 
 LBD <=  LBD & jld & tla  |  lbd & JLD  |  LAD & TLA  ; 
 ead <=  ied  ; 
 AAD <=  IAD & TAA  |  DAD & TBA  |  IED & TCA  |  WAD & TDA  |  TMA  ; 
 OHB <=  IAD & TAA  |  DAD & TBA  |  IED & TCA  |  WAD & TDA  |  TMA  ; 
 OAD <=  DAD & TEA  |  EAD & TEC  |  NAD & TEE  ; 
 OAL <=  DAL & TEA  |  ECL & TEC  |  WCN & TEE  ; 
 eal <=  iel  ; 
 ebl <=  iel  ; 
 ecl <=  iel  ; 
 DAD <= ICD ; 
 DAL <= ICL ; 
 EDD <= EAD ; 
 EDL <= EAL ; 
 AAL <=  IAL & TAB  |  DAL & TBB  |  IEL & TCB  |  WAL & TDA  |  TMB  ; 
 OGF <=  IAL & TAB  |  DAL & TBB  |  IEL & TCB  |  WAL & TDA  |  TMB  ; 
 DBD <= IDD ; 
 DBL <= IDL ; 
 ABD <=  IBD & TAC  |  DBD & TBC  |  EAD & TCC  |  WBD & TDC  |  TMC  ; 
 OGN <=  IBD & TAC  |  DBD & TBC  |  EAD & TCC  |  WBD & TDC  |  TMC  ; 
 ord <= gcl ; 
 MAB <=  MAB & tld  |  GAH & TLD  ; 
 ABL <=  IBL & TAD  |  DBL & TBD  |  ECL & TCD  |  WBL & TDD  |  TMD  ; 
 OGV <=  IBL & TAD  |  DBL & TBD  |  ECL & TCD  |  WBL & TDD  |  TMD  ; 
 OBD <=  DBD & TEB  |  EDD & TED  |  WDF & TEF  ; 
 OBL <=  DBL & TEB  |  EDL & TED  |  WDN & TEF  ; 
 QLR <= QLQ ; 
 QLS <= QLR ; 
 OLF <=  QFB & QLS  |  QFA & qls  ; 
 QFB <=  QFB & QLS  |  QFA & qls  ; 
 ocd <= pcd ; 
 ocl <= pcl ; 
 odd <= pdd ; 
 odl <= pdl ; 
 QCA <= IHA ; 
 QCC <= IHA ; 
 QRF <= QRE ; 
 RIX <= JRB ; 
 QRA <=  RIX  |  JRA  |  QHF  |  IJD  ; 
 OJC <=  RIX  |  JRA  |  IJD  |  JRE  |  QSA  ; 
 OMA <=  QLG & jrc  |  JRB  |  JRD  |  IJD  ; 
 OMB <=  QLG & jrc  |  JRB  |  JRD  |  IJD  ; 
 OTC <= QLQ ; 
 qib <= qia ; 
 qic <= qib ; 
 qid <= qic ; 
 qia <=  ijd & qhf  |  ijd & QRA  ; 
 OED <=  KAD  ; 
 oei <=  qfc  |  QSG  ; 
 KAD <=  KAD & tlc  |  MAB & QMG  |  JND  |  RSC & QSB  ; 
 OJE <=  JCO  ; 
 REB <=  JCO  ; 
 OJD <=  JCO  |  JJB  |  JCA  |  JCB  |  JCF  ; 
 LAD <=  IPD & tlb & jcr  |  IQD & TLB  ; 
 PAE <=  PAE & jge & tpa  |  pae & JGE  |  AAE & TPA  ; 
 PCE <=  PAE & jge & tpa  |  pae & JGE  |  AAE & TPA  ; 
 PEE <=  PAE & jge & tpa  |  pae & JGE  |  AAE & TPA  ; 
 PAM <=  PAM & jgm & tpb  |  pam & JGM  |  AAM & TPB  ; 
 PCM <=  PAM & jgm & tpb  |  pam & JGM  |  AAM & TPB  ; 
 PEM <=  PAM & jgm & tpb  |  pam & JGM  |  AAM & TPB  ; 
 qvc <=  quf  |  jfa  ; 
 BAM <=  BAM & jdm & tfb  |  bam & JDM  |  AAM & TFB  ; 
 BCM <=  BAM & jdm & tfb  |  bam & JDM  |  AAM & TFB  ; 
 BEM <=  BAM & jdm & tfb  |  bam & JDM  |  AAM & TFB  ; 
 qwe <=  jda  |  jdb  ; 
 PBE <=  PBE & jhe & tpc  |  pbe & JHE  |  ABE & TPC  ; 
 PDE <=  PBE & jhe & tpc  |  pbe & JHE  |  ABE & TPC  ; 
 PFE <=  PBE & jhe & tpc  |  pbe & JHE  |  ABE & TPC  ; 
 QUF <=  QPA & JPA  |  QPB  |  QUE  ; 
 BBE <=  BBE & jee & tfc  |  bbe & JEE  |  ABE & TFC  ; 
 BDE <=  BBE & jee & tfc  |  bbe & JEE  |  ABE & TFC  ; 
 BFE <=  BBE & jee & tfc  |  bbe & JEE  |  ABE & TFC  ; 
 PBM <=  PBM & jhm & tpd  |  pbm & JHE  |  ABM & TPD  ; 
 PDM <=  PBM & jhm & tpd  |  pbm & JHE  |  ABM & TPD  ; 
 PFM <=  PBM & jhm & tpd  |  pbm & JHE  |  ABM & TPD  ; 
 BBM <=  BBM & jem & tfd  |  bbm & JEM  |  ABM & TFD  ; 
 BDM <=  BBM & jem & tfd  |  bbm & JEM  |  ABM & TFD  ; 
 BFM <=  BBM & jem & tfd  |  bbm & JEM  |  ABM & TFD  ; 
 gae <=  FAB & TGA  |  GAE & tga  ; 
 gam <=  fad & TGA  |  gam & tga  |  FBE & TGB  ; 
 gbe <=  fae & TGC  |  fbb & TGD  |  gbe & tgc  ; 
 gbm <=  fah & TGC  |  fai & TGD  |  gbm & tgc  ; 
 gcm <=  eae & TGE  |  ZZO  |  gcm & tge  ; 
 qma <=  qac  |  jcl  ; 
 qme <=  qac  |  jcj  ; 
 qmb <= qma ; 
 qmc <= qmb ; 
 qmf <= qme ; 
 qmg <= qmf ; 
 RJK <=  RJK & rjl & jct  |  RJA  ; 
 RJA <=  QAC & GBA  ; 
 RJE <=  RJD & GBA  |  QZD  ; 
 RJB <= RJA ; 
 RJC <= RJB ; 
 RJD <= RJC ; 
 RJL <= RJC ; 
 RAA <=  QAC & GAC & gba  |  RJC  |  QYD  ; 
 RAF <= RAE ; 
 RAG <= RAF ; 
 LBE <=  LBE & jle & tla  |  lbe & JLE  |  LAE & TLA  ; 
 eae <=  iee  ; 
 AAE <=  IAE & TAE  |  DAE & TBE  |  IEE & TCE  |  WAE & TDE  |  TMA  ; 
 OHC <=  IAE & TAE  |  DAE & TBE  |  IEE & TCE  |  WAE & TDE  |  TMA  ; 
 OAE <=  DAE & TEA  |  EAE & TEC  |  WCG & TEE  ; 
 OAM <=  DAM & TEA  |  ECM & TEC  |  WCO & TEE  ; 
 eam <=  iem  ; 
 ecm <=  iem  ; 
 DAE <= ICE ; 
 DAM <= ICM ; 
 EDE <= EAE ; 
 EDM <= EAM ; 
 gbf <=  faf & TGC  |  FBE & TGD  |  gbf & tgc  ; 
 gbn <=  fah & TGC  |  faj & TGD  |  gbn & tgc  ; 
 QXA <=  REC  |  JJI  |  RAA  |  RBA  |  QZE  ; 
 QXB <=  REC  |  JJI  |  RAA  |  RBA  |  QZE  ; 
 DBE <= IDE ; 
 DBM <= IDM ; 
 ABE <=  IBE & TAG  |  DBE & TBG  |  EAE & TCG  |  WBE & TDG  |  TMC  ; 
 OGO <=  IBE & TAG  |  DBE & TBG  |  EAE & TCG  |  WBE & TDG  |  TMC  ; 
 ore <= gcm ; 
 MAC <=  MAC & tld  |  GAI & TLD  ; 
 ABM <=  IBM & TAH  |  DBM & TBH  |  ECM & TCH  |  WBM & TDH  |  TMD  ; 
 OGW <=  IBM & TAH  |  DBM & TBH  |  ECM & TCH  |  WBM & TDH  |  TMD  ; 
 OBE <=  DBE & TEB  |  EDE & TED  |  WDG & TEF  ; 
 OBM <=  DBM & TEB  |  EDM & TED  |  WDO & TEF  ; 
 RJF <= RJE ; 
 RJG <= RJF ; 
 RJH <= RJG ; 
 RJI <= RJH ; 
 OIA <=  JCA  |  JCB  |  JCC & qca  |  JCM  |  QQH  ; 
 REC <=  JCA  |  JCB  |  JCC & qca  |  JCM  |  QQH  ; 
 oce <= pce ; 
 ocm <= pcm ; 
 ode <= pde ; 
 odm <= pdm ; 
 RAB <= RAA ; 
 RAC <= RAB ; 
 RAD <= RAC ; 
 RAE <= RAD ; 
 OIC <=  JCP & QCA  |  JJC & QCA  ; 
 OIB <=  RAC & JJI  |  RBC  ; 
 OID <=  QQH & JJI  ; 
 OEE <= KAE ; 
 OIE <= JCM ; 
 OLC <= QTX ; 
 OTA <= QTX ; 
 KAE <=  KAE & tlc  |  MAC & QMG  |  JNE  ; 
 otd <= qrf ; 
 LAE <=  IPE & tlb & jcr  |  IQE & TLB  |  JCR  ; 
 PAF <=  PAF & jgf & tpa  |  paf & JGF  |  AAF & TPA  ; 
 PCF <=  PAF & jgf & tpa  |  paf & JGF  |  AAF & TPA  ; 
 PEF <=  PAF & jgf & tpa  |  paf & JGF  |  AAF & TPA  ; 
 PAN <=  PAN & jgn & tpb  |  pan & JGN  |  AAN & TPB  ; 
 PCN <=  PAN & jgn & tpb  |  pan & JGN  |  AAN & TPB  ; 
 PEN <=  PAN & jgn & tpb  |  pan & JGN  |  AAN & TPB  ; 
 qvd <=  quf  |  jfa  |  jfb  ; 
 BAN <=  BAN & jdn & tfb  |  ban & JDN  |  AAN & TFB  ; 
 BCN <=  BAN & jdn & tfb  |  ban & JDN  |  AAN & TFB  ; 
 BEN <=  BAN & jdn & tfb  |  ban & JDN  |  AAN & TFB  ; 
 qwf <=  jda  |  jdb  |  jdc  ; 
 PBF <=  PBF & jhf & tpc  |  pbf & JHF  |  ABF & TPC  ; 
 PDF <=  PBF & jhf & tpc  |  pbf & JHF  |  ABF & TPC  ; 
 PFF <=  PBF & jhf & tpc  |  pbf & JHF  |  ABF & TPC  ; 
 BBF <=  BBF & jef & tfc  |  bbf & JEF  |  ABF & TFC  ; 
 BDF <=  BBF & jef & tfc  |  bbf & JEF  |  ABF & TFC  ; 
 BFF <=  BBF & jef & tfc  |  bbf & JEF  |  ABF & TFC  ; 
 PBN <=  PBN & jhn & tpd  |  pbn & JHF  |  ABN & TPD  ; 
 PDN <=  PBN & jhn & tpd  |  pbn & JHF  |  ABN & TPD  ; 
 PFN <=  PBN & jhn & tpd  |  pbn & JHF  |  ABN & TPD  ; 
 BBN <=  BBN & jen & tfd  |  bbn & JEN  |  ABN & TFD  ; 
 BDN <=  BBN & jen & tfd  |  bbn & JEN  |  ABN & TFD  ; 
 BFN <=  BBN & jen & tfd  |  bbn & JEN  |  ABN & TFD  ; 
 QQL <=  JCC & QCC  |  JCG  ; 
 rqa <=  jqb  |  jqd  ; 
 QQM <=  QQL & JJJ  ; 
 QQI <=  RLA & QQD  ; 
 QQN <= QQL ; 
 RQB <= RQA ; 
 rqc <= rqb ; 
 gan <=  fad & TGA  |  gan & tga  |  fbe & TGB  ; 
 gaf <=  fag & TGA  |  gaf & tga  ; 
 AAM <=  IAM & TAF  |  DAM & TBF  |  IEM & TCF  |  WAM & TDF  |  TMB  ; 
 OGG <=  IAM & TAF  |  DAM & TBF  |  IEM & TCF  |  WAM & TDF  |  TMB  ; 
 gcn <=  eaf & TGE  |  ZZO  |  gcn & tge  ; 
 QMK <=  QMJ  |  QMK & jjm  ; 
 qmi <=  qaa  |  jfh & jjm  ; 
 qmj <= qmi ; 
 qqx <= qqd ; 
 QQH <=  QQH & qqc & qtq  |  JJD & qcc  |  JCQ & qcc  ; 
 QQJ <=  QQJ & qqk & qtq  |  JJD & qcc  |  JCQ & qcc  ; 
 QQD <= JJJ ; 
 QQE <= QQD ; 
 QQF <= JJE ; 
 QQG <= QQF ; 
 QQK <=  JJE & RLC & JLG  ; 
 LBF <=  LBF & jlf & tla  |  lbf & JLF  |  LAF & TLA  ; 
 eaf <=  ief  ; 
 AAF <=  IAF & TAE  |  DAF & TBE  |  IEF & TCE  |  WAF & TDE  |  TMA  ; 
 OHD <=  IAF & TAE  |  DAF & TBE  |  IEF & TCE  |  WAF & TDE  |  TMA  ; 
 OAF <=  DAF & TEA  |  EAF & TEC  |  WCH & TEE  ; 
 OAN <=  DAN & TEA  |  ECN & TEC  |  WCP & TEE  ; 
 ean <=  ien  ; 
 ecn <=  ien  ; 
 DAF <= ICF ; 
 DAN <= ICN ; 
 EDF <= EAF ; 
 EDN <= EAN ; 
 AAN <=  IAF & TAF  |  DAN & TBF  |  IEN & TCF  |  WAN & TDF  |  TMB  ; 
 OGH <=  IAF & TAF  |  DAN & TBF  |  IEN & TCF  |  WAN & TDF  |  TMB  ; 
 QXC <=  REC  |  JJJ  |  RAA  |  RBA  |  QZE  ; 
 QXD <=  REC  |  JJJ  |  RAA  |  RBA  |  QZE  ; 
 DBF <= IDF ; 
 DBN <= IDN ; 
 ABF <=  IBF & TAG  |  DBF & TBG  |  EAF & TCG  |  WBF & TDG  |  TMC  ; 
 OGP <=  IBF & TAG  |  DBF & TBG  |  EAF & TCG  |  WBF & TDG  |  TMC  ; 
 orf <= gcn ; 
 ABN <=  IBF & TAH  |  DBN & TBH  |  ECN & TCH  |  WBN & TDH  |  TMD  ; 
 OGX <=  IBF & TAH  |  DBN & TBH  |  ECN & TCH  |  WBN & TDH  |  TMD  ; 
 OBF <=  DBF & TEB  |  EDF & TED  |  WDH & TEF  ; 
 OBN <=  DBN & TEB  |  EDN & TED  |  WDP & TEF  ; 
 RBF <=  RBE & jce  ; 
 RBG <=  RBF & jce  ; 
 RBB <= jce & RBA ; 
 RBC <= jce & RBB ; 
 RBD <= jce & RBC ; 
 RBE <= jce & RBD ; 
 rba <=  ihb  |  JCB  |  JCD  |  JCH  ; 
 ocf <= pcf ; 
 ocn <= pcn ; 
 odf <= pdf ; 
 odn <= pdn ; 
 QQC <=  QQC & jjn & jjp  |  JQC & JQE  ; 
 QHE <= QHD ; 
 QHF <= QHE ; 
 qtq <= qtp ; 
 qtr <= qtp ; 
 QHC <=  IOA  |  IOB  |  IOC  |  IOD  ; 
 OEJ <=  IOA & RMA  |  IOB & RMI  |  IOC & RMI  |  IOD & RMI  |  RMN  ; 
 QHD <=  IOA & RMA  |  IOB & RMI  |  IOC & RMI  |  IOD & RMI  |  RMN  ; 
 QQA <=  QQA & jjl & qtr & qqc  |  ZZO & qtr & qqc  |  RAB & qqc  |  RBE & jce  ; 
 QQB <=  JQF & jjp & ihc  |  JQC & JQE  ; 
 QQW <=  JQF & jjp & ihc  |  JQC & JQE  ; 
 OEM <=  QMK  |  QNN  |  QNR  |  QSE  ; 
 OEF <= KAF ; 
 ote <= qqf ; 
 KAF <=  KAF & tlc  |  QMG  ; 
 OEP <=  QMK  |  QNB  |  QSE  |  JCS  ; 
 LAF <=  IPF & tlb & jcr  |  IQF & TLB  ; 
 PAG <=  PAG & jgg & tpa  |  pag & JGG  |  AAG & TPA  ; 
 PCG <=  PAG & jgg & tpa  |  pag & JGG  |  AAG & TPA  ; 
 PEG <=  PAG & jgg & tpa  |  pag & JGG  |  AAG & TPA  ; 
 BAG <=  BAG & jdg & tfa  |  bag & JDG  |  AAG & TFA  ; 
 BCG <=  BAG & jdg & tfa  |  bag & JDG  |  AAG & TFA  ; 
 BEG <=  BAG & jdg & tfa  |  bag & JDG  |  AAG & TFA  ; 
 PAO <=  PAO & jgo & tpb  |  pao & JGO  |  AAO & TPB  ; 
 PCO <=  PAO & jgo & tpb  |  pao & JGO  |  AAO & TPB  ; 
 PEO <=  PAO & jgo & tpb  |  pao & JGO  |  AAO & TPB  ; 
 qve <=  quf  |  jfa  |  jfb  |  jfc  ; 
 BAO <=  BAO & jdo & tfb  |  bao & JDO  |  AAO & TFB  ; 
 BCO <=  BAO & jdo & tfb  |  bao & JDO  |  AAO & TFB  ; 
 BEO <=  BAO & jdo & tfb  |  bao & JDO  |  AAO & TFB  ; 
 qwg <=  jda  |  jdb  |  jdc  |  jdd  ; 
 PBG <=  PBG & jhg & tpc  |  pbg & JHG  |  ABG & TPC  ; 
 PDG <=  PBG & jhg & tpc  |  pbg & JHG  |  ABG & TPC  ; 
 PFG <=  PBG & jhg & tpc  |  pbg & JHG  |  ABG & TPC  ; 
 BBG <=  BBG & jeg & tfc  |  bbg & JEG  |  ABG & TFC  ; 
 BDG <=  BBG & jeg & tfc  |  bbg & JEG  |  ABG & TFC  ; 
 BFG <=  BBG & jeg & tfc  |  bbg & JEG  |  ABG & TFC  ; 
 PBO <=  PBO & jho & tpd  |  pbo & JHG  |  ABO & TPD  ; 
 PDO <=  PBO & jho & tpd  |  pbo & JHG  |  ABO & TPD  ; 
 PFO <=  PBO & jho & tpd  |  pbo & JHG  |  ABO & TPD  ; 
 BBO <=  BBO & jeo & tfd  |  bbo & JEO  |  ABO & TFD  ; 
 BDO <=  BBO & jeo & tfd  |  bbo & JEO  |  ABO & TFD  ; 
 BFO <=  BBO & jeo & tfd  |  bbo & JEO  |  ABO & TFD  ; 
 gag <=  eag & TGA  |  gag & tga  ; 
 gao <=  fab & TGA  |  gao & tga  |  FBE & TGB  ; 
 gbg <=  fag & TGC  |  fbe & TGD  |  gbg & tgc  ; 
 gbo <=  fah & TGC  |  fak & TGD  |  gbo & tgc  ; 
 qna <=  qac  |  gaf  ; 
 qne <=  qac  |  gaf  |  GAA  ; 
 qnb <= qna ; 
 qnc <= qnb ; 
 qnf <= qne ; 
 qng <= qnf ; 
 eag <=  ieg  ; 
 AAG <=  IAG & TAE  |  DAG & TBE  |  IEG & TCE  |  WAG & TDE  |  TMA  ; 
 OGA <=  IAG & TAE  |  DAG & TBE  |  IEG & TCE  |  WAG & TDE  |  TMA  ; 
 OAG <=  DAG & TEA  |  EAG & TEC  |  WCI & TEE  ; 
 OAO <=  DAO & TEA  |  ECO & TEC  |  WDA & TEE  ; 
 eao <=  ieo  ; 
 eco <=  ieo  ; 
 DAG <= ICG ; 
 DAO <= ICO ; 
 EDG <= EAG ; 
 EDO <= EAO ; 
 AAO <=  IAG & TAF  |  DAO & TBF  |  IEO & TCF  |  WAO & TDF  |  TMB  ; 
 OGI <=  IAG & TAF  |  DAO & TBF  |  IEO & TCF  |  WAO & TDF  |  TMB  ; 
 DBG <= IDG ; 
 DBO <= IDO ; 
 ABG <=  IBG & TAG  |  DBG & TBG  |  EAG & TCG  |  WBG & TDG  |  TMC  ; 
 OGQ <=  IBG & TAG  |  DBG & TBG  |  EAG & TCG  |  WBG & TDG  |  TMC  ; 
 qsi <= iqi ; 
 ABO <=  IBG & TAH  |  DBO & TBH  |  ECO & TCH  |  WBO & TDH  |  TMD  ; 
 OBG <=  DBG & TEB  |  EDG & TED  |  WDI & TEF  ; 
 OBO <=  DBO & TEB  |  EDO & TED  ; 
 old <=  qaa  |  gch  ; 
 ocg <= pcg ; 
 oco <= pco ; 
 odg <= pdg ; 
 odo <= pdo ; 
 OES <=  JJK & QMK  |  JKE  |  JJF  ; 
 OFC <= QRD ; 
 OLB <= QKK ; 
 OQB <= JXA ; 
 otf <= qsd ; 
 OET <=  JKC  |  QMJ  |  QNA  |  RQB  ; 
 OEH <= QRF ; 
 OEQ <= QQF ; 
 oer <= rsa ; 
 OFA <=  RLB & QNB  ; 
 OLA <=  qkd & QKE  ; 
 ofb <=  rlb  |  qsh  |  QSB  ; 
 oqa <=  rla  |  qsh  |  QSB  ; 
 PAH <=  PAH & jgh & tpa  |  pah & JGH  |  AAH & TPA  ; 
 PCH <=  PAH & jgh & tpa  |  pah & JGH  |  AAH & TPA  ; 
 PEH <=  PAH & jgh & tpa  |  pah & JGH  |  AAH & TPA  ; 
 BAH <=  BAH & jdh & tfa  |  bah & JDH  |  AAH & TFA  ; 
 BCH <=  BAH & jdh & tfa  |  bah & JDH  |  AAH & TFA  ; 
 BEH <=  BAH & jdh & tfa  |  bah & JDH  |  AAH & TFA  ; 
 PAP <=  PAP & jgp & tpb  |  pap & JGP  |  AAP & TPB  ; 
 PCP <=  PAP & jgp & tpb  |  pap & JGP  |  AAP & TPB  ; 
 PEP <=  PAP & jgp & tpb  |  pap & JGP  |  AAP & TPB  ; 
 qvf <=  quf  |  jfa  |  jfb  |  jfc  |  jfd  ; 
 qvg <=  quf  |  jfa  |  jfb  |  jfc  |  jfd  ; 
 BAP <=  BAP & jdp & tfb  |  bap & JDP  |  AAP & TFB  ; 
 BCP <=  BAP & jdp & tfb  |  bap & JDP  |  AAP & TFB  ; 
 BEP <=  BAP & jdp & tfb  |  bap & JDP  |  AAP & TFB  ; 
 qwh <=  jda  |  jdb  |  jdc  |  jdd  |  jde  ; 
 PBH <=  PBH & jhh & tpc  |  pbh & JHH  |  ABH & TPC  ; 
 PDH <=  PBH & jhh & tpc  |  pbh & JHH  |  ABH & TPC  ; 
 PFH <=  PBH & jhh & tpc  |  pbh & JHH  |  ABH & TPC  ; 
 BBH <=  BBH & jeh & tfc  |  bbh & JEH  |  ABH & TFC  ; 
 BDH <=  BBH & jeh & tfc  |  bbh & JEH  |  ABH & TFC  ; 
 BFH <=  BBH & jeh & tfc  |  bbh & JEH  |  ABH & TFC  ; 
 PBP <=  PBP & jhp & tpd  |  pbp & JHH  |  ABP & TPD  ; 
 PDP <=  PBP & jhp & tpd  |  pbp & JHH  |  ABP & TPD  ; 
 PFP <=  PBP & jhp & tpd  |  pbp & JHH  |  ABP & TPD  ; 
 BBP <=  BBP & jep & tfd  |  bbp & JEP  |  ABP & TFD  ; 
 BDP <=  BBP & jep & tfd  |  bbp & JEP  |  ABP & TFD  ; 
 BFP <=  BBP & jep & tfd  |  bbp & JEP  |  ABP & TFD  ; 
 gah <=  eah & TGA  |  gah & tga  ; 
 gap <=  fab & TGA  |  gap & tga  |  fbe & TGB  ; 
 gbh <=  fae & TGC  |  fba & TGD  |  gbh & tgc  ; 
 gbp <=  fah & TGC  |  fal & TGD  |  gbp & tgc  ; 
 gch <=  faa & TGE  |  fba & TGF  |  gch & tge  ; 
 QSC <=  QSC & jxb  |  RRF  ; 
 QSD <=  QSD & jjm  |  RRH  ; 
 RSA <= RRH ; 
 RSB <= RSA ; 
 RSC <= RSB ; 
 QSE <= QSD ; 
 QSF <= QSE ; 
 QSG <= QSF ; 
 eah <=  ieh  ; 
 AAH <=  IAH & TAE  |  DAH & TBE  |  IEH & TCE  |  WAH & TDE  |  TMA  ; 
 OGB <=  IAH & TAE  |  DAH & TBE  |  IEH & TCE  |  WAH & TDE  |  TMA  ; 
 OAH <=  DAH & TEA  |  EAH & TEC  |  WCJ & TEE  ; 
 OAP <=  DAP & TEA  |  ECP & TEC  |  WDB & TEE  ; 
 eap <=  iep  ; 
 ebp <=  iep  ; 
 ecp <=  iep  ; 
 DAH <= ICH ; 
 DAP <= ICP ; 
 EDH <= EAH ; 
 EDP <= EAP ; 
 AAP <=  IAH & TAF  |  DAP & TBF  |  IEP & TCF  |  WAP & TDF  |  TMB  ; 
 OGJ <=  IAH & TAF  |  DAP & TBF  |  IEP & TCF  |  WAP & TDF  |  TMB  ; 
 DBH <= IDH ; 
 DBP <= IDP ; 
 QBA <= IJC ; 
 ABH <=  IBH & TAG  |  DBH & TBG  |  EAH & TCG  |  WBH & TDG  |  TMC  ; 
 OGR <=  IBH & TAG  |  DBH & TBG  |  EAH & TCG  |  WBH & TDG  |  TMC  ; 
 ABP <=  IBH & TAH  |  DBP & TBH  |  ECP & TCH  |  WBP & TDH  |  TMD  ; 
 OBH <=  DBH & TEB  |  EDH & TED  |  WDJ & TEF  ; 
 OBP <=  DBP & TEB  |  EDP & TED  ; 
 QSB <=  QSB & jxa & qtp  |  IQH  ; 
 QSA <=  QSA & jxa & qtp  |  IQG  ; 
 QAA <= IJB & IJA ; 
 QAB <= IJB & IJA ; 
 QAC <= IJB & IJA ; 
 QAD <= IJB & IJA ; 
 och <= pch ; 
 ocp <= pcp ; 
 odh <= pdh ; 
 odp <= pdp ; 
 RRE <= RRD ; 
 RRF <= RRE ; 
 RRG <= JXB ; 
 RRH <= RRG ; 
 RRA <= IQG ; 
 RRB <= RRA ; 
 RRC <= RRB ; 
 RRD <= RRC ; 
 OEG <=  RLD & qqg  |  RLD & QQJ  ; 
 qfc <=  RLD & qqg  |  RLD & QQJ  ; 
 QSH <= QSD & QSF ; 
 OEL <=  RKA  |  QLJ  |  JKD  ; 
 OEV <=  QNQ  |  QNU  |  QQD  ; 
 OEN <= JKC ; 
 OEO <= JKC ; 
 OEX <= QYB ; 
 OEY <= QYC ; 
 OEK <=  JJK & QSG  ; 
 OEU <=  QMI  |  QNI  ; 
 OEW <=  QMK  |  QMJ  ; 
end
endmodule;
