module kc( IZZ,
 IAA, 
 IAB, 
 IAC, 
 IAD, 
 IAE, 
 IAF, 
 IAG, 
 IAH, 
 IAI, 
 IAJ, 
 IAK, 
 IAL, 
 IAM, 
 IAN, 
 IAO, 
 IAP, 
 IBA, 
 IBB, 
 IBC, 
 IBD, 
 IBE, 
 IBF, 
 IBG, 
 IBH, 
 IBI, 
 IBJ, 
 IBK, 
 IBL, 
 IBM, 
 IBN, 
 IBO, 
 IBP, 
 ICA, 
 ICB, 
 ICC, 
 ICD, 
 ICE, 
 ICF, 
 ICG, 
 ICH, 
 ICI, 
 ICJ, 
 ICK, 
 ICL, 
 ICM, 
 ICN, 
 ICO, 
 ICP, 
 IDA, 
 IDB, 
 IDC, 
 IDD, 
 IDE, 
 IDF, 
 IDG, 
 IDH, 
 IDI, 
 IDJ, 
 IDK, 
 IDL, 
 IDM, 
 IDN, 
 IDO, 
 IDP, 
 IFA, 
 IFB, 
 IFC, 
 IFD, 
 IFE, 
 IFFF , 
 IFG, 
 IFH, 
 IFI, 
 IFJ, 
 IFK, 
 IFL, 
 OAA, 
 OAB, 
 OAC, 
 OAD, 
 OAE, 
 OAF, 
 OAG, 
 OAH, 
 OAI, 
 OAJ, 
 OAK, 
 OAL, 
 OAM, 
 OAN, 
 OAO, 
 OAP, 
 OBA, 
 OBB, 
 OBC, 
 OBD, 
 OBE, 
 OBF, 
 OBG, 
 OBH, 
 OBI, 
 OBJ, 
 OBK, 
 OBL, 
 OBM, 
 OBN, 
 OBO, 
 OBP, 
 OCA, 
 OCB, 
 OCC, 
 OCD, 
 OCE, 
 OCF, 
 OCG, 
 OCH, 
 OCI, 
 OCJ, 
 OCK, 
 OCL, 
 OCM, 
 OCN, 
 OCO, 
 OCP, 
 ODA, 
 ODB, 
 ODC, 
 ODD, 
 ODE, 
 ODF, 
 ODG, 
 ODH, 
 ODI, 
 ODJ, 
 ODK, 
 ODL, 
 ODM, 
 ODN, 
 ODO, 
 ODP, 
 OEA, 
 OEB, 
OEC ); 
    
 input IZZ; 
 input IAA; 
 input IAB; 
 input IAC; 
 input IAD; 
 input IAE; 
 input IAF; 
 input IAG; 
 input IAH; 
 input IAI; 
 input IAJ; 
 input IAK; 
 input IAL; 
 input IAM; 
 input IAN; 
 input IAO; 
 input IAP; 
 input IBA; 
 input IBB; 
 input IBC; 
 input IBD; 
 input IBE; 
 input IBF; 
 input IBG; 
 input IBH; 
 input IBI; 
 input IBJ; 
 input IBK; 
 input IBL; 
 input IBM; 
 input IBN; 
 input IBO; 
 input IBP; 
 input ICA; 
 input ICB; 
 input ICC; 
 input ICD; 
 input ICE; 
 input ICF; 
 input ICG; 
 input ICH; 
 input ICI; 
 input ICJ; 
 input ICK; 
 input ICL; 
 input ICM; 
 input ICN; 
 input ICO; 
 input ICP; 
 input IDA; 
 input IDB; 
 input IDC; 
 input IDD; 
 input IDE; 
 input IDF; 
 input IDG; 
 input IDH; 
 input IDI; 
 input IDJ; 
 input IDK; 
 input IDL; 
 input IDM; 
 input IDN; 
 input IDO; 
 input IDP; 
 input IFA; 
 input IFB; 
 input IFC; 
 input IFD; 
 input IFE; 
 input IFFF ; 
 input IFG; 
 input IFH; 
 input IFI; 
 input IFJ; 
 input IFK; 
 input IFL; 
 output OAA; 
 output OAB; 
 output OAC; 
 output OAD; 
 output OAE; 
 output OAF; 
 output OAG; 
 output OAH; 
 output OAI; 
 output OAJ; 
 output OAK; 
 output OAL; 
 output OAM; 
 output OAN; 
 output OAO; 
 output OAP; 
 output OBA; 
 output OBB; 
 output OBC; 
 output OBD; 
 output OBE; 
 output OBF; 
 output OBG; 
 output OBH; 
 output OBI; 
 output OBJ; 
 output OBK; 
 output OBL; 
 output OBM; 
 output OBN; 
 output OBO; 
 output OBP; 
 output OCA; 
 output OCB; 
 output OCC; 
 output OCD; 
 output OCE; 
 output OCF; 
 output OCG; 
 output OCH; 
 output OCI; 
 output OCJ; 
 output OCK; 
 output OCL; 
 output OCM; 
 output OCN; 
 output OCO; 
 output OCP; 
 output ODA; 
 output ODB; 
 output ODC; 
 output ODD; 
 output ODE; 
 output ODF; 
 output ODG; 
 output ODH; 
 output ODI; 
 output ODJ; 
 output ODK; 
 output ODL; 
 output ODM; 
 output ODN; 
 output ODO; 
 output ODP; 
 output OEA; 
 output OEB; 
 output OEC; 
  
  
reg  AAA ;
reg  AAB ;
reg  AAC ;
reg  AAD ;
reg  AAE ;
reg  AAF ;
reg  AAG ;
reg  AAH ;
reg  AAI ;
reg  AAJ ;
reg  AAK ;
reg  AAL ;
reg  AAM ;
reg  AAN ;
reg  AAO ;
reg  AAP ;
reg  ABA ;
reg  ABB ;
reg  ABC ;
reg  ABD ;
reg  ABE ;
reg  ABF ;
reg  ABG ;
reg  ABH ;
reg  ABI ;
reg  ABJ ;
reg  ABK ;
reg  ABL ;
reg  ABM ;
reg  ABN ;
reg  ABO ;
reg  ABP ;
reg  BAA ;
reg  BAB ;
reg  BAC ;
reg  BAD ;
reg  BAE ;
reg  BAF ;
reg  BAG ;
reg  BAH ;
reg  BAI ;
reg  BAJ ;
reg  BAK ;
reg  BAL ;
reg  BAM ;
reg  BAN ;
reg  BAO ;
reg  BAP ;
reg  BBA ;
reg  BBB ;
reg  BBC ;
reg  BBD ;
reg  BBE ;
reg  BBF ;
reg  BBG ;
reg  BBH ;
reg  BBI ;
reg  BBJ ;
reg  BBK ;
reg  BBL ;
reg  BBM ;
reg  BBN ;
reg  BBO ;
reg  BBP ;
reg  BCA ;
reg  BCB ;
reg  BCC ;
reg  BCD ;
reg  BCE ;
reg  BCF ;
reg  BCG ;
reg  BCH ;
reg  BCI ;
reg  BCJ ;
reg  BCK ;
reg  BCL ;
reg  BCM ;
reg  BCN ;
reg  BCO ;
reg  BCP ;
reg  BDA ;
reg  BDB ;
reg  BDC ;
reg  BDD ;
reg  BDE ;
reg  BDF ;
reg  BDG ;
reg  BDH ;
reg  BDI ;
reg  BDJ ;
reg  BDK ;
reg  BDL ;
reg  BDM ;
reg  BDN ;
reg  BDO ;
reg  BDP ;
reg  EAA ;
reg  EAB ;
reg  EAC ;
reg  EAD ;
reg  EBA ;
reg  EBB ;
reg  EBC ;
reg  EBD ;
reg  ECA ;
reg  ECB ;
reg  ECC ;
reg  ECD ;
reg  EDA ;
reg  EDB ;
reg  EDC ;
reg  EDD ;
reg  EEA ;
reg  EEB ;
reg  EEC ;
reg  EED ;
reg  EFA ;
reg  EFB ;
reg  EFC ;
reg  EFD ;
reg  EGA ;
reg  EGB ;
reg  EGC ;
reg  EGD ;
reg  EHA ;
reg  EHB ;
reg  EHC ;
reg  EHD ;
reg  eia ;
reg  eib ;
reg  eic ;
reg  eid ;
reg  eja ;
reg  ejb ;
reg  ejc ;
reg  ejd ;
reg  eka ;
reg  ekb ;
reg  ekc ;
reg  ekd ;
reg  ela ;
reg  elb ;
reg  elc ;
reg  eld ;
reg  ema ;
reg  emb ;
reg  emc ;
reg  emd ;
reg  ena ;
reg  enb ;
reg  enc ;
reg  endd ;
reg  eoa ;
reg  eob ;
reg  eoc ;
reg  eod ;
reg  epa ;
reg  epb ;
reg  epc ;
reg  epd ;
reg  HAA ;
reg  HAB ;
reg  HAC ;
reg  HAD ;
reg  HAE ;
reg  haf ;
reg  HAG ;
reg  hah ;
reg  hai ;
reg  HAJ ;
reg  HAK ;
reg  HBA ;
reg  HBB ;
reg  HBC ;
reg  HBD ;
reg  HCA ;
reg  HCB ;
reg  HCC ;
reg  HCD ;
reg  HDA ;
reg  HDB ;
reg  HDC ;
reg  HDD ;
reg  HEA ;
reg  HEB ;
reg  HEC ;
reg  HED ;
reg  HFA ;
reg  HFB ;
reg  HFC ;
reg  HFD ;
reg  HGA ;
reg  HGB ;
reg  HGC ;
reg  HGD ;
reg  HHA ;
reg  HHB ;
reg  HHC ;
reg  HHD ;
reg  HIA ;
reg  HIB ;
reg  HIC ;
reg  HID ;
reg  HJA ;
reg  HJB ;
reg  HJC ;
reg  HJD ;
reg  HKA ;
reg  HKB ;
reg  HKC ;
reg  HKD ;
reg  HLA ;
reg  HLB ;
reg  HLC ;
reg  HLD ;
reg  HMA ;
reg  HMB ;
reg  HMC ;
reg  HMD ;
reg  HNA ;
reg  HNB ;
reg  HNC ;
reg  HND ;
reg  HOA ;
reg  HOB ;
reg  HOC ;
reg  HOD ;
reg  HPA ;
reg  HPB ;
reg  HPC ;
reg  HPD ;
reg  HQA ;
reg  HQB ;
reg  HQC ;
reg  HQD ;
reg  KAA ;
reg  KAB ;
reg  KAC ;
reg  KAD ;
reg  KAE ;
reg  KAF ;
reg  KAG ;
reg  KAH ;
reg  KAI ;
reg  KAJ ;
reg  KAK ;
reg  KAL ;
reg  KAM ;
reg  KAN ;
reg  KAO ;
reg  KAP ;
reg  KBA ;
reg  KBB ;
reg  KBC ;
reg  KBD ;
reg  KBE ;
reg  KBF ;
reg  KBG ;
reg  KBH ;
reg  KBI ;
reg  KBJ ;
reg  KBK ;
reg  KBL ;
reg  KBM ;
reg  KBN ;
reg  KBO ;
reg  KBP ;
reg  KKA ;
reg  LAA ;
reg  LAB ;
reg  LAC ;
reg  LAE ;
reg  LAF ;
reg  LAG ;
reg  LAH ;
reg  LAI ;
reg  LAJ ;
reg  LAK ;
reg  LAL ;
reg  LAM ;
reg  LAN ;
reg  LAO ;
reg  LAP ;
reg  LBA ;
reg  LBB ;
reg  LBC ;
reg  LBD ;
reg  LBE ;
reg  LBF ;
reg  LBG ;
reg  LBH ;
reg  LBI ;
reg  LBJ ;
reg  LBK ;
reg  LBL ;
reg  LBM ;
reg  LBN ;
reg  LBO ;
reg  LBP ;
reg  MAA ;
reg  MAB ;
reg  MAC ;
reg  MAD ;
reg  MAE ;
reg  MAF ;
reg  MAG ;
reg  MAH ;
reg  MAI ;
reg  MAJ ;
reg  MAK ;
reg  MAL ;
reg  MAM ;
reg  MAN ;
reg  MAO ;
reg  MAP ;
reg  MBA ;
reg  MBB ;
reg  MBC ;
reg  MBD ;
reg  MBE ;
reg  MBF ;
reg  MBG ;
reg  MBH ;
reg  MBI ;
reg  MBJ ;
reg  MBK ;
reg  MBL ;
reg  MBM ;
reg  MBN ;
reg  MBO ;
reg  MBP ;
reg  OAA ;
reg  OAB ;
reg  OAC ;
reg  OAD ;
reg  OAE ;
reg  OAF ;
reg  OAG ;
reg  OAH ;
reg  OAI ;
reg  OAJ ;
reg  OAK ;
reg  OAL ;
reg  OAM ;
reg  OAN ;
reg  OAO ;
reg  OAP ;
reg  OBA ;
reg  OBB ;
reg  OBC ;
reg  OBD ;
reg  OBE ;
reg  OBF ;
reg  OBG ;
reg  OBH ;
reg  OBI ;
reg  OBJ ;
reg  OBK ;
reg  OBL ;
reg  OBM ;
reg  OBN ;
reg  OBO ;
reg  OBP ;
reg  OCA ;
reg  OCB ;
reg  OCC ;
reg  OCD ;
reg  OCE ;
reg  OCF ;
reg  OCG ;
reg  OCH ;
reg  OCI ;
reg  OCJ ;
reg  OCK ;
reg  OCL ;
reg  OCM ;
reg  OCN ;
reg  OCO ;
reg  OCP ;
reg  ODA ;
reg  ODB ;
reg  ODC ;
reg  ODD ;
reg  ODE ;
reg  ODF ;
reg  ODG ;
reg  ODH ;
reg  ODI ;
reg  ODJ ;
reg  ODK ;
reg  ODL ;
reg  ODM ;
reg  ODN ;
reg  ODO ;
reg  ODP ;
reg  oea ;
reg  oeb ;
reg  OEC ;
reg  QAA ;
reg  QAB ;
reg  QAC ;
reg  QAD ;
reg  QAE ;
reg  QAF ;
reg  QAG ;
reg  QAH ;
reg  QAI ;
reg  QAJ ;
reg  QAK ;
reg  QAL ;
reg  QAP ;
reg  QAQ ;
reg  QBA ;
reg  QBB ;
reg  QBC ;
reg  QBD ;
reg  QBH ;
reg  QBI ;
reg  QBJ ;
reg  QBK ;
reg  QBL ;
reg  QDA ;
reg  QDB ;
reg  QDC ;
reg  qdd ;
reg  QEA ;
reg  QEB ;
reg  QEC ;
reg  QFA ;
reg  QFB ;
reg  QFC ;
reg  QFD ;
reg  QGE ;
reg  taa ;
reg  tab ;
reg  TBA ;
reg  TBB ;
reg  TCA ;
reg  TCB ;
reg  TDA ;
reg  TDB ;
reg  tea ;
reg  teb ;
reg  TFA ;
reg  TFB ;
reg  TGA ;
reg  TGB ;
reg  TIA ;
reg  TIB ;
reg  TJA ;
reg  TJB ;
reg  TLA ;
reg  TLB ;
reg  TLC ;
reg  TMA ;
reg  TMB ;
reg  TMC ;
reg  TNA ;
reg  TNB ;
reg  TOA ;
reg  TOB ;
reg  TPA ;
reg  TPB ;
reg  TPC ;
reg  TPD ;
reg  TPE ;
reg  TPF ;
reg  TPG ;
reg  TPH ;
reg  TQA ;
reg  TQB ;
reg  TQC ;
reg  TQD ;
reg  TQE ;
reg  TQF ;
reg  TQG ;
reg  TQH ;
reg  TRA ;
reg  TRB ;
reg  TSA ;
reg  TSB ;
reg  TSC ;
reg  TSD ;
reg  TTA ;
reg  TTB ;
wire  aaa ;
wire  aab ;
wire  aac ;
wire  aad ;
wire  aae ;
wire  aaf ;
wire  aag ;
wire  aah ;
wire  aai ;
wire  aaj ;
wire  aak ;
wire  aal ;
wire  aam ;
wire  aan ;
wire  aao ;
wire  aap ;
wire  aba ;
wire  abb ;
wire  abc ;
wire  abd ;
wire  abe ;
wire  abf ;
wire  abg ;
wire  abh ;
wire  abi ;
wire  abj ;
wire  abk ;
wire  abl ;
wire  abm ;
wire  abn ;
wire  abo ;
wire  abp ;
wire  aca ;
wire  ACA ;
wire  acb ;
wire  ACB ;
wire  acc ;
wire  ACC ;
wire  acd ;
wire  ACD ;
wire  ace ;
wire  ACE ;
wire  acf ;
wire  ACF ;
wire  acg ;
wire  ACG ;
wire  ach ;
wire  ACH ;
wire  aci ;
wire  ACI ;
wire  acj ;
wire  ACJ ;
wire  ack ;
wire  ACK ;
wire  acl ;
wire  ACL ;
wire  acm ;
wire  ACM ;
wire  acn ;
wire  ACN ;
wire  aco ;
wire  ACO ;
wire  acp ;
wire  ACP ;
wire  ada ;
wire  ADA ;
wire  adb ;
wire  ADB ;
wire  adc ;
wire  ADC ;
wire  add ;
wire  ADD ;
wire  ade ;
wire  ADE ;
wire  adf ;
wire  ADF ;
wire  adg ;
wire  ADG ;
wire  adh ;
wire  ADH ;
wire  adi ;
wire  ADI ;
wire  adj ;
wire  ADJ ;
wire  adk ;
wire  ADK ;
wire  adl ;
wire  ADL ;
wire  adm ;
wire  ADM ;
wire  adn ;
wire  ADN ;
wire  ado ;
wire  ADO ;
wire  adp ;
wire  ADP ;
wire  baa ;
wire  bab ;
wire  bac ;
wire  bad ;
wire  bae ;
wire  baf ;
wire  bag ;
wire  bah ;
wire  bai ;
wire  baj ;
wire  bak ;
wire  bal ;
wire  bam ;
wire  ban ;
wire  bao ;
wire  bap ;
wire  bba ;
wire  bbb ;
wire  bbc ;
wire  bbd ;
wire  bbe ;
wire  bbf ;
wire  bbg ;
wire  bbh ;
wire  bbi ;
wire  bbj ;
wire  bbk ;
wire  bbl ;
wire  bbm ;
wire  bbn ;
wire  bbo ;
wire  bbp ;
wire  bca ;
wire  bcb ;
wire  bcc ;
wire  bcd ;
wire  bce ;
wire  bcf ;
wire  bcg ;
wire  bch ;
wire  bci ;
wire  bcj ;
wire  bck ;
wire  bcl ;
wire  bcm ;
wire  bcn ;
wire  bco ;
wire  bcp ;
wire  bda ;
wire  bdb ;
wire  bdc ;
wire  bdd ;
wire  bde ;
wire  bdf ;
wire  bdg ;
wire  bdh ;
wire  bdi ;
wire  bdj ;
wire  bdk ;
wire  bdl ;
wire  bdm ;
wire  bdn ;
wire  bdo ;
wire  bdp ;
wire  daa ;
wire  DAA ;
wire  dab ;
wire  DAB ;
wire  dac ;
wire  DAC ;
wire  dad ;
wire  DAD ;
wire  dae ;
wire  DAE ;
wire  daf ;
wire  DAF ;
wire  dag ;
wire  DAG ;
wire  dah ;
wire  DAH ;
wire  dai ;
wire  DAI ;
wire  daj ;
wire  DAJ ;
wire  dak ;
wire  DAK ;
wire  dal ;
wire  DAL ;
wire  dam ;
wire  DAM ;
wire  dan ;
wire  DAN ;
wire  dao ;
wire  DAO ;
wire  dap ;
wire  DAP ;
wire  dba ;
wire  DBA ;
wire  dbb ;
wire  DBB ;
wire  dbc ;
wire  DBC ;
wire  dbd ;
wire  DBD ;
wire  dbe ;
wire  DBE ;
wire  dbf ;
wire  DBF ;
wire  dbg ;
wire  DBG ;
wire  dbh ;
wire  DBH ;
wire  dbi ;
wire  DBI ;
wire  dbj ;
wire  DBJ ;
wire  dbk ;
wire  DBK ;
wire  dbl ;
wire  DBL ;
wire  dbm ;
wire  DBM ;
wire  dbn ;
wire  DBN ;
wire  dbo ;
wire  DBO ;
wire  dbp ;
wire  DBP ;
wire  eaa ;
wire  eab ;
wire  eac ;
wire  ead ;
wire  eba ;
wire  ebb ;
wire  ebc ;
wire  ebd ;
wire  eca ;
wire  ecb ;
wire  ecc ;
wire  ecd ;
wire  eda ;
wire  edb ;
wire  edc ;
wire  edd ;
wire  eea ;
wire  eeb ;
wire  eec ;
wire  eed ;
wire  efa ;
wire  efb ;
wire  efc ;
wire  efd ;
wire  ega ;
wire  egb ;
wire  egc ;
wire  egd ;
wire  eha ;
wire  ehb ;
wire  ehc ;
wire  ehd ;
wire  EIA ;
wire  EIB ;
wire  EIC ;
wire  EID ;
wire  EJA ;
wire  EJB ;
wire  EJC ;
wire  EJD ;
wire  EKA ;
wire  EKB ;
wire  EKC ;
wire  EKD ;
wire  ELA ;
wire  ELB ;
wire  ELC ;
wire  ELD ;
wire  EMA ;
wire  EMB ;
wire  EMC ;
wire  EMD ;
wire  ENA ;
wire  ENB ;
wire  ENC ;
wire  ENDD  ;
wire  EOA ;
wire  EOB ;
wire  EOC ;
wire  EOD ;
wire  EPA ;
wire  EPB ;
wire  EPC ;
wire  EPD ;
wire  gab ;
wire  GAB ;
wire  gac ;
wire  GAC ;
wire  gad ;
wire  GAD ;
wire  gae ;
wire  GAE ;
wire  gaf ;
wire  GAF ;
wire  gag ;
wire  GAG ;
wire  gah ;
wire  GAH ;
wire  gbb ;
wire  GBB ;
wire  gbc ;
wire  GBC ;
wire  gbd ;
wire  GBD ;
wire  gbe ;
wire  GBE ;
wire  gbf ;
wire  GBF ;
wire  gbg ;
wire  GBG ;
wire  gbh ;
wire  GBH ;
wire  gcb ;
wire  GCB ;
wire  gcc ;
wire  GCC ;
wire  gcd ;
wire  GCD ;
wire  gce ;
wire  GCE ;
wire  gcf ;
wire  GCF ;
wire  gcg ;
wire  GCG ;
wire  gch ;
wire  GCH ;
wire  gdb ;
wire  GDB ;
wire  gdc ;
wire  GDC ;
wire  gdd ;
wire  GDD ;
wire  gde ;
wire  GDE ;
wire  gdf ;
wire  GDF ;
wire  gdg ;
wire  GDG ;
wire  gdh ;
wire  GDH ;
wire  geb ;
wire  GEB ;
wire  gec ;
wire  GEC ;
wire  ged ;
wire  GED ;
wire  gee ;
wire  GEE ;
wire  gef ;
wire  GEF ;
wire  geg ;
wire  GEG ;
wire  geh ;
wire  GEH ;
wire  gfb ;
wire  GFB ;
wire  gfc ;
wire  GFC ;
wire  gfd ;
wire  GFD ;
wire  gfe ;
wire  GFE ;
wire  gff ;
wire  GFF ;
wire  gfg ;
wire  GFG ;
wire  gfh ;
wire  GFH ;
wire  ggb ;
wire  GGB ;
wire  ggc ;
wire  GGC ;
wire  ggd ;
wire  GGD ;
wire  gge ;
wire  GGE ;
wire  ggf ;
wire  GGF ;
wire  ggg ;
wire  GGG ;
wire  ggh ;
wire  GGH ;
wire  ghb ;
wire  GHB ;
wire  ghc ;
wire  GHC ;
wire  ghd ;
wire  GHD ;
wire  ghf ;
wire  GHF ;
wire  ghg ;
wire  GHG ;
wire  ghh ;
wire  GHH ;
wire  gia ;
wire  GIA ;
wire  gja ;
wire  GJA ;
wire  gka ;
wire  GKA ;
wire  gla ;
wire  GLA ;
wire  gma ;
wire  GMA ;
wire  gna ;
wire  GNA ;
wire  gpa ;
wire  GPA ;
wire  gqa ;
wire  GQA ;
wire  haa ;
wire  hab ;
wire  hac ;
wire  had ;
wire  hae ;
wire  HAF ;
wire  hag ;
wire  HAH ;
wire  HAI ;
wire  haj ;
wire  hak ;
wire  hba ;
wire  hbb ;
wire  hbc ;
wire  hbd ;
wire  hca ;
wire  hcb ;
wire  hcc ;
wire  hcd ;
wire  hda ;
wire  hdb ;
wire  hdc ;
wire  hdd ;
wire  hea ;
wire  heb ;
wire  hec ;
wire  hed ;
wire  hfa ;
wire  hfb ;
wire  hfc ;
wire  hfd ;
wire  hga ;
wire  hgb ;
wire  hgc ;
wire  hgd ;
wire  hha ;
wire  hhb ;
wire  hhc ;
wire  hhd ;
wire  hia ;
wire  hib ;
wire  hic ;
wire  hid ;
wire  hja ;
wire  hjb ;
wire  hjc ;
wire  hjd ;
wire  hka ;
wire  hkb ;
wire  hkc ;
wire  hkd ;
wire  hla ;
wire  hlb ;
wire  hlc ;
wire  hld ;
wire  hma ;
wire  hmb ;
wire  hmc ;
wire  hmd ;
wire  hna ;
wire  hnb ;
wire  hnc ;
wire  hnd ;
wire  hoa ;
wire  hob ;
wire  hoc ;
wire  hod ;
wire  hpa ;
wire  hpb ;
wire  hpc ;
wire  hpd ;
wire  hqa ;
wire  hqb ;
wire  hqc ;
wire  hqd ;
wire  iaa ;
wire  iab ;
wire  iac ;
wire  iad ;
wire  iae ;
wire  iaf ;
wire  iag ;
wire  iah ;
wire  iai ;
wire  iaj ;
wire  iak ;
wire  ial ;
wire  iam ;
wire  ian ;
wire  iao ;
wire  iap ;
wire  iba ;
wire  ibb ;
wire  ibc ;
wire  ibd ;
wire  ibe ;
wire  ibf ;
wire  ibg ;
wire  ibh ;
wire  ibi ;
wire  ibj ;
wire  ibk ;
wire  ibl ;
wire  ibm ;
wire  ibn ;
wire  ibo ;
wire  ibp ;
wire  ica ;
wire  icb ;
wire  icc ;
wire  icd ;
wire  ice ;
wire  icf ;
wire  icg ;
wire  ich ;
wire  ici ;
wire  icj ;
wire  ick ;
wire  icl ;
wire  icm ;
wire  icn ;
wire  ico ;
wire  icp ;
wire  ida ;
wire  idb ;
wire  idc ;
wire  idd ;
wire  ide ;
wire  idf ;
wire  idg ;
wire  idh ;
wire  idi ;
wire  idj ;
wire  idk ;
wire  idl ;
wire  idm ;
wire  idn ;
wire  ido ;
wire  idp ;
wire  ifa ;
wire  ifb ;
wire  ifc ;
wire  ifd ;
wire  ife ;
wire  ifff  ;
wire  ifg ;
wire  ifh ;
wire  ifi ;
wire  ifj ;
wire  ifk ;
wire  ifl ;
wire  jaa ;
wire  JAA ;
wire  jab ;
wire  JAB ;
wire  jac ;
wire  JAC ;
wire  jad ;
wire  JAD ;
wire  jae ;
wire  JAE ;
wire  jaf ;
wire  JAF ;
wire  jag ;
wire  JAG ;
wire  jah ;
wire  JAH ;
wire  jai ;
wire  JAI ;
wire  jaj ;
wire  JAJ ;
wire  jak ;
wire  JAK ;
wire  jal ;
wire  JAL ;
wire  jam ;
wire  JAM ;
wire  jan ;
wire  JAN ;
wire  jao ;
wire  JAO ;
wire  jap ;
wire  JAP ;
wire  jba ;
wire  JBA ;
wire  jbb ;
wire  JBB ;
wire  jbc ;
wire  JBC ;
wire  jbd ;
wire  JBD ;
wire  jbe ;
wire  JBE ;
wire  jbf ;
wire  JBF ;
wire  jbg ;
wire  JBG ;
wire  jbh ;
wire  JBH ;
wire  jbi ;
wire  JBI ;
wire  jbj ;
wire  JBJ ;
wire  jbk ;
wire  JBK ;
wire  jbl ;
wire  JBL ;
wire  jbm ;
wire  JBM ;
wire  jbn ;
wire  JBN ;
wire  jbo ;
wire  JBO ;
wire  jbp ;
wire  JBP ;
wire  jca ;
wire  JCA ;
wire  jcb ;
wire  JCB ;
wire  jcc ;
wire  JCC ;
wire  jcd ;
wire  JCD ;
wire  jda ;
wire  JDA ;
wire  jdb ;
wire  JDB ;
wire  jdc ;
wire  JDC ;
wire  jdd ;
wire  JDD ;
wire  kaa ;
wire  kab ;
wire  kac ;
wire  kad ;
wire  kae ;
wire  kaf ;
wire  kag ;
wire  kah ;
wire  kai ;
wire  kaj ;
wire  kak ;
wire  kal ;
wire  kam ;
wire  kan ;
wire  kao ;
wire  kap ;
wire  kba ;
wire  kbb ;
wire  kbc ;
wire  kbd ;
wire  kbe ;
wire  kbf ;
wire  kbg ;
wire  kbh ;
wire  kbi ;
wire  kbj ;
wire  kbk ;
wire  kbl ;
wire  kbm ;
wire  kbn ;
wire  kbo ;
wire  kbp ;
wire  kka ;
wire  laa ;
wire  lab ;
wire  lac ;
wire  lad ;
wire  LAD ;
wire  lae ;
wire  laf ;
wire  lag ;
wire  lah ;
wire  lai ;
wire  laj ;
wire  lak ;
wire  lal ;
wire  lam ;
wire  lan ;
wire  lao ;
wire  lap ;
wire  lba ;
wire  lbb ;
wire  lbc ;
wire  lbd ;
wire  lbe ;
wire  lbf ;
wire  lbg ;
wire  lbh ;
wire  lbi ;
wire  lbj ;
wire  lbk ;
wire  lbl ;
wire  lbm ;
wire  lbn ;
wire  lbo ;
wire  lbp ;
wire  maa ;
wire  mab ;
wire  mac ;
wire  mad ;
wire  mae ;
wire  maf ;
wire  mag ;
wire  mah ;
wire  mai ;
wire  maj ;
wire  mak ;
wire  mal ;
wire  mam ;
wire  man ;
wire  mao ;
wire  map ;
wire  mba ;
wire  mbb ;
wire  mbc ;
wire  mbd ;
wire  mbe ;
wire  mbf ;
wire  mbg ;
wire  mbh ;
wire  mbi ;
wire  mbj ;
wire  mbk ;
wire  mbl ;
wire  mbm ;
wire  mbn ;
wire  mbo ;
wire  mbp ;
wire  naa ;
wire  NAA ;
wire  nab ;
wire  NAB ;
wire  nac ;
wire  NAC ;
wire  nad ;
wire  NAD ;
wire  nae ;
wire  NAE ;
wire  naf ;
wire  NAF ;
wire  nag ;
wire  NAG ;
wire  nah ;
wire  NAH ;
wire  nai ;
wire  NAI ;
wire  naj ;
wire  NAJ ;
wire  nak ;
wire  NAK ;
wire  nal ;
wire  NAL ;
wire  nam ;
wire  NAM ;
wire  nan ;
wire  NAN ;
wire  nao ;
wire  NAO ;
wire  nap ;
wire  NAP ;
wire  nba ;
wire  NBA ;
wire  nbb ;
wire  NBB ;
wire  nbc ;
wire  NBC ;
wire  nbd ;
wire  NBD ;
wire  nbe ;
wire  NBE ;
wire  nbf ;
wire  NBF ;
wire  nbg ;
wire  NBG ;
wire  nbh ;
wire  NBH ;
wire  nbi ;
wire  NBI ;
wire  nbj ;
wire  NBJ ;
wire  nbk ;
wire  NBK ;
wire  nbl ;
wire  NBL ;
wire  nbm ;
wire  NBM ;
wire  nbn ;
wire  NBN ;
wire  nbo ;
wire  NBO ;
wire  nbp ;
wire  NBP ;
wire  oaa ;
wire  oab ;
wire  oac ;
wire  oad ;
wire  oae ;
wire  oaf ;
wire  oag ;
wire  oah ;
wire  oai ;
wire  oaj ;
wire  oak ;
wire  oal ;
wire  oam ;
wire  oan ;
wire  oao ;
wire  oap ;
wire  oba ;
wire  obb ;
wire  obc ;
wire  obd ;
wire  obe ;
wire  obf ;
wire  obg ;
wire  obh ;
wire  obi ;
wire  obj ;
wire  obk ;
wire  obl ;
wire  obm ;
wire  obn ;
wire  obo ;
wire  obp ;
wire  oca ;
wire  ocb ;
wire  occ ;
wire  ocd ;
wire  oce ;
wire  ocf ;
wire  ocg ;
wire  och ;
wire  oci ;
wire  ocj ;
wire  ock ;
wire  ocl ;
wire  ocm ;
wire  ocn ;
wire  oco ;
wire  ocp ;
wire  oda ;
wire  odb ;
wire  odc ;
wire  odd ;
wire  ode ;
wire  odf ;
wire  odg ;
wire  odh ;
wire  odi ;
wire  odj ;
wire  odk ;
wire  odl ;
wire  odm ;
wire  odn ;
wire  odo ;
wire  odp ;
wire  OEA ;
wire  OEB ;
wire  oec ;
wire  qaa ;
wire  qab ;
wire  qac ;
wire  qad ;
wire  qae ;
wire  qaf ;
wire  qag ;
wire  qah ;
wire  qai ;
wire  qaj ;
wire  qak ;
wire  qal ;
wire  qap ;
wire  qaq ;
wire  qba ;
wire  qbb ;
wire  qbc ;
wire  qbd ;
wire  qbh ;
wire  qbi ;
wire  qbj ;
wire  qbk ;
wire  qbl ;
wire  qda ;
wire  qdb ;
wire  qdc ;
wire  QDD ;
wire  qea ;
wire  qeb ;
wire  qec ;
wire  qfa ;
wire  qfb ;
wire  qfc ;
wire  qfd ;
wire  qfe ;
wire  QFE ;
wire  qge ;
wire  TAA ;
wire  TAB ;
wire  tba ;
wire  tbb ;
wire  tca ;
wire  tcb ;
wire  tda ;
wire  tdb ;
wire  TEA ;
wire  TEB ;
wire  tfa ;
wire  tfb ;
wire  tga ;
wire  tgb ;
wire  tia ;
wire  tib ;
wire  tja ;
wire  tjb ;
wire  tla ;
wire  tlb ;
wire  tlc ;
wire  tma ;
wire  tmb ;
wire  tmc ;
wire  tna ;
wire  tnb ;
wire  toa ;
wire  tob ;
wire  tpa ;
wire  tpb ;
wire  tpc ;
wire  tpd ;
wire  tpe ;
wire  tpf ;
wire  tpg ;
wire  tph ;
wire  tqa ;
wire  tqb ;
wire  tqc ;
wire  tqd ;
wire  tqe ;
wire  tqf ;
wire  tqg ;
wire  tqh ;
wire  tra ;
wire  trb ;
wire  tsa ;
wire  tsb ;
wire  tsc ;
wire  tsd ;
wire  tta ;
wire  ttb ;
wire  ZZI ;
wire  ZZO ;
assign ZZI = 1'b1;
assign ZZO = 1'b0;
assign baa = ~BAA;  //complement 
assign bai = ~BAI;  //complement 
assign bba = ~BBA;  //complement 
assign bbi = ~BBI;  //complement 
assign bca = ~BCA;  //complement 
assign bcb = ~BCB;  //complement 
assign bcc = ~BCC;  //complement 
assign bcd = ~BCD;  //complement 
assign eaa = ~EAA;  //complement 
assign eab = ~EAB;  //complement 
assign eac = ~EAC;  //complement 
assign ead = ~EAD;  //complement 
assign maa = ~MAA;  //complement 
assign mai = ~MAI;  //complement 
assign mba = ~MBA;  //complement 
assign mbi = ~MBI;  //complement 
assign qaa = ~QAA;  //complement 
assign qab = ~QAB;  //complement 
assign qac = ~QAC;  //complement 
assign qad = ~QAD;  //complement 
assign qae = ~QAE;  //complement 
assign qaf = ~QAF;  //complement 
assign qag = ~QAG;  //complement 
assign qah = ~QAH;  //complement 
assign qai = ~QAI;  //complement 
assign qaj = ~QAJ;  //complement 
assign qak = ~QAK;  //complement 
assign qal = ~QAL;  //complement 
assign qda = ~QDA;  //complement 
assign qdb = ~QDB;  //complement 
assign qdc = ~QDC;  //complement 
assign NAA =  TOA & DAA  ; 
assign naa = ~NAA;  //complement 
assign NAB =  TOA & DAB  ; 
assign nab = ~NAB;  //complement 
assign NAC =  TOA & DAC  ; 
assign nac = ~NAC;  //complement 
assign NAD =  TOA & DAD  ; 
assign nad = ~NAD;  //complement 
assign NAE =  TOA & DAE  ; 
assign nae = ~NAE;  //complement 
assign NAF =  TOA & DAF  ; 
assign naf = ~NAF;  //complement 
assign NAG =  TOA & DAG  ; 
assign nag = ~NAG;  //complement 
assign NAH =  TOA & DAH  ; 
assign nah = ~NAH;  //complement 
assign NAI =  TOA & DAI  ; 
assign nai = ~NAI;  //complement 
assign NAJ =  TOA & DAJ  ; 
assign naj = ~NAJ;  //complement 
assign NAK =  TOA & DAK  ; 
assign nak = ~NAK;  //complement 
assign NAL =  TOA & DAL  ; 
assign nal = ~NAL;  //complement 
assign NAM =  TOA & DAM  ; 
assign nam = ~NAM;  //complement 
assign NAN =  TOA & DAN  ; 
assign nan = ~NAN;  //complement 
assign NAO =  TOA & DAO  ; 
assign nao = ~NAO;  //complement 
assign JCA =  BAA & BAB & BAC & BAD  ; 
assign jca = ~JCA;  //complement  
assign JCB =  BAE & BAF & BAG & BAH  ; 
assign jcb = ~JCB;  //complement 
assign JCC =  BAI & BAJ & BAK & BAL  ; 
assign jcc = ~JCC;  //complement  
assign JCD =  BAM & BAN & BAO & BAP  ; 
assign jcd = ~JCD;  //complement 
assign JDA =  BBA & BBB & BBC & BBD  ; 
assign jda = ~JDA;  //complement  
assign JDB =  BBE & BBF & BBG & BBH  ; 
assign jdb = ~JDB;  //complement 
assign JDC =  BBI & BBJ & BBK & BBL  ; 
assign jdc = ~JDC;  //complement  
assign JDD =  BBM & BBN & BBO & BBP  ; 
assign jdd = ~JDD;  //complement 
assign aaa = ~AAA;  //complement 
assign aai = ~AAI;  //complement 
assign aba = ~ABA;  //complement 
assign abi = ~ABI;  //complement 
assign NBD =  TOB & DBD  ; 
assign nbd = ~NBD;  //complement 
assign NBE =  TOB & DBE  ; 
assign nbe = ~NBE;  //complement 
assign NBF =  TOB & DBF  ; 
assign nbf = ~NBF;  //complement 
assign NBG =  TOB & DBG  ; 
assign nbg = ~NBG;  //complement 
assign NBH =  TOB & DBH  ; 
assign nbh = ~NBH;  //complement 
assign NBI =  TOB & DBI  ; 
assign nbi = ~NBI;  //complement 
assign NBJ =  TOB & DBJ  ; 
assign nbj = ~NBJ;  //complement 
assign NBK =  TOB & DBK  ; 
assign nbk = ~NBK;  //complement 
assign NBL =  TOB & DBL  ; 
assign nbl = ~NBL;  //complement 
assign NBM =  TOB & DBM  ; 
assign nbm = ~NBM;  //complement 
assign NBN =  TOB & DBN  ; 
assign nbn = ~NBN;  //complement 
assign NBO =  TOB & DBO  ; 
assign nbo = ~NBO;  //complement 
assign NAP =  TOA & DAP  ; 
assign nap = ~NAP;  //complement 
assign NBP =  TOB & DBP  ; 
assign nbp = ~NBP;  //complement 
assign NBA =  TOB & DBA  ; 
assign nba = ~NBA;  //complement 
assign NBB =  TOB & DBB  ; 
assign nbb = ~NBB;  //complement 
assign NBC =  TOB & DBC  ; 
assign nbc = ~NBC;  //complement 
assign EIA = ~eia;  //complement 
assign EIB = ~eib;  //complement 
assign EIC = ~eic;  //complement 
assign EID = ~eid;  //complement 
assign qea = ~QEA;  //complement 
assign qeb = ~QEB;  //complement 
assign qec = ~QEC;  //complement 
assign QDD = ~qdd;  //complement 
assign tba = ~TBA;  //complement 
assign tbb = ~TBB;  //complement 
assign tca = ~TCA;  //complement 
assign tcb = ~TCB;  //complement 
assign qfa = ~QFA;  //complement 
assign qfb = ~QFB;  //complement 
assign qfc = ~QFC;  //complement 
assign qfd = ~QFD;  //complement 
assign QFE =  IAE  ; 
assign qfe = ~QFE;  //complement 
assign qba = ~QBA;  //complement 
assign qbb = ~QBB;  //complement 
assign qbc = ~QBC;  //complement 
assign qbd = ~QBD;  //complement 
assign qbh = ~QBH;  //complement 
assign tfa = ~TFA;  //complement 
assign tfb = ~TFB;  //complement 
assign tga = ~TGA;  //complement 
assign tgb = ~TGB;  //complement 
assign JAA =  AAA & TPA  |  AAB & TPB  |  AAC & TPC  |  AAD & TPD  ; 
assign jaa = ~JAA;  //complement 
assign JAI =  AAI & TPA  |  AAJ & TPB  |  AAK & TPC  |  AAL & TPD  ; 
assign jai = ~JAI;  //complement 
assign JBA =  ABA & TPE  |  ABB & TPF  |  ABC & TPG  |  ABD & TPH  ; 
assign jba = ~JBA;  //complement 
assign JBI =  ABI & TPE  |  ABJ & TPF  |  ABK & TPG  |  ABL & TPH  ; 
assign jbi = ~JBI;  //complement 
assign kaa = ~KAA;  //complement 
assign kai = ~KAI;  //complement 
assign kba = ~KBA;  //complement 
assign kbi = ~KBI;  //complement 
assign ACA =  MAA & TIA  |  AAA & TJA  ; 
assign aca = ~ACA;  //complement 
assign ACI =  MAI & TIA  |  AAI & TJA  ; 
assign aci = ~ACI;  //complement 
assign ADA =  MBA & TIB  |  ABA & TJB  ; 
assign ada = ~ADA;  //complement 
assign ADI =  MBI & TIB  |  ABI & TJB  ; 
assign adi = ~ADI;  //complement 
assign tpe = ~TPE;  //complement 
assign tpf = ~TPF;  //complement 
assign tpg = ~TPG;  //complement 
assign tph = ~TPH;  //complement 
assign oaa = ~OAA;  //complement 
assign oai = ~OAI;  //complement 
assign oec = ~OEC;  //complement 
assign qap = ~QAP;  //complement 
assign qbi = ~QBI;  //complement 
assign qbj = ~QBJ;  //complement 
assign qbk = ~QBK;  //complement 
assign qbl = ~QBL;  //complement 
assign oba = ~OBA;  //complement 
assign obi = ~OBI;  //complement 
assign qaq = ~QAQ;  //complement 
assign OEA = ~oea;  //complement 
assign OEB = ~oeb;  //complement 
assign oca = ~OCA;  //complement 
assign oci = ~OCI;  //complement 
assign tia = ~TIA;  //complement 
assign tib = ~TIB;  //complement 
assign tja = ~TJA;  //complement 
assign tjb = ~TJB;  //complement 
assign tna = ~TNA;  //complement 
assign tnb = ~TNB;  //complement 
assign tsa = ~TSA;  //complement 
assign tsb = ~TSB;  //complement 
assign tsc = ~TSC;  //complement 
assign tsd = ~TSD;  //complement 
assign oda = ~ODA;  //complement 
assign odi = ~ODI;  //complement 
assign TAA = ~taa;  //complement 
assign qge = ~QGE;  //complement 
assign kka = ~KKA;  //complement 
assign TAB = ~tab;  //complement 
assign toa = ~TOA;  //complement 
assign tob = ~TOB;  //complement 
assign hak = ~HAK;  //complement 
assign tla = ~TLA;  //complement 
assign tlb = ~TLB;  //complement 
assign tlc = ~TLC;  //complement 
assign gah =  eia & eab & eac  |  eib & eac  |  eic  ; 
assign GAH = ~gah; //complement 
assign GAE =  EIA & EAB & EAC & EAD  |  EIB & EAC & EAD  |  EIC & EAD  |  EID  ; 
assign gae = ~GAE;  //complement 
assign GAD =  EIA & EAB & EAC  |  EIB & EAC  |  EIC  ; 
assign gad = ~GAD; //complement 
assign DAA = ZZO & ~aaa & ~baa  |  QDC & ~aaa & baa  |  QDB & aaa & ~baa  |  QDA & aaa & baa; 
assign daa = ~DAA;  //complement 
assign DAI = ZZO & ~aai & ~bai  |         QDC & ~aai & bai  |  QDB & aai & ~bai  |  QDA & aai & bai ; 
assign dai = ~DAI;  //complement 
assign DBA = ZZO & ~aba & ~bba  |  QEC & ~aba & bba  |  QEB & aba & ~bba  |  QEA & aba & bba; 
assign dba = ~DBA;  //complement 
assign DBI = ZZO & ~abi & ~bbi  |         QEC & ~abi & bbi  |  QEB & abi & ~bbi  |  QEA & abi & bbi ; 
assign dbi = ~DBI;  //complement 
assign laa = ~LAA;  //complement 
assign lab = ~LAB;  //complement 
assign lac = ~LAC;  //complement 
assign lba = ~LBA;  //complement 
assign lbb = ~LBB;  //complement 
assign lbc = ~LBC;  //complement 
assign tpa = ~TPA;  //complement 
assign tpb = ~TPB;  //complement 
assign tpc = ~TPC;  //complement 
assign tpd = ~TPD;  //complement 
assign eba = ~EBA;  //complement 
assign ebb = ~EBB;  //complement 
assign ebc = ~EBC;  //complement 
assign tra = ~TRA;  //complement 
assign trb = ~TRB;  //complement 
assign ebd = ~EBD;  //complement 
assign mab = ~MAB;  //complement 
assign maj = ~MAJ;  //complement 
assign mbb = ~MBB;  //complement 
assign mbj = ~MBJ;  //complement 
assign tda = ~TDA;  //complement 
assign tdb = ~TDB;  //complement 
assign gbh =  eja & ebb & ebc  |  ejb & ebc  |  ejc  ; 
assign GBH = ~gbh; //complement 
assign gch =  eka & ecb & ecc  |  ekb & ecc  |  ekc  ; 
assign GCH = ~gch; //complement 
assign gdh =  ela & edb & edc  |  elb & edc  |  elc  ; 
assign GDH = ~gdh; //complement 
assign geh =  ema & eeb & eec  |  emb & eec  |  emc  ; 
assign GEH = ~geh; //complement 
assign gfh =  ena & efb & efc  |  enb & efc  |  enc  ; 
assign GFH = ~gfh; //complement 
assign ggh =  eoa & egb & egc  |  eob & egc  |  eoc  ; 
assign GGH = ~ggh; //complement 
assign ghh =  epa & ehb & ehc  |  epb & ehc  |  epc  ; 
assign GHH = ~ghh; //complement 
assign hac = ~HAC;  //complement 
assign had = ~HAD;  //complement 
assign tma = ~TMA;  //complement 
assign tmb = ~TMB;  //complement 
assign tmc = ~TMC;  //complement 
assign gag =  eia & eab  |  eib  ; 
assign GAG = ~gag;  //complement 
assign gcg =  eka & ecb  |  ekb  ; 
assign GCG = ~gcg;  //complement 
assign geg =  ema & eeb  |  emb  ; 
assign GEG = ~geg;  //complement 
assign ggg =  eoa & egb  |  eob  ; 
assign GGG = ~ggg;  //complement 
assign aab = ~AAB;  //complement 
assign aaj = ~AAJ;  //complement 
assign abb = ~ABB;  //complement 
assign abj = ~ABJ;  //complement 
assign bab = ~BAB;  //complement 
assign baj = ~BAJ;  //complement 
assign bbb = ~BBB;  //complement 
assign bbj = ~BBJ;  //complement 
assign EJA = ~eja;  //complement 
assign EJB = ~ejb;  //complement 
assign EJC = ~ejc;  //complement 
assign EJD = ~ejd;  //complement 
assign TEA = ~tea;  //complement 
assign TEB = ~teb;  //complement 
assign GAB =  EIA  ; 
assign gab = ~GAB;  //complement 
assign GBB =  EJA  ; 
assign gbb = ~GBB;  //complement 
assign GCB =  EKA  ; 
assign gcb = ~GCB;  //complement 
assign GDB =  ELA  ; 
assign gdb = ~GDB;  //complement 
assign GEB =  EMA  ; 
assign geb = ~GEB;  //complement 
assign GFB =  ENA  ; 
assign gfb = ~GFB;  //complement 
assign GHB =  EPA  ; 
assign ghb = ~GHB;  //complement 
assign GGB =  EOA  ; 
assign ggb = ~GGB;  //complement 
assign gaf =  eia  ; 
assign GAF = ~gaf;  //complement 
assign gbf =  eja  ; 
assign GBF = ~gbf;  //complement 
assign gcf =  eka  ; 
assign GCF = ~gcf;  //complement 
assign gdf =  ela  ; 
assign GDF = ~gdf;  //complement 
assign gef =  ema  ; 
assign GEF = ~gef;  //complement 
assign gff =  ena  ; 
assign GFF = ~gff;  //complement 
assign ggf =  eoa  ; 
assign GGF = ~ggf;  //complement 
assign ghf =  epa  ; 
assign GHF = ~ghf;  //complement 
assign hae = ~HAE;  //complement 
assign HAF = ~haf;  //complement 
assign JAB =  AAB & TPA  |  AAC & TPB  |  AAD & TPC  |  AAE & TPD  ; 
assign jab = ~JAB;  //complement 
assign JAJ =  AAJ & TPA  |  AAK & TPB  |  AAL & TPC  |  AAM & TPD  ; 
assign jaj = ~JAJ;  //complement 
assign JBB =  ABB & TPE  |  ABC & TPF  |  ABD & TPG  |  ABE & TPH  ; 
assign jbb = ~JBB;  //complement 
assign JBJ =  ABJ & TPE  |  ABK & TPF  |  ABL & TPG  |  ABM & TPH  ; 
assign jbj = ~JBJ;  //complement 
assign kab = ~KAB;  //complement 
assign kaj = ~KAJ;  //complement 
assign kbb = ~KBB;  //complement 
assign kbj = ~KBJ;  //complement 
assign ACB =  MAB & TIA  |  AAB & TJA  ; 
assign acb = ~ACB;  //complement 
assign ACJ =  MAJ & TIA  |  AAJ & TJA  ; 
assign acj = ~ACJ;  //complement 
assign ADB =  MBB & TIB  |  ABB & TJB  ; 
assign adb = ~ADB;  //complement 
assign ADJ =  MBJ & TIB  |  ABJ & TJB  ; 
assign adj = ~ADJ;  //complement 
assign tqc = ~TQC;  //complement 
assign tqd = ~TQD;  //complement 
assign tqe = ~TQE;  //complement 
assign tqf = ~TQF;  //complement 
assign tqh = ~TQH;  //complement 
assign tqg = ~TQG;  //complement 
assign oab = ~OAB;  //complement 
assign oaj = ~OAJ;  //complement 
assign lbd = ~LBD;  //complement 
assign haa = ~HAA;  //complement 
assign hba = ~HBA;  //complement 
assign hca = ~HCA;  //complement 
assign hda = ~HDA;  //complement 
assign hab = ~HAB;  //complement 
assign obb = ~OBB;  //complement 
assign obj = ~OBJ;  //complement 
assign hea = ~HEA;  //complement 
assign hfa = ~HFA;  //complement 
assign hga = ~HGA;  //complement 
assign hha = ~HHA;  //complement 
assign hbb = ~HBB;  //complement 
assign hbc = ~HBC;  //complement 
assign ocb = ~OCB;  //complement 
assign ocj = ~OCJ;  //complement 
assign hbd = ~HBD;  //complement 
assign hcb = ~HCB;  //complement 
assign hcc = ~HCC;  //complement 
assign odb = ~ODB;  //complement 
assign odj = ~ODJ;  //complement 
assign hcd = ~HCD;  //complement 
assign hhb = ~HHB;  //complement 
assign hhc = ~HHC;  //complement 
assign hhd = ~HHD;  //complement 
assign hag = ~HAG;  //complement 
assign GBE =  EJA & EBB & EBC & EBD  |  EJB & EBC & EBD  |  EJC & EBD  |  EJD  ; 
assign gbe = ~GBE;  //complement 
assign GBD =  EJA & EBB & EBC  |  EJB & EBC  |  EJC  ; 
assign gbd = ~GBD; //complement 
assign DAB = ZZO & ~aab & ~bab  |  QDC & ~aab & bab  |  QDB & aab & ~bab  |  QDA & aab & bab; 
assign dab = ~DAB;  //complement 
assign DAJ = ZZO & ~aaj & ~baj  |         QDC & ~aaj & baj  |  QDB & aaj & ~baj  |  QDA & aaj & baj ; 
assign daj = ~DAJ;  //complement 
assign DBB = ZZO & ~abb & ~bbb  |  QEC & ~abb & bbb  |  QEB & abb & ~bbb  |  QEA & abb & bbb; 
assign dbb = ~DBB;  //complement 
assign DBJ = ZZO & ~abj & ~bbj  |         QEC & ~abj & bbj  |  QEB & abj & ~bbj  |  QEA & abj & bbj ; 
assign dbj = ~DBJ;  //complement 
assign lae = ~LAE;  //complement 
assign laf = ~LAF;  //complement 
assign lbe = ~LBE;  //complement 
assign lbf = ~LBF;  //complement 
assign LAD =  HBD & qbb  |  HJD & QBB  ; 
assign lad = ~LAD;  //complement 
assign tqa = ~TQA;  //complement 
assign tqb = ~TQB;  //complement 
assign bbc = ~BBC;  //complement 
assign bbk = ~BBK;  //complement 
assign eca = ~ECA;  //complement 
assign bda = ~BDA;  //complement 
assign bdb = ~BDB;  //complement 
assign bdc = ~BDC;  //complement 
assign bdd = ~BDD;  //complement 
assign ecb = ~ECB;  //complement 
assign ecc = ~ECC;  //complement 
assign ecd = ~ECD;  //complement 
assign mac = ~MAC;  //complement 
assign mak = ~MAK;  //complement 
assign mbc = ~MBC;  //complement 
assign mbk = ~MBK;  //complement 
assign GMA =  EFA & EFB & EFC & EFD  ; 
assign gma = ~GMA;  //complement  
assign GNA =  EGA & EGB & EGC & EGD  ; 
assign gna = ~GNA;  //complement 
assign GPA =  EDA & EDB & EDC & EDD & EEA & EEB  ; 
assign gpa = ~GPA;  //complement  
assign aac = ~AAC;  //complement 
assign aak = ~AAK;  //complement 
assign abc = ~ABC;  //complement 
assign abk = ~ABK;  //complement 
assign bac = ~BAC;  //complement 
assign GIA =  EBA & EBB & EBC & EBD  ; 
assign gia = ~GIA;  //complement  
assign GJA =  ECA & ECB & ECC & ECD  ; 
assign gja = ~GJA;  //complement 
assign GKA =  EDA & EDB & EDC & EDD  ; 
assign gka = ~GKA;  //complement  
assign GLA =  EEA & EEB & EEC & EED  ; 
assign gla = ~GLA;  //complement 
assign bak = ~BAK;  //complement 
assign EKA = ~eka;  //complement 
assign EKB = ~ekb;  //complement 
assign EKC = ~ekc;  //complement 
assign EKD = ~ekd;  //complement 
assign GAC =  EIA & EAB  |  EAB  ; 
assign gac = ~GAC;  //complement 
assign GCC =  EKA & ECB  |  EKB  ; 
assign gcc = ~GCC;  //complement 
assign GEC =  EMA & EEB  |  EMB  ; 
assign gec = ~GEC;  //complement 
assign GGC =  EOA & EGB  |  EOB  ; 
assign ggc = ~GGC;  //complement 
assign tta = ~TTA;  //complement 
assign ttb = ~TTB;  //complement 
assign hia = ~HIA;  //complement 
assign hja = ~HJA;  //complement 
assign hka = ~HKA;  //complement 
assign hla = ~HLA;  //complement 
assign hma = ~HMA;  //complement 
assign hna = ~HNA;  //complement 
assign hoa = ~HOA;  //complement 
assign hpa = ~HPA;  //complement 
assign hqa = ~HQA;  //complement 
assign hqb = ~HQB;  //complement 
assign hqc = ~HQC;  //complement 
assign JAC =  AAC & TPA  |  AAD & TPB  |  AAE & TPC  |  AAF & TPD  ; 
assign jac = ~JAC;  //complement 
assign hqd = ~HQD;  //complement 
assign JAK =  AAK & TPA  |  AAL & TPB  |  AAM & TPC  |  AAN & TPD  ; 
assign jak = ~JAK;  //complement 
assign JBC =  ABC & TPE  |  ABD & TPF  |  ABE & TPG  |  ABF & TPH  ; 
assign jbc = ~JBC;  //complement 
assign JBK =  ABK & TPE  |  ABL & TPF  |  ABM & TPG  |  ABN & TPH  ; 
assign jbk = ~JBK;  //complement 
assign kac = ~KAC;  //complement 
assign kak = ~KAK;  //complement 
assign kbc = ~KBC;  //complement 
assign kbk = ~KBK;  //complement 
assign ACC =  MAC & TIA  |  AAC & TJA  ; 
assign acc = ~ACC;  //complement 
assign ACK =  MAK & TIA  |  AAK & TJA  ; 
assign ack = ~ACK;  //complement 
assign ADC =  MBC & TIB  |  ABC & TJB  ; 
assign adc = ~ADC;  //complement 
assign ADK =  MBK & TIB  |  ABK & TJB  ; 
assign adk = ~ADK;  //complement 
assign lbj = ~LBJ;  //complement 
assign laj = ~LAJ;  //complement 
assign lak = ~LAK;  //complement 
assign lal = ~LAL;  //complement 
assign HAH = ~hah;  //complement 
assign oac = ~OAC;  //complement 
assign oak = ~OAK;  //complement 
assign lai = ~LAI;  //complement 
assign lbk = ~LBK;  //complement 
assign lbl = ~LBL;  //complement 
assign obc = ~OBC;  //complement 
assign obk = ~OBK;  //complement 
assign hdb = ~HDB;  //complement 
assign hdc = ~HDC;  //complement 
assign hdd = ~HDD;  //complement 
assign occ = ~OCC;  //complement 
assign ock = ~OCK;  //complement 
assign GQA =  EEC & EED & EFA & EFB & EFC & EFD  ; 
assign gqa = ~GQA;  //complement  
assign HAI = ~hai;  //complement 
assign haj = ~HAJ;  //complement 
assign odc = ~ODC;  //complement 
assign odk = ~ODK;  //complement 
assign GBC =  EJA & EBB  |  EJB  ; 
assign gbc = ~GBC;  //complement 
assign GDC =  ELA & EDB  |  ELB  ; 
assign gdc = ~GDC;  //complement 
assign GFC =  ENA & EFB  |  ENB  ; 
assign gfc = ~GFC;  //complement 
assign GHC =  EPA & EHB  |  EPB  ; 
assign ghc = ~GHC;  //complement 
assign gbg =  eja & ebb  |  ejb  ; 
assign GBG = ~gbg;  //complement 
assign gdg =  ela & edb  |  elb  ; 
assign GDG = ~gdg;  //complement 
assign gfg =  ena & efb  |  enb  ; 
assign GFG = ~gfg;  //complement 
assign GCE =  EKA & ECB & ECC & ECD  |  EKB & ECC & ECD  |  EKC & ECD  |  EKD  ; 
assign gce = ~GCE;  //complement 
assign GCD =  EKA & ECB & ECC  |  EKB & ECC  |  EKC  ; 
assign gcd = ~GCD; //complement 
assign DAC = ZZO & ~aac & ~bac  |  QDC & ~aac & bac  |  QDB & aac & ~bac  |  QDA & aac & bac; 
assign dac = ~DAC;  //complement 
assign DAK = ZZO & ~aak & ~bak  |         QDC & ~aak & bak  |  QDB & aak & ~bak  |  QDA & aak & bak ; 
assign dak = ~DAK;  //complement 
assign DBC = ZZO & ~abc & ~bbc  |  QEC & ~abc & bbc  |  QEB & abc & ~bbc  |  QEA & abc & bbc; 
assign dbc = ~DBC;  //complement 
assign DBK = ZZO & ~abk & ~bbk  |         QEC & ~abk & bbk  |  QEB & abk & ~bbk  |  QEA & abk & bbk ; 
assign dbk = ~DBK;  //complement 
assign lag = ~LAG;  //complement 
assign lah = ~LAH;  //complement 
assign lbg = ~LBG;  //complement 
assign lbh = ~LBH;  //complement 
assign lbi = ~LBI;  //complement 
assign eda = ~EDA;  //complement 
assign edb = ~EDB;  //complement 
assign edc = ~EDC;  //complement 
assign bde = ~BDE;  //complement 
assign bdf = ~BDF;  //complement 
assign bdg = ~BDG;  //complement 
assign bdh = ~BDH;  //complement 
assign edd = ~EDD;  //complement 
assign mad = ~MAD;  //complement 
assign mal = ~MAL;  //complement 
assign mbd = ~MBD;  //complement 
assign mbl = ~MBL;  //complement 
assign ghg =  epa & ehb  |  epb  ; 
assign GHG = ~ghg;  //complement 
assign aad = ~AAD;  //complement 
assign aal = ~AAL;  //complement 
assign abd = ~ABD;  //complement 
assign abl = ~ABL;  //complement 
assign bad = ~BAD;  //complement 
assign bal = ~BAL;  //complement 
assign bbd = ~BBD;  //complement 
assign bbl = ~BBL;  //complement 
assign ELA = ~ela;  //complement 
assign ELB = ~elb;  //complement 
assign ELC = ~elc;  //complement 
assign ELD = ~eld;  //complement 
assign JAD =  AAD & TPA  |  AAE & TPB  |  AAF & TPC  |  AAG & TPD  ; 
assign jad = ~JAD;  //complement 
assign JAL =  AAL & TPA  |  AAM & TPB  |  AAN & TPC  |  AAO & TPD  ; 
assign jal = ~JAL;  //complement 
assign JBD =  ABD & TPE  |  ABE & TPF  |  ABF & TPG  |  ABG & TPH  ; 
assign jbd = ~JBD;  //complement 
assign JBL =  ABL & TPE  |  ABM & TPF  |  ABN & TPG  |  ABO & TPH  ; 
assign jbl = ~JBL;  //complement 
assign kad = ~KAD;  //complement 
assign kal = ~KAL;  //complement 
assign kbd = ~KBD;  //complement 
assign kbl = ~KBL;  //complement 
assign ACD =  MAD & TIA  |  AAD & TJA  ; 
assign acd = ~ACD;  //complement 
assign ACL =  MAL & TIA  |  AAL & TJA  ; 
assign acl = ~ACL;  //complement 
assign ADD =  MBD & TIB  |  ABD & TJB  ; 
assign add = ~ADD;  //complement 
assign ADL =  MBL & TIB  |  ABL & TJB  ; 
assign adl = ~ADL;  //complement 
assign oad = ~OAD;  //complement 
assign oal = ~OAL;  //complement 
assign obd = ~OBD;  //complement 
assign obl = ~OBL;  //complement 
assign ocd = ~OCD;  //complement 
assign ocl = ~OCL;  //complement 
assign odd = ~ODD;  //complement 
assign odl = ~ODL;  //complement 
assign GDE =  ELA & EDB & EDC & EDD  |  ELB & EDC & EDD  |  ELC & EDD  |  ELD  ; 
assign gde = ~GDE;  //complement 
assign GDD =  ELA & EDB & EDC  |  ELB & EDC  |  ELC  ; 
assign gdd = ~GDD; //complement 
assign DAD = ZZO & ~aad & ~bad  |  QDC & ~aad & bad  |  QDB & aad & ~bad  |  QDA & aad & bad; 
assign dad = ~DAD;  //complement 
assign DAL = ZZO & ~aal & ~bal  |         QDC & ~aal & bal  |  QDB & aal & ~bal  |  QDA & aal & bal ; 
assign dal = ~DAL;  //complement 
assign DBD = ZZO & ~abd & ~bbd  |  QEC & ~abd & bbd  |  QEB & abd & ~bbd  |  QEA & abd & bbd; 
assign dbd = ~DBD;  //complement 
assign DBL = ZZO & ~abl & ~bbl  |         QEC & ~abl & bbl  |  QEB & abl & ~bbl  |  QEA & abl & bbl ; 
assign dbl = ~DBL;  //complement 
assign heb = ~HEB;  //complement 
assign hec = ~HEC;  //complement 
assign hed = ~HED;  //complement 
assign eea = ~EEA;  //complement 
assign eeb = ~EEB;  //complement 
assign eec = ~EEC;  //complement 
assign bce = ~BCE;  //complement 
assign bcf = ~BCF;  //complement 
assign bcg = ~BCG;  //complement 
assign bch = ~BCH;  //complement 
assign eed = ~EED;  //complement 
assign mae = ~MAE;  //complement 
assign mam = ~MAM;  //complement 
assign mbe = ~MBE;  //complement 
assign mbm = ~MBM;  //complement 
assign aae = ~AAE;  //complement 
assign aam = ~AAM;  //complement 
assign abe = ~ABE;  //complement 
assign abm = ~ABM;  //complement 
assign bae = ~BAE;  //complement 
assign bam = ~BAM;  //complement 
assign bbe = ~BBE;  //complement 
assign bbm = ~BBM;  //complement 
assign EMA = ~ema;  //complement 
assign EMB = ~emb;  //complement 
assign EMC = ~emc;  //complement 
assign EMD = ~emd;  //complement 
assign hfb = ~HFB;  //complement 
assign hfc = ~HFC;  //complement 
assign hfd = ~HFD;  //complement 
assign JAE =  AAE & TPA  |  AAF & TPB  |  AAG & TPC  |  AAH & TPD  ; 
assign jae = ~JAE;  //complement 
assign JAM =  AAM & TPA  |  AAN & TPB  |  AAO & TPC  |  AAP & TPD  ; 
assign jam = ~JAM;  //complement 
assign JBE =  ABE & TPE  |  ABF & TPF  |  ABG & TPG  |  ABH & TPH  ; 
assign jbe = ~JBE;  //complement 
assign JBM =  ABM & TPE  |  ABN & TPF  |  ABO & TPG  |  ABP & TPH  ; 
assign jbm = ~JBM;  //complement 
assign kae = ~KAE;  //complement 
assign kam = ~KAM;  //complement 
assign kbe = ~KBE;  //complement 
assign kbm = ~KBM;  //complement 
assign ACE =  MAE & TIA  |  AAE & TJA  ; 
assign ace = ~ACE;  //complement 
assign ACM =  MAM & TIA  |  AAM & TJA  ; 
assign acm = ~ACM;  //complement 
assign ADE =  MBE & TIB  |  ABE & TJB  ; 
assign ade = ~ADE;  //complement 
assign ADM =  MBM & TIB  |  ABM & TJB  ; 
assign adm = ~ADM;  //complement 
assign oae = ~OAE;  //complement 
assign oam = ~OAM;  //complement 
assign obe = ~OBE;  //complement 
assign obm = ~OBM;  //complement 
assign oce = ~OCE;  //complement 
assign ocm = ~OCM;  //complement 
assign ode = ~ODE;  //complement 
assign odm = ~ODM;  //complement 
assign GEE =  EMA & EEB & EEC & EED  |  EMB & EEC & EED  |  EMC & EED  |  EMD  ; 
assign gee = ~GEE;  //complement 
assign GED =  EMA & EEB & EEC  |  EMB & EEC  |  EMC  ; 
assign ged = ~GED; //complement 
assign DAE = ZZO & ~aae & ~bae  |  QDC & ~aae & bae  |  QDB & aae & ~bae  |  QDA & aae & bae; 
assign dae = ~DAE;  //complement 
assign DAM = ZZO & ~aam & ~bam  |         QDC & ~aam & bam  |  QDB & aam & ~bam  |  QDA & aam & bam ; 
assign dam = ~DAM;  //complement 
assign DBE = ZZO & ~abe & ~bbe  |  QEC & ~abe & bbe  |  QEB & abe & ~bbe  |  QEA & abe & bbe; 
assign dbe = ~DBE;  //complement 
assign DBM = ZZO & ~abm & ~bbm  |         QEC & ~abm & bbm  |  QEB & abm & ~bbm  |  QEA & abm & bbm ; 
assign dbm = ~DBM;  //complement 
assign lam = ~LAM;  //complement 
assign lan = ~LAN;  //complement 
assign lao = ~LAO;  //complement 
assign lbm = ~LBM;  //complement 
assign lbn = ~LBN;  //complement 
assign lbo = ~LBO;  //complement 
assign lap = ~LAP;  //complement 
assign lbp = ~LBP;  //complement 
assign efa = ~EFA;  //complement 
assign efb = ~EFB;  //complement 
assign efc = ~EFC;  //complement 
assign bci = ~BCI;  //complement 
assign bcj = ~BCJ;  //complement 
assign bck = ~BCK;  //complement 
assign bcl = ~BCL;  //complement 
assign efd = ~EFD;  //complement 
assign maf = ~MAF;  //complement 
assign man = ~MAN;  //complement 
assign mbf = ~MBF;  //complement 
assign mbn = ~MBN;  //complement 
assign aaf = ~AAF;  //complement 
assign aan = ~AAN;  //complement 
assign abf = ~ABF;  //complement 
assign abn = ~ABN;  //complement 
assign baf = ~BAF;  //complement 
assign ban = ~BAN;  //complement 
assign bbf = ~BBF;  //complement 
assign bbn = ~BBN;  //complement 
assign ENA = ~ena;  //complement 
assign ENB = ~enb;  //complement 
assign ENC = ~enc;  //complement 
assign ENDD  = ~endd;  //complement 
assign hib = ~HIB;  //complement 
assign hic = ~HIC;  //complement 
assign hid = ~HID;  //complement 
assign hjb = ~HJB;  //complement 
assign hjc = ~HJC;  //complement 
assign hjd = ~HJD;  //complement 
assign hkb = ~HKB;  //complement 
assign hkc = ~HKC;  //complement 
assign hkd = ~HKD;  //complement 
assign hlb = ~HLB;  //complement 
assign hlc = ~HLC;  //complement 
assign hld = ~HLD;  //complement 
assign JAF =  AAF & TPA  |  AAG & TPB  |  AAH & TPC  |  AAI & TPD  ; 
assign jaf = ~JAF;  //complement 
assign JAN =  AAN & TPA  |  AAO & TPB  |  AAP & TPC  |  ABA & TPD  ; 
assign jan = ~JAN;  //complement 
assign JBF =  ABF & TPE  |  ABG & TPF  |  ABH & TPG  |  ABI & TPH  ; 
assign jbf = ~JBF;  //complement 
assign JBN =  ABN & TPE  |  ABO & TPF  |  ABP & TPG  ; 
assign jbn = ~JBN;  //complement 
assign kaf = ~KAF;  //complement 
assign kan = ~KAN;  //complement 
assign kbf = ~KBF;  //complement 
assign kbn = ~KBN;  //complement 
assign ACF =  MAF & TIA  |  AAF & TJA  ; 
assign acf = ~ACF;  //complement 
assign ACN =  MAN & TIA  |  AAN & TJA  ; 
assign acn = ~ACN;  //complement 
assign ADF =  MBF & TIB  |  ABF & TJB  ; 
assign adf = ~ADF;  //complement 
assign ADN =  MBN & TIB  |  ABN & TJB  ; 
assign adn = ~ADN;  //complement 
assign oaf = ~OAF;  //complement 
assign oan = ~OAN;  //complement 
assign obf = ~OBF;  //complement 
assign obn = ~OBN;  //complement 
assign ocf = ~OCF;  //complement 
assign ocn = ~OCN;  //complement 
assign odf = ~ODF;  //complement 
assign odn = ~ODN;  //complement 
assign GFE =  ENA & EFB & EFC & EFD  |  ENB & EFC & EFD  |  ENC & EFD  |  ENDD   ; 
assign gfe = ~GFE;  //complement 
assign GFD =  ENA & EFB & EFC  |  ENB & EFC  |  ENC  ; 
assign gfd = ~GFD; //complement 
assign DAF = ZZO & ~aaf & ~baf  |  QDC & ~aaf & baf  |  QDB & aaf & ~baf  |  QDA & aaf & baf; 
assign daf = ~DAF;  //complement 
assign DAN = ZZO & ~aan & ~ban  |         QDC & ~aan & ban  |  QDB & aan & ~ban  |  QDA & aan & ban ; 
assign dan = ~DAN;  //complement 
assign DBF = ZZO & ~abf & ~bbf  |  QEC & ~abf & bbf  |  QEB & abf & ~bbf  |  QEA & abf & bbf; 
assign dbf = ~DBF;  //complement 
assign DBN = ZZO & ~abn & ~bbn  |         QEC & ~abn & bbn  |  QEB & abn & ~bbn  |  QEA & abn & bbn ; 
assign dbn = ~DBN;  //complement 
assign hgb = ~HGB;  //complement 
assign hgc = ~HGC;  //complement 
assign hgd = ~HGD;  //complement 
assign ega = ~EGA;  //complement 
assign egb = ~EGB;  //complement 
assign egc = ~EGC;  //complement 
assign bcm = ~BCM;  //complement 
assign bcn = ~BCN;  //complement 
assign bco = ~BCO;  //complement 
assign bcp = ~BCP;  //complement 
assign egd = ~EGD;  //complement 
assign mag = ~MAG;  //complement 
assign mao = ~MAO;  //complement 
assign mbg = ~MBG;  //complement 
assign mbo = ~MBO;  //complement 
assign aag = ~AAG;  //complement 
assign aao = ~AAO;  //complement 
assign abg = ~ABG;  //complement 
assign abo = ~ABO;  //complement 
assign bag = ~BAG;  //complement 
assign bao = ~BAO;  //complement 
assign bbg = ~BBG;  //complement 
assign bbo = ~BBO;  //complement 
assign EOA = ~eoa;  //complement 
assign EOB = ~eob;  //complement 
assign EOC = ~eoc;  //complement 
assign EOD = ~eod;  //complement 
assign JAG =  AAG & TPA  |  AAH & TPB  |  AAI & TPC  |  AAJ & TPD  ; 
assign jag = ~JAG;  //complement 
assign JAO =  AAO & TPA  |  AAP & TPB  |  ABA & TPC  |  ABB & TPD  ; 
assign jao = ~JAO;  //complement 
assign JBG =  ABG & TPE  |  ABH & TPF  |  ABI & TPG  |  ABJ & TPH  ; 
assign jbg = ~JBG;  //complement 
assign JBO =  ABO & TPE  |  ABP & TPF  ; 
assign jbo = ~JBO;  //complement 
assign kag = ~KAG;  //complement 
assign kao = ~KAO;  //complement 
assign kbg = ~KBG;  //complement 
assign kbo = ~KBO;  //complement 
assign ACG =  MAG & TIA  |  AAG & TJA  ; 
assign acg = ~ACG;  //complement 
assign ACO =  MAO & TIA  |  AAO & TJA  ; 
assign aco = ~ACO;  //complement 
assign ADG =  MBG & TIB  |  ABG & TJB  ; 
assign adg = ~ADG;  //complement 
assign ADO =  MBO & TIB  |  ABO & TJB  ; 
assign ado = ~ADO;  //complement 
assign oag = ~OAG;  //complement 
assign oao = ~OAO;  //complement 
assign obg = ~OBG;  //complement 
assign obo = ~OBO;  //complement 
assign ocg = ~OCG;  //complement 
assign oco = ~OCO;  //complement 
assign odg = ~ODG;  //complement 
assign odo = ~ODO;  //complement 
assign GGE =  EOA & EGB & EGC & EGD  |  EOB & EGC & EGD  |  EOC & EGD  |  EOD  ; 
assign gge = ~GGE;  //complement 
assign GGD =  EOA & EGB & EGC  |  EOB & EGC  |  EOC  ; 
assign ggd = ~GGD; //complement 
assign DAG = ZZO & ~aag & ~bag  |  QDC & ~aag & bag  |  QDB & aag & ~bag  |  QDA & aag & bag; 
assign dag = ~DAG;  //complement 
assign DAO = ZZO & ~aao & ~bao  |         QDC & ~aao & bao  |  QDB & aao & ~bao  |  QDA & aao & bao ; 
assign dao = ~DAO;  //complement 
assign DBG = ZZO & ~abg & ~bbg  |  QEC & ~abg & bbg  |  QEB & abg & ~bbg  |  QEA & abg & bbg; 
assign dbg = ~DBG;  //complement 
assign DBO = ZZO & ~abo & ~bbo  |         QEC & ~abo & bbo  |  QEB & abo & ~bbo  |  QEA & abo & bbo ; 
assign dbo = ~DBO;  //complement 
assign eha = ~EHA;  //complement 
assign ehb = ~EHB;  //complement 
assign ehc = ~EHC;  //complement 
assign bdi = ~BDI;  //complement 
assign bdj = ~BDJ;  //complement 
assign bdk = ~BDK;  //complement 
assign bdl = ~BDL;  //complement 
assign ehd = ~EHD;  //complement 
assign mah = ~MAH;  //complement 
assign map = ~MAP;  //complement 
assign mbh = ~MBH;  //complement 
assign mbp = ~MBP;  //complement 
assign bdm = ~BDM;  //complement 
assign bdn = ~BDN;  //complement 
assign bdo = ~BDO;  //complement 
assign bdp = ~BDP;  //complement 
assign aah = ~AAH;  //complement 
assign aap = ~AAP;  //complement 
assign abh = ~ABH;  //complement 
assign abp = ~ABP;  //complement 
assign bah = ~BAH;  //complement 
assign bap = ~BAP;  //complement 
assign bbh = ~BBH;  //complement 
assign bbp = ~BBP;  //complement 
assign EPA = ~epa;  //complement 
assign EPB = ~epb;  //complement 
assign EPC = ~epc;  //complement 
assign EPD = ~epd;  //complement 
assign JAH =  AAH & TPA  |  AAI & TPB  |  AAJ & TPC  |  AAK & TPD  ; 
assign jah = ~JAH;  //complement 
assign JAP =  AAP & TPA  |  ABA & TPB  |  ABB & TPC  |  ABC & TPD  ; 
assign jap = ~JAP;  //complement 
assign JBH =  ABH & TPE  |  ABI & TPF  |  ABJ & TPG  |  ABK & TPH  ; 
assign jbh = ~JBH;  //complement 
assign JBP =  ABP & TPE  ; 
assign jbp = ~JBP;  //complement 
assign kah = ~KAH;  //complement 
assign kap = ~KAP;  //complement 
assign kbh = ~KBH;  //complement 
assign kbp = ~KBP;  //complement 
assign ACH =  MAH & TIA  |  AAH & TJA  ; 
assign ach = ~ACH;  //complement 
assign ACP =  MAP & TIA  |  AAP & TJA  ; 
assign acp = ~ACP;  //complement 
assign ADH =  MBH & TIB  |  ABH & TJB  ; 
assign adh = ~ADH;  //complement 
assign ADP =  MBP & TIB  |  ABP & TJB  ; 
assign adp = ~ADP;  //complement 
assign hnc = ~HNC;  //complement 
assign hnd = ~HND;  //complement 
assign hob = ~HOB;  //complement 
assign oah = ~OAH;  //complement 
assign oap = ~OAP;  //complement 
assign hoc = ~HOC;  //complement 
assign hod = ~HOD;  //complement 
assign hpb = ~HPB;  //complement 
assign obh = ~OBH;  //complement 
assign obp = ~OBP;  //complement 
assign hpc = ~HPC;  //complement 
assign hpd = ~HPD;  //complement 
assign och = ~OCH;  //complement 
assign ocp = ~OCP;  //complement 
assign odh = ~ODH;  //complement 
assign odp = ~ODP;  //complement 
assign GHD =  EPA & EHB & EHC  |  EPB & EHC  |  EPC  ; 
assign ghd = ~GHD; //complement 
assign DAH = ZZO & ~aah & ~bah  |  QDC & ~aah & bah  |  QDB & aah & ~bah  |  QDA & aah & bah; 
assign dah = ~DAH;  //complement 
assign DAP = ZZO & ~aap & ~bap  |         QDC & ~aap & bap  |  QDB & aap & ~bap  |  QDA & aap & bap ; 
assign dap = ~DAP;  //complement 
assign DBH = ZZO & ~abh & ~bbh  |  QEC & ~abh & bbh  |  QEB & abh & ~bbh  |  QEA & abh & bbh; 
assign dbh = ~DBH;  //complement 
assign DBP = ZZO & ~abp & ~bbp  |         QEC & ~abp & bbp  |  QEB & abp & ~bbp  |  QEA & abp & bbp ; 
assign dbp = ~DBP;  //complement 
assign hmb = ~HMB;  //complement 
assign hmc = ~HMC;  //complement 
assign hmd = ~HMD;  //complement 
assign hnb = ~HNB;  //complement 
assign iaa = ~IAA; //complement 
assign iab = ~IAB; //complement 
assign iac = ~IAC; //complement 
assign iad = ~IAD; //complement 
assign iae = ~IAE; //complement 
assign iaf = ~IAF; //complement 
assign iag = ~IAG; //complement 
assign iah = ~IAH; //complement 
assign iai = ~IAI; //complement 
assign iaj = ~IAJ; //complement 
assign iak = ~IAK; //complement 
assign ial = ~IAL; //complement 
assign iam = ~IAM; //complement 
assign ian = ~IAN; //complement 
assign iao = ~IAO; //complement 
assign iap = ~IAP; //complement 
assign iba = ~IBA; //complement 
assign ibb = ~IBB; //complement 
assign ibc = ~IBC; //complement 
assign ibd = ~IBD; //complement 
assign ibe = ~IBE; //complement 
assign ibf = ~IBF; //complement 
assign ibg = ~IBG; //complement 
assign ibh = ~IBH; //complement 
assign ibi = ~IBI; //complement 
assign ibj = ~IBJ; //complement 
assign ibk = ~IBK; //complement 
assign ibl = ~IBL; //complement 
assign ibm = ~IBM; //complement 
assign ibn = ~IBN; //complement 
assign ibo = ~IBO; //complement 
assign ibp = ~IBP; //complement 
assign ica = ~ICA; //complement 
assign icb = ~ICB; //complement 
assign icc = ~ICC; //complement 
assign icd = ~ICD; //complement 
assign ice = ~ICE; //complement 
assign icf = ~ICF; //complement 
assign icg = ~ICG; //complement 
assign ich = ~ICH; //complement 
assign ici = ~ICI; //complement 
assign icj = ~ICJ; //complement 
assign ick = ~ICK; //complement 
assign icl = ~ICL; //complement 
assign icm = ~ICM; //complement 
assign icn = ~ICN; //complement 
assign ico = ~ICO; //complement 
assign icp = ~ICP; //complement 
assign ida = ~IDA; //complement 
assign idb = ~IDB; //complement 
assign idc = ~IDC; //complement 
assign idd = ~IDD; //complement 
assign ide = ~IDE; //complement 
assign idf = ~IDF; //complement 
assign idg = ~IDG; //complement 
assign idh = ~IDH; //complement 
assign idi = ~IDI; //complement 
assign idj = ~IDJ; //complement 
assign idk = ~IDK; //complement 
assign idl = ~IDL; //complement 
assign idm = ~IDM; //complement 
assign idn = ~IDN; //complement 
assign ido = ~IDO; //complement 
assign idp = ~IDP; //complement 
assign ifa = ~IFA; //complement 
assign ifb = ~IFB; //complement 
assign ifc = ~IFC; //complement 
assign ifd = ~IFD; //complement 
assign ife = ~IFE; //complement 
assign ifff  = ~IFFF ; //complement 
assign ifg = ~IFG; //complement 
assign ifh = ~IFH; //complement 
assign ifi = ~IFI; //complement 
assign ifj = ~IFJ; //complement 
assign ifk = ~IFK; //complement 
assign ifl = ~IFL; //complement 
always@(posedge IZZ )
   begin 
 BAA <=  BAA & TEA  |  IAA & TFA  |  ICA & TGA  |  ACA  ; 
 BAI <=  BAI & TEA  |  IAI & TFA  |  ICI & TGA  |  ACI  ; 
 BBA <=  BBA & TEB  |  IBA & TFB  |  IDA & TGB  |  ADA  ; 
 BBI <=  BBI & TEB  |  IBI & TFB  |  IDI & TGB  |  ADI  ; 
 BCA <= TDA & BAA ; 
 BCB <= TDA & BAB ; 
 BCC <= TDA & BAC ; 
 BCD <= TDA & BAD ; 
 EAA <=  TSA & baa  |  tsa & BAA  |  AAA  ; 
 EAB <=  TSA & bab  |  tsa & BAB  |  AAB  ; 
 EAC <=  TSA & bac  |  tsa & BAC  |  AAC  ; 
 EAD <=  TSA & bad  |  tsa & BAD  |  AAD  ; 
 MAA <=  TLA & KAA  |  TMA & KBP  |  TLC & KBA  |  TNA & LAA  |  NAA  ; 
 MAI <=  TLA & KAI  |  TMA & KBH  |  TLC & KBI  |  TNA & LAI  |  NAI  ; 
 MBA <=  TLB & KBA  |  TMB & KAP  |  TMC & KBP  |  TNB & LBA  |  NBA  ; 
 MBI <=  TLB & KBI  |  TMB & KAH  |  TMC & KBH  |  TNB & LBI  |  NBI  ; 
 QAA <= IFA ; 
 QAB <= IFB ; 
 QAC <= IFC ; 
 QAD <= IFD ; 
 QAE <= IFE ; 
 QAF <= IFFF  ; 
 QAG <= IFG ; 
 QAH <= IFH ; 
 QAI <= IFI ; 
 QAJ <= IFJ ; 
 QAK <= IFK ; 
 QAL <= IFL ; 
 QDA <=  QAE  |  QAG  ; 
 QDB <=  QAF  |  QAG  ; 
 QDC <=  QAF  |  QAG  ; 
 AAA <=  AAA & TAA  |  IAA & TBA  |  ICA & TCA  |  BCA  ; 
 AAI <=  AAI & TAA  |  IAI & TBA  |  ICI & TCA  |  BCI  ; 
 ABA <=  ABA & TAB  |  IBA & TBB  |  IDA & TCB  |  BDA  ; 
 ABI <=  ABI & TAB  |  IBI & TBB  |  IDI & TCB  |  BDI  ; 
 eia <=  TSC & baa  |  tsc & BAA  |  aaa  ; 
 eib <=  TSC & bab  |  tsc & BAB  |  aab  ; 
 eic <=  TSC & bac  |  tsc & BAC  |  aac  ; 
 eid <=  TSC & bad  |  tsc & BAD  |  aad  ; 
 QEA <= QAG; 
 QEB <=  QAF  |  QAG  ; 
 QEC <=  QAF  |  QAG  ; 
 qdd <=  qae & qaf & qag  ; 
 TBA <= QAI ; 
 TBB <= QAI ; 
 TCA <= QAK ; 
 TCB <= QAK ; 
 QFA <= IAA ; 
 QFB <= IAB ; 
 QFC <= IAC ; 
 QFD <= IAD ; 
 QBA <= QAA ; 
 QBB <= QAB ; 
 QBC <= QAC ; 
 QBD <= QAD ; 
 QBH <= QAH ; 
 TFA <= QAJ ; 
 TFB <= QAJ ; 
 TGA <= QAL ; 
 TGB <= QAL ; 
 KAA <=  JAA & TQA  |  JAE & TQB  |  JAI & TQC  |  JAM & TQD  ; 
 KAI <=  JAI & TQA  |  JAM & TQB  |  JBA & TQC  |  JBE & TQD  ; 
 KBA <=  JBA & TQE  |  JBE & TQF  |  JBI & TQG  |  JBM & TQH  ; 
 KBI <=  JBI & TQE  |  JBM & TQF  ; 
 TPE <= iab & iaa ; 
 TPF <= iab & IAA ; 
 TPG <= IAB & iaa ; 
 TPH <= IAB & IAA ; 
 OAA <= AAA & TRA |  BAA & tra ; 
 OAI <= AAI & TRA |  BAI & tra ; 
 OEC <= BBP ; 
 QAP <=  IFA  |  IFB  |  IFC  |  IFD  ; 
 QBI <= QAI ; 
 QBJ <= QAJ ; 
 QBK <= QAK ; 
 QBL <= QAL ; 
 OBA <= ABA & TRB |  BBA & trb ; 
 OBI <= ABI & TRB |  BBI & trb ; 
 QAQ <=  IFE  |  IFFF   |  IFG  |  IFH  ; 
 oea <=  jca  |  jcb  |  jcc  |  jcd  ; 
 oeb <=  jda  |  jdb  |  jdc  |  jdd  ; 
 OCA <= AAA & TTA |  BAA & tta ; 
 OCI <= AAI & TTA |  BAI & tta ; 
 TIA <= QDD ; 
 TIB <= QDD ; 
 TJA <= QAH ; 
 TJB <= QAH ; 
 TNA <=  QAA  |  QAB  ; 
 TNB <=  QAA  |  QAB  ; 
 TSA <= QAA ; 
 TSB <= QAA ; 
 TSC <= QAA ; 
 TSD <= QAA ; 
 ODA <= ABA & TTB |  BBA & ttb ; 
 ODI <= ABI & TTB |  BBI & ttb ; 
 taa <=  QAI  |  QAK  |  QAH  ; 
 QGE <= QFE ; 
 KKA <=  HAH & HAK  |  HAI & HAK  |  HAJ  ; 
 tab <=  QAI  |  QAK  |  QAH  ; 
 TOA <= QDD ; 
 TOB <= QDD ; 
 HAK <= GNA ; 
 TLA <= QBC & qfe ; 
 TLB <= QBC & qfe ; 
 TLC <= QBC & QFE ; 
 LAA <= HBA & qbb |  HJA & QBB ; 
 LAB <= HBB & qbb |  HJB & QBB ; 
 LAC <= HBC & qbb |  HJC & QBB ; 
 LBA <= HFA & had |  HNA & HAD ; 
 LBB <= HFB & had |  HNB & HAD ; 
 LBC <= HFC & had |  HNC & HAD ; 
 TPA <= iab & iaa ; 
 TPB <= iab & IAA ; 
 TPC <= IAB & iaa ; 
 TPD <= IAB & IAA ; 
 EBA <=  TSA & bae  |  tsa & BAE  |  AAE  ; 
 EBB <=  TSA & baf  |  tsa & BAF  |  AAF  ; 
 EBC <=  TSA & bag  |  tsa & BAG  |  AAG  ; 
 TRA <= QAJ ; 
 TRB <= QAJ ; 
 EBD <=  TSA & bah  |  tsa & BAH  |  AAH  ; 
 MAB <=  TLA & KAB  |  TMA & KBO  |  TLC & KBB  |  TNA & LAB  |  NAB  ; 
 MAJ <=  TLA & KAJ  |  TMA & KBG  |  TLC & KBJ  |  TNA & LAJ  |  NAJ  ; 
 MBB <=  TLB & KBB  |  TMB & KAO  |  TMC & KBO  |  TNB & LBB  |  NBB  ; 
 MBJ <=  TLB & KBJ  |  TMB & KAG  |  TMC & KBG  |  TNB & LBJ  |  NBJ  ; 
 TDA <= QAH ; 
 TDB <= QAH ; 
 HAC <=  GAE & GIA & GJA  |  GBE & GJA  |  GCE  ; 
 HAD <=  GAE & GIA & GJA & GKA  |  GBE & GJA & GKA  |  GCE & GKA  |  GDE  ; 
 TMA <= QBD & qfe ; 
 TMB <= QBD & qfe ; 
 TMC <= QBD & QFE ; 
 AAB <=  AAB & TAA  |  IAB & TBA  |  ICB & TCA  |  BCB  ; 
 AAJ <=  AAJ & TAA  |  IAJ & TBA  |  ICJ & TCA  |  BCJ  ; 
 ABB <=  ABB & TAB  |  IBB & TBB  |  IDB & TCB  |  BDB  ; 
 ABJ <=  ABJ & TAB  |  IBJ & TBB  |  IDJ & TCB  |  BDJ  ; 
 BAB <=  BAB & TEA  |  IAB & TFA  |  ICB & TGA  |  ACB  ; 
 BAJ <=  BAJ & TEA  |  IAJ & TFA  |  ICJ & TGA  |  ACJ  ; 
 BBB <=  BBB & TEB  |  IBB & TFB  |  IDB & TGB  |  ADB  ; 
 BBJ <=  BBJ & TEB  |  IBJ & TFB  |  IDJ & TGB  |  ADJ  ; 
 eja <=  TSC & bae  |  tsc & BAE  |  aae  ; 
 ejb <=  TSC & baf  |  tsc & BAF  |  aaf  ; 
 ejc <=  TSC & bag  |  tsc & BAG  |  aag  ; 
 ejd <=  TSC & bah  |  tsc & BAH  |  aah  ; 
 tea <=  QAJ  |  QAL  |  QAP  |  QAQ  ; 
 teb <=  QAJ  |  QAL  |  QAP  |  QAQ  ; 
 HAE <=  GAE & GIA & GJA & GKA & GLA  |  GBE & GJA & GKA & GLA  |  GCE & GKA & GLA  |  ZZI & GDE & GLA  |  GEE  ; 
 haf <=  gae  |  gia  |  gja  |  gpa  |  gqa  ; 
 KAB <=  JAB & TQA  |  JAF & TQB  |  JAJ & TQC  |  JAN & TQD  ; 
 KAJ <=  JAJ & TQA  |  JAN & TQB  |  JBB & TQC  |  JBF & TQD  ; 
 KBB <=  JBB & TQE  |  JBF & TQF  |  JBJ & TQG  |  JBN & TQH  ; 
 KBJ <=  JBJ & TQE  |  JBN & TQF  ; 
 TQC <= QFD & qfc ; 
 TQD <= QFD & QFC ; 
 TQE <= qfd & qfc ; 
 TQF <= qfd & QFC ; 
 TQH <= QFD & QFC ; 
 TQG <= QFD & qfc ; 
 OAB <= AAB & TRA |  BAB & tra ; 
 OAJ <= AAJ & TRA |  BAJ & tra ; 
 LBD <= HFD & had |  HND & HAD ; 
 HAA <= GAE ; 
 HBA <= EAA ; 
 HCA <= EBA ; 
 HDA <= ECA ; 
 HAB <=  GAE & GIA  |  GBE  ; 
 OBB <= ABB & TRB |  BBB & trb ; 
 OBJ <= ABJ & TRB |  BBJ & trb ; 
 HEA <= EDA ; 
 HFA <= EEA ; 
 HGA <= EFA ; 
 HHA <= EGA ; 
 HBB <= EAB & gab |  eab & GAB ; 
 HBC <= EAC & gac |  eac & GAC ; 
 OCB <= AAB & TTA |  BAB & tta ; 
 OCJ <= AAJ & TTA |  BAJ & tta ; 
 HBD <= EAD & gad |  ead & GAD ; 
 HCB <= EBB & gbb |  ebb & GBB ; 
 HCC <= EBC & gbc |  ebc & GBC ; 
 ODB <= ABB & TTB |  BBB & ttb ; 
 ODJ <= ABJ & TTB |  BBJ & ttb ; 
 HCD <= EBD & gbd |  ebd & GBD ; 
 HHB <= EGB & ggb |  egb & GGB ; 
 HHC <= EGC & ggc |  egc & GGC ; 
 HHD <= EGD & ggd |  egd & GGD ; 
 HAG <=  GBE & GJA & GKA & GLA & GMA  |  GCE & GKA & GLA & GMA  |  GDE & GLA & GMA  |  ZZI & GEE & GMA  |  GFE  ; 
 LAE <= HCA & haa |  HKA & HAA ; 
 LAF <= HCB & haa |  HKB & HAA ; 
 LBE <= HGA & hae |  HOA & HAE ; 
 LBF <= HGB & hae |  HOB & HAE ; 
 TQA <= qfd & qfc ; 
 TQB <= qfd & QFC ; 
 BBC <=  BBC & TEB  |  IBC & TFB  |  IDC & TGB  |  ADC  ; 
 BBK <=  BBK & TEB  |  IBK & TFB  |  IDK & TGB  |  ADK  ; 
 ECA <=  TSA & bai  |  tsa & BAI  |  AAI  ; 
 BDA <= TDB & BBA ; 
 BDB <= TDB & BBB ; 
 BDC <= TDB & BBC ; 
 BDD <= TDB & BBD ; 
 ECB <=  TSA & baj  |  tsa & BAJ  |  AAJ  ; 
 ECC <=  TSA & bak  |  tsa & BAK  |  AAK  ; 
 ECD <=  TSA & bal  |  tsa & BAL  |  AAL  ; 
 MAC <=  TLA & KAC  |  TMA & KBN  |  TLC & KBC  |  TNA & LAC  |  NAC  ; 
 MAK <=  TLA & KAK  |  TMA & KBF  |  TLC & KBK  |  TNA & LAK  |  NAK  ; 
 MBC <=  TLB & KBC  |  TMB & KAN  |  TMC & KBN  |  TNB & LBC  |  NBC  ; 
 MBK <=  TLB & KBK  |  TMB & KAF  |  TMC & KBF  |  TNB & LBK  |  NBK  ; 
 AAC <=  AAC & TAA  |  IAC & TBA  |  ICC & TCA  |  BCC  ; 
 AAK <=  AAK & TAA  |  IAK & TBA  |  ICK & TCA  |  BCK  ; 
 ABC <=  ABC & TAB  |  IBC & TBB  |  IDC & TCB  |  BDC  ; 
 ABK <=  ABK & TAB  |  IBK & TBB  |  IDK & TCB  |  BDK  ; 
 BAC <=  BAC & TEA  |  IAC & TFA  |  ICC & TGA  |  ACC  ; 
 BAK <=  BAK & TEA  |  IAK & TFA  |  ICK & TGA  |  ACK  ; 
 eka <=  TSC & bai  |  tsc & BAI  |  aai  ; 
 ekb <=  TSC & baj  |  tsc & BAJ  |  aaj  ; 
 ekc <=  TSC & bak  |  tsc & BAK  |  aak  ; 
 ekd <=  TSC & bal  |  tsc & BAL  |  aal  ; 
 TTA <= QAI ; 
 TTB <= QAI ; 
 HIA <= EHA ; 
 HJA <= eaa ; 
 HKA <= eba ; 
 HLA <= eca ; 
 HMA <= eda ; 
 HNA <= eea ; 
 HOA <= efa ; 
 HPA <= ega ; 
 HQA <= eha ; 
 HQB <= EHB & ghf |  ehb & GHF ; 
 HQC <= EHC & ghg |  ehc & GHG ; 
 HQD <= EHD & ghh |  ehd & GHH ; 
 KAC <=  JAC & TQA  |  JAG & TQB  |  JAK & TQC  |  JAO & TQD  ; 
 KAK <=  JAK & TQA  |  JAO & TQB  |  JBC & TQC  |  JBG & TQD  ; 
 KBC <=  JBC & TQE  |  JBG & TQF  |  JBK & TQG  |  JBO & TQH  ; 
 KBK <=  JBK & TQE  |  JBO & TQF  ; 
 LBJ <=  HHB & haf & hag  |  HPB & HAF  |  HPB & HAG  ; 
 LAJ <= HDB & hab |  HLB & HAB ; 
 LAK <= HDC & hab |  HLC & HAB ; 
 LAL <= HDD & hab |  HLD & HAB ; 
 hah <=  gae  |  gia  |  gja  |  gpa  |  gqa  ; 
 OAC <= AAC & TRA |  BAC & tra ; 
 OAK <= AAK & TRA |  BAK & tra ; 
 LAI <= HDA & hab |  HLA & HAB ; 
 LBK <=  HHC & haf & hag  |  HPC & HAF  |  HPC & HAG  ; 
 LBL <=  HHD & haf & hag  |  HPD & HAF  |  HPD & HAG  ; 
 OBC <= ABC & TRB |  BBC & trb ; 
 OBK <= ABK & TRB |  BBK & trb ; 
 HDB <= ECB & gcb |  ecb & GCB ; 
 HDC <= ECC & gcc |  ecc & GCC ; 
 HDD <= ECD & gcd |  ecd & GCD ; 
 OCC <= AAC & TTA |  BAC & tta ; 
 OCK <= AAK & TTA |  BAK & tta ; 
 hai <=  gbe  |  gja  |  gka  |  gla  |  gma  ; 
 HAJ <=  GCE & GKA & GLA & GMA & GNA  |  GDE & GLA & GMA & GNA  |  GEE & GMA & GNA  |  ZZI & GFE & GNA  |  GGE  ; 
 ODC <= ABC & TTB |  BBC & ttb ; 
 ODK <= ABK & TTB |  BBK & ttb ; 
 LAG <= HCC & haa |  HKC & HAA ; 
 LAH <= HCD & haa |  HKD & HAA ; 
 LBG <= HGC & hae |  HOC & HAE ; 
 LBH <= HGD & hae |  HOD & HAE ; 
 LBI <=  HHA & haf & hag  |  HPA & HAF  |  HPA & HAG  ; 
 EDA <=  TSA & bam  |  tsa & BAM  |  AAM  ; 
 EDB <=  TSA & ban  |  tsa & BAN  |  AAN  ; 
 EDC <=  TSA & bao  |  tsa & BAO  |  AAO  ; 
 BDE <= TDB & BBE ; 
 BDF <= TDB & BBF ; 
 BDG <= TDB & BBG ; 
 BDH <= TDB & BBH ; 
 EDD <=  TSA & bap  |  tsa & BAP  |  AAP  ; 
 MAD <=  TLA & KAD  |  TMA & KBM  |  TLC & KBD  |  TNA & LAD  |  NAD  ; 
 MAL <=  TLA & KAL  |  TMA & KBE  |  TLC & KBL  |  TNA & LAL  |  NAL  ; 
 MBD <=  TLB & KBD  |  TMB & KAM  |  TMC & KBM  |  TNB & LBD  |  NBD  ; 
 MBL <=  TLB & KBL  |  TMB & KAE  |  TMC & KBE  |  TNB & LBL  |  NBL  ; 
 AAD <=  AAD & TAA  |  IAD & TBA  |  ICD & TCA  |  BCD  ; 
 AAL <=  AAL & TAA  |  IAL & TBA  |  ICL & TCA  |  BCL  ; 
 ABD <=  ABD & TAB  |  IBD & TBB  |  IDD & TCB  |  BDD  ; 
 ABL <=  ABL & TAB  |  IBL & TBB  |  IDL & TCB  |  BDL  ; 
 BAD <=  BAD & TEA  |  IAD & TFA  |  ICD & TGA  |  ACD  ; 
 BAL <=  BAL & TEA  |  IAL & TFA  |  ICL & TGA  |  ACL  ; 
 BBD <=  BBD & TEB  |  IBD & TFB  |  IDD & TGB  |  ADD  ; 
 BBL <=  BBL & TEB  |  IBL & TFB  |  IDL & TGB  |  ADL  ; 
 ela <=  TSC & bam  |  tsc & BAM  |  aam  ; 
 elb <=  TSC & ban  |  tsc & BAN  |  aan  ; 
 elc <=  TSC & bao  |  tsc & BAO  |  aao  ; 
 eld <=  TSC & bap  |  tsc & BAP  |  aap  ; 
 KAD <=  JAD & TQA  |  JAH & TQB  |  JAL & TQC  |  JAP & TQD  ; 
 KAL <=  JAL & TQA  |  JAP & TQB  |  JBD & TQC  |  JBH & TQD  ; 
 KBD <=  JBD & TQE  |  JBH & TQF  |  JBL & TQG  |  JBP & TQH  ; 
 KBL <=  JBL & TQE  |  JBP & TQF  ; 
 OAD <= AAD & TRA |  BAD & tra ; 
 OAL <= AAL & TRA |  BAL & tra ; 
 OBD <= ABD & TRB |  BBD & trb ; 
 OBL <= ABL & TRB |  BBL & trb ; 
 OCD <= AAD & TTA |  BAD & tta ; 
 OCL <= AAL & TTA |  BAL & tta ; 
 ODD <= ABD & TTB |  BBD & ttb ; 
 ODL <= ABL & TTB |  BBL & ttb ; 
 HEB <= EDB & gdb |  edb & GDB ; 
 HEC <= EDC & gdc |  edc & GDC ; 
 HED <= EDD & gdd |  edd & GDD ; 
 EEA <=  TSB & bba  |  tsb & BBA  |  ABA  ; 
 EEB <=  TSB & bbb  |  tsb & BBB  |  ABB  ; 
 EEC <=  TSB & bbc  |  tsb & BBC  |  ABC  ; 
 BCE <= TDA & BAE ; 
 BCF <= TDA & BAF ; 
 BCG <= TDA & BAG ; 
 BCH <= TDA & BAH ; 
 EED <=  TSB & bbd  |  tsb & BBD  |  ABD  ; 
 MAE <=  TLA & KAE  |  TMA & KBL  |  TLC & KBE  |  TNA & LAE  |  NAE  ; 
 MAM <=  TLA & KAM  |  TMA & KBD  |  TLC & KBM  |  TNA & LAM  |  NAM  ; 
 MBE <=  TLB & KBE  |  TMB & KAL  |  TMC & KBL  |  TNB & LBE  |  NBE  ; 
 MBM <=  TLB & KBM  |  TMB & KAD  |  TMC & KBD  |  TNB & LBM  |  NBM  ; 
 AAE <=  AAE & TAA  |  IAE & TBA  |  ICE & TCA  |  BCE  ; 
 AAM <=  AAM & TAA  |  IAM & TBA  |  ICM & TCA  |  BCM  ; 
 ABE <=  ABE & TAB  |  IBE & TBB  |  IDE & TCB  |  BDE  ; 
 ABM <=  ABM & TAB  |  IBM & TBB  |  IDM & TCB  |  BDM  ; 
 BAE <=  BAE & TEA  |  IAE & TFA  |  ICE & TGA  |  ACE  ; 
 BAM <=  BAM & TEA  |  IAM & TFA  |  ICM & TGA  |  ACM  ; 
 BBE <=  BBE & TEB  |  IBE & TFB  |  IDE & TGB  |  ADE  ; 
 BBM <=  BBM & TEB  |  IBM & TFB  |  IDM & TGB  |  ADM  ; 
 ema <=  TSD & bba  |  tsd & BBA  |  aba  ; 
 emb <=  TSD & bbb  |  tsd & BBB  |  abb  ; 
 emc <=  TSD & bbc  |  tsd & BBC  |  abc  ; 
 emd <=  TSD & bbd  |  tsd & BBD  |  abd  ; 
 HFB <= EEB & geb |  eeb & GEB ; 
 HFC <= EEC & gec |  eec & GEC ; 
 HFD <= EED & ged |  eed & GED ; 
 KAE <=  JAE & TQA  |  JAI & TQB  |  JAM & TQC  |  JBA & TQD  ; 
 KAM <=  JAM & TQA  |  JBA & TQB  |  JBE & TQC  |  JBI & TQD  ; 
 KBE <=  JBE & TQE  |  JBI & TQF  |  JBM & TQG  ; 
 KBM <=  JBM & TQE  ; 
 OAE <= AAE & TRA |  BAE & tra ; 
 OAM <= AAM & TRA |  BAM & tra ; 
 OBE <= ABE & TRB |  BBE & trb ; 
 OBM <= ABM & TRB |  BBM & trb ; 
 OCE <= AAE & TTA |  BAE & tta ; 
 OCM <= AAM & TTA |  BAM & tta ; 
 ODE <= ABE & TTB |  BBE & ttb ; 
 ODM <= ABM & TTB |  BBM & ttb ; 
 LAM <= HEA & hac |  HMA & HAC ; 
 LAN <= HEB & hac |  HMB & HAC ; 
 LAO <= HEC & hac |  HMC & HAC ; 
 LBM <= HIA & kka |  HQA & KKA ; 
 LBN <= HIB & kka |  HQB & KKA ; 
 LBO <= HIC & kka |  HQC & KKA ; 
 LAP <= HED & hac |  HMD & HAC ; 
 LBP <= HID & kka |  HQD & KKA ; 
 EFA <=  TSB & bbe  |  tsb & BBE  |  ABE  ; 
 EFB <=  TSB & bbf  |  tsb & BBF  |  ABF  ; 
 EFC <=  TSB & bbg  |  tsb & BBG  |  ABG  ; 
 BCI <= TDA & BAI ; 
 BCJ <= TDA & BAJ ; 
 BCK <= TDA & BAK ; 
 BCL <= TDA & BAL ; 
 EFD <=  TSB & bbh  |  tsb & BBH  |  ABH  ; 
 MAF <=  TLA & KAF  |  TMA & KBK  |  TLC & KBF  |  TNA & LAF  |  NAF  ; 
 MAN <=  TLA & KAN  |  TMA & KBC  |  TLC & KBN  |  TNA & LAN  |  NAN  ; 
 MBF <=  TLB & KBF  |  TMB & KAK  |  TMC & KBK  |  TNB & LBF  |  NBF  ; 
 MBN <=  TLB & KBN  |  TMB & KAC  |  TMC & KBC  |  TNB & LBN  |  NBN  ; 
 AAF <=  AAF & TAA  |  IAF & TBA  |  ICF & TCA  |  BCF  ; 
 AAN <=  AAN & TAA  |  IAN & TBA  |  ICN & TCA  |  BCN  ; 
 ABF <=  ABF & TAB  |  IBF & TBB  |  IDF & TCB  |  BDF  ; 
 ABN <=  ABN & TAB  |  IBN & TBB  |  IDN & TCB  |  BDN  ; 
 BAF <=  BAF & TEA  |  IAF & TFA  |  ICF & TGA  |  ACF  ; 
 BAN <=  BAN & TEA  |  IAN & TFA  |  ICN & TGA  |  ACN  ; 
 BBF <=  BBF & TEB  |  IBF & TFB  |  IDF & TGB  |  ADF  ; 
 BBN <=  BBN & TEB  |  IBN & TFB  |  IDN & TGB  |  ADN  ; 
 ena <=  TSD & bbe  |  tsd & BBE  |  abe  ; 
 enb <=  TSD & bbf  |  tsd & BBF  |  abf  ; 
 enc <=  TSD & bbg  |  tsd & BBG  |  abg  ; 
 endd <=  TSD & bbh  |  tsd & BBH  |  abh  ; 
 HIB <= EHB & ghb |  ehb & GHB ; 
 HIC <= EHC & ghc |  ehc & GHC ; 
 HID <= EHD & ghd |  ehd & GHD ; 
 HJB <= EAB & gaf |  eab & GAF ; 
 HJC <= EAC & gag |  eac & GAG ; 
 HJD <= EAD & gah |  ead & GAH ; 
 HKB <= EBB & gbf |  ebb & GBF ; 
 HKC <= EBC & gbg |  ebc & GBG ; 
 HKD <= EBD & gbh |  ebd & GBH ; 
 HLB <= ECB & gcf |  ecb & GCF ; 
 HLC <= ECC & gcg |  ecc & GCG ; 
 HLD <= ECD & gch |  ecd & GCH ; 
 KAF <=  JAF & TQA  |  JAJ & TQB  |  JAN & TQC  |  JBB & TQD  ; 
 KAN <=  JAN & TQA  |  JBB & TQB  |  JBF & TQC  |  JBJ & TQD  ; 
 KBF <=  JBF & TQE  |  JBJ & TQF  |  JBN & TQG  ; 
 KBN <=  JBN & TQE  ; 
 OAF <= AAF & TRA |  BAF & tra ; 
 OAN <= AAN & TRA |  BAN & tra ; 
 OBF <= ABF & TRB |  BBF & trb ; 
 OBN <= ABN & TRB |  BBN & trb ; 
 OCF <= AAF & TTA |  BAF & tta ; 
 OCN <= AAN & TTA |  BAN & tta ; 
 ODF <= ABF & TTB |  BBF & ttb ; 
 ODN <= ABN & TTB |  BBN & ttb ; 
 HGB <= EFB & gfb |  efb & GFB ; 
 HGC <= EFC & gfc |  efc & GFC ; 
 HGD <= EFD & gfd |  efd & GFD ; 
 EGA <=  TSB & bbi  |  tsb & BBI  |  ABI  ; 
 EGB <=  TSB & bbj  |  tsb & BBJ  |  ABJ  ; 
 EGC <=  TSB & bbk  |  tsb & BBK  |  ABK  ; 
 BCM <= TDA & BAM ; 
 BCN <= TDA & BAN ; 
 BCO <= TDA & BAO ; 
 BCP <= TDA & BAP ; 
 EGD <=  TSB & bbl  |  tsb & BBL  |  ABL  ; 
 MAG <=  TLA & KAG  |  TMA & KBJ  |  TLC & KBG  |  TNA & LAG  |  NAG  ; 
 MAO <=  TLA & KAO  |  TMA & KBB  |  TLC & KBO  |  TNA & LAO  |  NAO  ; 
 MBG <=  TLB & KBG  |  TMB & KAJ  |  TMC & KBJ  |  TNB & LBG  |  NBG  ; 
 MBO <=  TLB & KBO  |  TMB & KAB  |  TMC & KBB  |  TNB & LBO  |  NBO  ; 
 AAG <=  AAG & TAA  |  IAG & TBA  |  ICG & TCA  |  BCG  ; 
 AAO <=  AAO & TAA  |  IAO & TBA  |  ICO & TCA  |  BCO  ; 
 ABG <=  ABG & TAB  |  IBG & TBB  |  IDG & TCB  |  BDG  ; 
 ABO <=  ABO & TAB  |  IBO & TBB  |  IDO & TCB  |  BDO  ; 
 BAG <=  BAG & TEA  |  IAH & TFA  |  ICG & TGA  |  ACG  ; 
 BAO <=  BAO & TEA  |  IAO & TFA  |  ICO & TGA  |  ACO  ; 
 BBG <=  BBG & TEB  |  IBH & TFB  |  IDG & TGB  |  ADG  ; 
 BBO <=  BBO & TEB  |  IBO & TFB  |  IDO & TGB  |  ADO  ; 
 eoa <=  TSD & bbi  |  tsd & BBI  |  abi  ; 
 eob <=  TSD & bbj  |  tsd & BBJ  |  abj  ; 
 eoc <=  TSD & bbk  |  tsd & BBK  |  abk  ; 
 eod <=  TSD & bbl  |  tsd & BBL  |  abl  ; 
 KAG <=  JAG & TQA  |  JAK & TQB  |  JAO & TQC  |  JBC & TQD  ; 
 KAO <=  JAO & TQA  |  JBC & TQB  |  JBG & TQC  |  JBK & TQD  ; 
 KBG <=  JBG & TQE  |  JBK & TQF  |  JBO & TQG  ; 
 KBO <=  JBO & TQE  ; 
 OAG <= AAG & TRA |  BAG & tra ; 
 OAO <= AAO & TRA |  BAO & tra ; 
 OBG <= ABG & TRB |  BBG & trb ; 
 OBO <= ABO & TRB |  BBO & trb ; 
 OCG <= AAG & TTA |  BAG & tta ; 
 OCO <= AAO & TTA |  BAO & tta ; 
 ODG <= ABG & TTB |  BBG & ttb ; 
 ODO <= ABO & TTB |  BBO & ttb ; 
 EHA <=  TSB & bbm  |  tsb & BBM  |  ABM  ; 
 EHB <=  TSB & bbn  |  tsb & BBN  |  ABN  ; 
 EHC <=  TSB & bbo  |  tsb & BBO  |  ABO  ; 
 BDI <= TDB & BBI ; 
 BDJ <= TDB & BBJ ; 
 BDK <= TDB & BBK ; 
 BDL <= TDB & BBL ; 
 EHD <=  TSB & bbp  |  tsb & BBP  |  ABP  ; 
 MAH <=  TLA & KAH  |  TMA & KBI  |  TLC & KBH  |  TNA & LAH  |  NAH  ; 
 MAP <=  TLA & KAP  |  TMA & KBA  |  TLC & KBP  |  TNA & LAP  |  NAP  ; 
 MBH <=  TLB & KBH  |  TMB & KAI  |  TMC & KBI  |  TNB & LBH  |  NBH  ; 
 MBP <=  TLB & KBP  |  TMB & KAA  |  TMC & KBA  |  TNB & LBP  |  NBP  ; 
 BDM <= TDB & BBM ; 
 BDN <= TDB & BBN ; 
 BDO <= TDB & BBO ; 
 BDP <= TDB & BBP ; 
 AAH <=  AAH & TAA  |  IAH & TBA  |  ICH & TCA  |  BCH  ; 
 AAP <=  AAP & TAA  |  IAP & TBA  |  ICP & TCA  |  BCP  ; 
 ABH <=  ABH & TAB  |  IBH & TBB  |  IDH & TCB  |  BDH  ; 
 ABP <=  ABP & TAB  |  IBP & TBB  |  IDP & TCB  |  BDP  ; 
 BAH <=  BAH & TEA  |  IAH & TFA  |  ICH & TGA  |  ACH  ; 
 BAP <=  BAP & TEA  |  IAP & TFA  |  ICP & TGA  |  ACP  ; 
 BBH <=  BBH & TEB  |  IBH & TFB  |  IDH & TGB  |  ADH  ; 
 BBP <=  BBP & TEB  |  IBP & TFB  |  IDP & TGB  |  ADP  ; 
 epa <=  TSD & bbm  |  tsd & BBM  |  abm  ; 
 epb <=  TSD & bbn  |  tsd & BBN  |  abn  ; 
 epc <=  TSD & bbo  |  tsd & BBO  |  abo  ; 
 epd <=  TSD & bbp  |  tsd & BBP  |  abp  ; 
 KAH <=  JAH & TQA  |  JAL & TQB  |  JAP & TQC  |  JBD & TQD  ; 
 KAP <=  JAP & TQA  |  JBD & TQB  |  JBH & TQC  |  JBL & TQD  ; 
 KBH <=  JBH & TQE  |  JBL & TQF  |  JBP & TQG  ; 
 KBP <=  JBP & TQE  ; 
 HNC <= EEC & geg |  eec & GEG ; 
 HND <= EED & geh |  eed & GEH ; 
 HOB <= EFB & gff |  efb & GFF ; 
 OAH <= AAH & TRA |  BAH & tra ; 
 OAP <= AAP & TRA |  BAP & tra ; 
 HOC <= EFC & gfg |  efc & GFG ; 
 HOD <= EFD & gfh |  efd & GFH ; 
 HPB <= EGB & ggf |  egb & GGF ; 
 OBH <= ABH & TRB |  BBH & trb ; 
 OBP <= ABP & TRB |  BBP & trb ; 
 HPC <= EGC & ggg |  egc & GGG ; 
 HPD <= EGD & ggh |  egd & GGH ; 
 OCH <= AAH & TTA |  BAH & tta ; 
 OCP <= AAP & TTA |  BAP & tta ; 
 ODH <= ABH & TTB |  BBH & ttb ; 
 ODP <= ABP & TTB |  BBP & ttb ; 
 HMB <= EDB & gdf |  edb & GDF ; 
 HMC <= EDC & gdg |  edc & GDG ; 
 HMD <= EDD & gdh |  edd & GDH ; 
 HNB <= EEB & gef |  eeb & GEF ; 
end
endmodule;
