module kb( IZZ,
 IAA, 
 IAB, 
 IAC, 
 IAD, 
 IAE, 
 IAF, 
 IAG, 
 IAH, 
 IAI, 
 IAJ, 
 IAK, 
 IAL, 
 IAM, 
 IAN, 
 IAO, 
 IAP, 
 IAQ, 
 IAS, 
 IAT, 
 IBA, 
 IBB, 
 IBC, 
 IBD, 
 IBE, 
 IBF, 
 IBG, 
 IBH, 
 IBI, 
 IBJ, 
 IBK, 
 IBL, 
 IBM, 
 IBN, 
 IBO, 
 IBP, 
 IBQ, 
 IBS, 
 IBT, 
 ICA, 
 ICB, 
 ICC, 
 ICD, 
 ICE, 
 ICF, 
 ICG, 
 ICH, 
 ICI, 
 ICJ, 
 ICK, 
 ICL, 
 ICM, 
 ICN, 
 ICO, 
 ICP, 
 ICQ, 
 ICS, 
 ICT, 
 IDA, 
 IDB, 
 IDC, 
 IDD, 
 IDE, 
 IDF, 
 IDG, 
 IDH, 
 IDI, 
 IDJ, 
 IDK, 
 IDL, 
 IDM, 
 IDN, 
 IDO, 
 IDP, 
 IDQ, 
 IDS, 
 IDT, 
 IEA, 
 IEB, 
 IEC, 
 IED, 
 IEE, 
 IEF, 
 IEG, 
 IEH, 
 IEI, 
 IEJ, 
 IEK, 
 IEL, 
 IEM, 
 IEN, 
 IEO, 
 IEP, 
 IFA, 
 IFB, 
 IFC, 
 IFD, 
 IFE, 
 IFFF , 
 IFG, 
 IFH, 
 IFI, 
 IFJ, 
 IFK, 
 IFL, 
 IFM, 
 IFN, 
 IFO, 
 IFP, 
 IGA, 
 IGB, 
 IGC, 
 IGD, 
 IGE, 
 IGF, 
 IGG, 
 IGH, 
 IGI, 
 IGJ, 
 IGK, 
 IGL, 
 IHA, 
 IHB, 
 IHC, 
 IHD, 
 IHE, 
 IHF, 
 IHG, 
 IHH, 
 IHI, 
 IHJ, 
 IHK, 
 IHL, 
 OAA, 
 OAB, 
 OAC, 
 OAD, 
 OAE, 
 OAF, 
 OAG, 
 OAH, 
 OAI, 
 OAJ, 
 OAK, 
 OAL, 
 OAM, 
 OAN, 
 OAO, 
 OAP, 
 OAQ, 
 OAR, 
 OAS, 
 OAT, 
 OBA, 
 OBB, 
 OBC, 
 OBD, 
 OBE, 
 OBF, 
 OBG, 
 OBH, 
 OBI, 
 OBJ, 
 OBK, 
 OBL, 
 OBM, 
 OBN, 
 OBO, 
 OBP, 
 OBQ, 
 OBR, 
 OBS, 
 OBT, 
 OCA, 
 OCB, 
 OCC, 
 OCD, 
 OCE, 
 OCF, 
 OCG, 
 OCH, 
 OCI, 
 OCJ, 
 OCK, 
 OCL, 
 OCM, 
 OCN, 
 OCO, 
 OCP, 
 OCQ, 
 OCR, 
 OCS, 
 OCT, 
 ODA, 
 ODB, 
 ODC, 
 ODD, 
 ODE, 
 ODF, 
 ODG, 
 ODH, 
 ODI, 
 ODJ, 
 ODK, 
 ODL, 
 ODM, 
 ODN, 
 ODO, 
 ODP, 
 ODQ, 
 ODR, 
 ODS, 
 ODT, 
 OEA, 
 OEB, 
 OEC, 
 OED, 
 OEE, 
 OEF, 
 OEG, 
 OEH, 
 OEI, 
 OEJ, 
 OEK, 
 OEL, 
 OEM, 
 OEN, 
 OEO, 
 OEP, 
 OFA, 
 OFB, 
 OFC, 
 OFD, 
 OFE, 
 OFF, 
 OFG, 
 OFH, 
 OFI, 
 OFJ, 
 OFK, 
 OFL, 
 OFM, 
 OFN, 
 OFO, 
 OFP, 
 OGA, 
 OGB, 
 OGC, 
 OGD, 
OHA ); 
    
 input IZZ; 
 input IAA; 
 input IAB; 
 input IAC; 
 input IAD; 
 input IAE; 
 input IAF; 
 input IAG; 
 input IAH; 
 input IAI; 
 input IAJ; 
 input IAK; 
 input IAL; 
 input IAM; 
 input IAN; 
 input IAO; 
 input IAP; 
 input IAQ; 
 input IAS; 
 input IAT; 
 input IBA; 
 input IBB; 
 input IBC; 
 input IBD; 
 input IBE; 
 input IBF; 
 input IBG; 
 input IBH; 
 input IBI; 
 input IBJ; 
 input IBK; 
 input IBL; 
 input IBM; 
 input IBN; 
 input IBO; 
 input IBP; 
 input IBQ; 
 input IBS; 
 input IBT; 
 input ICA; 
 input ICB; 
 input ICC; 
 input ICD; 
 input ICE; 
 input ICF; 
 input ICG; 
 input ICH; 
 input ICI; 
 input ICJ; 
 input ICK; 
 input ICL; 
 input ICM; 
 input ICN; 
 input ICO; 
 input ICP; 
 input ICQ; 
 input ICS; 
 input ICT; 
 input IDA; 
 input IDB; 
 input IDC; 
 input IDD; 
 input IDE; 
 input IDF; 
 input IDG; 
 input IDH; 
 input IDI; 
 input IDJ; 
 input IDK; 
 input IDL; 
 input IDM; 
 input IDN; 
 input IDO; 
 input IDP; 
 input IDQ; 
 input IDS; 
 input IDT; 
 input IEA; 
 input IEB; 
 input IEC; 
 input IED; 
 input IEE; 
 input IEF; 
 input IEG; 
 input IEH; 
 input IEI; 
 input IEJ; 
 input IEK; 
 input IEL; 
 input IEM; 
 input IEN; 
 input IEO; 
 input IEP; 
 input IFA; 
 input IFB; 
 input IFC; 
 input IFD; 
 input IFE; 
 input IFFF ; 
 input IFG; 
 input IFH; 
 input IFI; 
 input IFJ; 
 input IFK; 
 input IFL; 
 input IFM; 
 input IFN; 
 input IFO; 
 input IFP; 
 input IGA; 
 input IGB; 
 input IGC; 
 input IGD; 
 input IGE; 
 input IGF; 
 input IGG; 
 input IGH; 
 input IGI; 
 input IGJ; 
 input IGK; 
 input IGL; 
 input IHA; 
 input IHB; 
 input IHC; 
 input IHD; 
 input IHE; 
 input IHF; 
 input IHG; 
 input IHH; 
 input IHI; 
 input IHJ; 
 input IHK; 
 input IHL; 
 output OAA; 
 output OAB; 
 output OAC; 
 output OAD; 
 output OAE; 
 output OAF; 
 output OAG; 
 output OAH; 
 output OAI; 
 output OAJ; 
 output OAK; 
 output OAL; 
 output OAM; 
 output OAN; 
 output OAO; 
 output OAP; 
 output OAQ; 
 output OAR; 
 output OAS; 
 output OAT; 
 output OBA; 
 output OBB; 
 output OBC; 
 output OBD; 
 output OBE; 
 output OBF; 
 output OBG; 
 output OBH; 
 output OBI; 
 output OBJ; 
 output OBK; 
 output OBL; 
 output OBM; 
 output OBN; 
 output OBO; 
 output OBP; 
 output OBQ; 
 output OBR; 
 output OBS; 
 output OBT; 
 output OCA; 
 output OCB; 
 output OCC; 
 output OCD; 
 output OCE; 
 output OCF; 
 output OCG; 
 output OCH; 
 output OCI; 
 output OCJ; 
 output OCK; 
 output OCL; 
 output OCM; 
 output OCN; 
 output OCO; 
 output OCP; 
 output OCQ; 
 output OCR; 
 output OCS; 
 output OCT; 
 output ODA; 
 output ODB; 
 output ODC; 
 output ODD; 
 output ODE; 
 output ODF; 
 output ODG; 
 output ODH; 
 output ODI; 
 output ODJ; 
 output ODK; 
 output ODL; 
 output ODM; 
 output ODN; 
 output ODO; 
 output ODP; 
 output ODQ; 
 output ODR; 
 output ODS; 
 output ODT; 
 output OEA; 
 output OEB; 
 output OEC; 
 output OED; 
 output OEE; 
 output OEF; 
 output OEG; 
 output OEH; 
 output OEI; 
 output OEJ; 
 output OEK; 
 output OEL; 
 output OEM; 
 output OEN; 
 output OEO; 
 output OEP; 
 output OFA; 
 output OFB; 
 output OFC; 
 output OFD; 
 output OFE; 
 output OFF; 
 output OFG; 
 output OFH; 
 output OFI; 
 output OFJ; 
 output OFK; 
 output OFL; 
 output OFM; 
 output OFN; 
 output OFO; 
 output OFP; 
 output OGA; 
 output OGB; 
 output OGC; 
 output OGD; 
 output OHA; 
  
  
reg  AAA ;
reg  AAB ;
reg  AAC ;
reg  AAD ;
reg  AAE ;
reg  AAF ;
reg  AAG ;
reg  AAH ;
reg  AAI ;
reg  AAJ ;
reg  AAK ;
reg  AAL ;
reg  AAM ;
reg  AAN ;
reg  AAO ;
reg  AAP ;
reg  ABA ;
reg  ABB ;
reg  ABC ;
reg  ABD ;
reg  ABE ;
reg  ABF ;
reg  ABG ;
reg  ABH ;
reg  ABI ;
reg  ABJ ;
reg  ABK ;
reg  ABL ;
reg  ABM ;
reg  ABN ;
reg  ABO ;
reg  ABP ;
reg  ACA ;
reg  ACB ;
reg  ACC ;
reg  ACD ;
reg  ACE ;
reg  ACF ;
reg  ACG ;
reg  ACH ;
reg  ACI ;
reg  ACJ ;
reg  ACK ;
reg  ACL ;
reg  ACM ;
reg  ACN ;
reg  ACO ;
reg  ACP ;
reg  ADA ;
reg  ADB ;
reg  ADC ;
reg  ADD ;
reg  ADE ;
reg  ADF ;
reg  ADG ;
reg  ADH ;
reg  ADI ;
reg  ADJ ;
reg  ADK ;
reg  ADL ;
reg  ADM ;
reg  ADN ;
reg  ADO ;
reg  ADP ;
reg  AEA ;
reg  AEB ;
reg  AEC ;
reg  AED ;
reg  AEE ;
reg  AEF ;
reg  AEG ;
reg  AEH ;
reg  AEI ;
reg  AEJ ;
reg  AEK ;
reg  AEL ;
reg  AEM ;
reg  AEN ;
reg  AEO ;
reg  AEP ;
reg  AFA ;
reg  AFB ;
reg  AFC ;
reg  AFD ;
reg  AFE ;
reg  AFF ;
reg  AFG ;
reg  AFH ;
reg  AFI ;
reg  AFJ ;
reg  AFK ;
reg  AFL ;
reg  AFM ;
reg  AFN ;
reg  AFO ;
reg  AFP ;
reg  BAA ;
reg  BAB ;
reg  BAC ;
reg  BAD ;
reg  BAE ;
reg  BAF ;
reg  BAG ;
reg  BAH ;
reg  BAI ;
reg  BAJ ;
reg  BAK ;
reg  BAL ;
reg  BAM ;
reg  BAN ;
reg  BAO ;
reg  BAP ;
reg  BBA ;
reg  BBB ;
reg  BBC ;
reg  BBD ;
reg  BBE ;
reg  BBF ;
reg  BBG ;
reg  BBH ;
reg  BBI ;
reg  BBJ ;
reg  BBK ;
reg  BBL ;
reg  BBM ;
reg  BBN ;
reg  BBO ;
reg  BBP ;
reg  BCA ;
reg  BCB ;
reg  BCC ;
reg  BCD ;
reg  BCE ;
reg  BCF ;
reg  BCG ;
reg  BCH ;
reg  BCI ;
reg  BCJ ;
reg  BCK ;
reg  BCL ;
reg  BCM ;
reg  BCN ;
reg  BCO ;
reg  BCP ;
reg  BDA ;
reg  BDB ;
reg  BDC ;
reg  BDD ;
reg  BDE ;
reg  BDF ;
reg  BDG ;
reg  BDH ;
reg  BDI ;
reg  BDJ ;
reg  BDK ;
reg  BDL ;
reg  BDM ;
reg  BDN ;
reg  BDO ;
reg  BDP ;
reg  BEA ;
reg  BEB ;
reg  BEC ;
reg  BED ;
reg  BEE ;
reg  BEF ;
reg  BEG ;
reg  BEH ;
reg  BEI ;
reg  BEJ ;
reg  BEK ;
reg  BEL ;
reg  BEM ;
reg  BEN ;
reg  BEO ;
reg  BEP ;
reg  BFA ;
reg  BFB ;
reg  BFC ;
reg  BFD ;
reg  BFE ;
reg  BFF ;
reg  BFG ;
reg  BFH ;
reg  BFI ;
reg  BFJ ;
reg  BFK ;
reg  BFL ;
reg  BFM ;
reg  BFN ;
reg  BFO ;
reg  BFP ;
reg  BGA ;
reg  BGB ;
reg  BGC ;
reg  BGD ;
reg  BGE ;
reg  BGF ;
reg  BGG ;
reg  BGH ;
reg  BGI ;
reg  BGJ ;
reg  BGK ;
reg  BGL ;
reg  BGM ;
reg  BGN ;
reg  BGO ;
reg  BGP ;
reg  BHA ;
reg  BHB ;
reg  BHC ;
reg  BHD ;
reg  BHE ;
reg  BHF ;
reg  BHG ;
reg  BHH ;
reg  BHI ;
reg  BHJ ;
reg  BHK ;
reg  BHL ;
reg  BHM ;
reg  BHN ;
reg  BHO ;
reg  BHP ;
reg  CAA ;
reg  CAB ;
reg  CAC ;
reg  CAD ;
reg  CAE ;
reg  CAF ;
reg  CAG ;
reg  CAH ;
reg  CAI ;
reg  CAJ ;
reg  CAK ;
reg  CAL ;
reg  CAM ;
reg  CAN ;
reg  CAO ;
reg  CAP ;
reg  CBA ;
reg  CBB ;
reg  CBC ;
reg  CBD ;
reg  CBE ;
reg  CBF ;
reg  CBG ;
reg  CBH ;
reg  CBI ;
reg  CBJ ;
reg  CBK ;
reg  CBL ;
reg  CBM ;
reg  CBN ;
reg  CBO ;
reg  CBP ;
reg  CCA ;
reg  CCB ;
reg  CCC ;
reg  CCD ;
reg  CCE ;
reg  CCF ;
reg  CCG ;
reg  CCH ;
reg  CCI ;
reg  CCJ ;
reg  CCK ;
reg  CCL ;
reg  CCM ;
reg  CCN ;
reg  CCO ;
reg  CCP ;
reg  CDA ;
reg  CDB ;
reg  CDC ;
reg  CDD ;
reg  CDE ;
reg  CDF ;
reg  CDG ;
reg  CDH ;
reg  CDI ;
reg  CDJ ;
reg  CDK ;
reg  CDL ;
reg  CDM ;
reg  CDN ;
reg  CDO ;
reg  CDP ;
reg  EAA ;
reg  EAB ;
reg  EAC ;
reg  EAD ;
reg  EAE ;
reg  EAF ;
reg  EAG ;
reg  EAH ;
reg  EAI ;
reg  EAJ ;
reg  EAK ;
reg  EAL ;
reg  gaa ;
reg  gab ;
reg  gac ;
reg  gad ;
reg  gae ;
reg  gaf ;
reg  gag ;
reg  gah ;
reg  gai ;
reg  gaj ;
reg  gak ;
reg  gal ;
reg  gba ;
reg  gbb ;
reg  gbc ;
reg  gbd ;
reg  gbe ;
reg  gbf ;
reg  gbg ;
reg  gbh ;
reg  gbi ;
reg  gbj ;
reg  gbk ;
reg  gbl ;
reg  HAA ;
reg  HAB ;
reg  HAC ;
reg  had ;
reg  hae ;
reg  haf ;
reg  hag ;
reg  HBA ;
reg  HBB ;
reg  HBC ;
reg  KBA ;
reg  KBB ;
reg  KBC ;
reg  KBD ;
reg  KBE ;
reg  KBF ;
reg  KBG ;
reg  KBH ;
reg  KDA ;
reg  LBA ;
reg  LBB ;
reg  LBC ;
reg  LBD ;
reg  LBE ;
reg  LBF ;
reg  LBG ;
reg  LBH ;
reg  LDA ;
reg  OAA ;
reg  OAB ;
reg  OAC ;
reg  OAD ;
reg  OAE ;
reg  OAF ;
reg  OAG ;
reg  OAH ;
reg  OAI ;
reg  OAJ ;
reg  OAK ;
reg  OAL ;
reg  OAM ;
reg  OAN ;
reg  OAO ;
reg  OAP ;
reg  oaq ;
reg  oar ;
reg  oas ;
reg  oat ;
reg  OBA ;
reg  OBB ;
reg  OBC ;
reg  OBD ;
reg  OBE ;
reg  OBF ;
reg  OBG ;
reg  OBH ;
reg  OBI ;
reg  OBJ ;
reg  OBK ;
reg  OBL ;
reg  OBM ;
reg  OBN ;
reg  OBO ;
reg  OBP ;
reg  obq ;
reg  obr ;
reg  obs ;
reg  obt ;
reg  OCA ;
reg  OCB ;
reg  OCC ;
reg  OCD ;
reg  OCE ;
reg  OCF ;
reg  OCG ;
reg  OCH ;
reg  OCI ;
reg  OCJ ;
reg  OCK ;
reg  OCL ;
reg  OCM ;
reg  OCN ;
reg  OCO ;
reg  OCP ;
reg  ocq ;
reg  ocr ;
reg  ocs ;
reg  oct ;
reg  ODA ;
reg  ODB ;
reg  ODC ;
reg  ODD ;
reg  ODE ;
reg  ODF ;
reg  ODG ;
reg  ODH ;
reg  ODI ;
reg  ODJ ;
reg  ODK ;
reg  ODL ;
reg  ODM ;
reg  ODN ;
reg  ODO ;
reg  ODP ;
reg  odq ;
reg  odr ;
reg  ods ;
reg  odt ;
reg  OEA ;
reg  OEB ;
reg  OEC ;
reg  OED ;
reg  OEE ;
reg  OEF ;
reg  OEG ;
reg  OEH ;
reg  OEI ;
reg  OEJ ;
reg  OEK ;
reg  OEL ;
reg  OEM ;
reg  OEN ;
reg  OEO ;
reg  OEP ;
reg  OFA ;
reg  OFB ;
reg  OFC ;
reg  OFD ;
reg  OFE ;
reg  OFF ;
reg  OFG ;
reg  OFH ;
reg  OFI ;
reg  OFJ ;
reg  OFK ;
reg  OFL ;
reg  OFM ;
reg  OFN ;
reg  OFO ;
reg  OFP ;
reg  OGA ;
reg  OGB ;
reg  OGC ;
reg  OGD ;
reg  OHA ;
reg  PAA ;
reg  PAB ;
reg  PAC ;
reg  PAD ;
reg  PAE ;
reg  PAF ;
reg  PAG ;
reg  PAH ;
reg  PAI ;
reg  PAJ ;
reg  PAK ;
reg  PAL ;
reg  PAM ;
reg  PAN ;
reg  PAO ;
reg  PAP ;
reg  PBA ;
reg  PBB ;
reg  PBC ;
reg  PBD ;
reg  PBE ;
reg  PBF ;
reg  PBG ;
reg  PBH ;
reg  PBI ;
reg  PBJ ;
reg  PBK ;
reg  PBL ;
reg  PBM ;
reg  PBN ;
reg  PBO ;
reg  PBP ;
reg  PBQ ;
reg  QAA ;
reg  QAB ;
reg  QAE ;
reg  QAF ;
reg  QAG ;
reg  QAH ;
reg  QAI ;
reg  QAJ ;
reg  QAK ;
reg  QAL ;
reg  qba ;
reg  qbb ;
reg  qbc ;
reg  qbd ;
reg  qbe ;
reg  qbf ;
reg  qbg ;
reg  qbh ;
reg  QCA ;
reg  QCB ;
reg  qcc ;
reg  qcd ;
reg  qce ;
reg  qcf ;
reg  QCG ;
reg  QCH ;
reg  qda ;
reg  qdb ;
reg  qdc ;
reg  qdd ;
reg  QEA ;
reg  QEB ;
reg  QEC ;
reg  QED ;
reg  qee ;
reg  qef ;
reg  qeg ;
reg  qeh ;
reg  QFA ;
reg  QFB ;
reg  QFC ;
reg  QFD ;
reg  qfe ;
reg  qff ;
reg  qfg ;
reg  qfh ;
reg  QGA ;
reg  QGB ;
reg  QGC ;
reg  QGD ;
reg  qge ;
reg  qgf ;
reg  qgg ;
reg  qgh ;
reg  QHA ;
reg  QHB ;
reg  QHC ;
reg  QHD ;
reg  qhe ;
reg  qhf ;
reg  qhg ;
reg  qhh ;
reg  QIA ;
reg  QIB ;
reg  QIC ;
reg  QID ;
reg  QIE ;
reg  QIF ;
reg  QIG ;
reg  QIH ;
reg  QJA ;
reg  QJB ;
reg  QJC ;
reg  QJD ;
reg  QJE ;
reg  QJF ;
reg  QJG ;
reg  QJH ;
reg  QKA ;
reg  QKB ;
reg  QKC ;
reg  QKD ;
reg  QKE ;
reg  QKF ;
reg  QKG ;
reg  QKH ;
reg  QLA ;
reg  QLB ;
reg  QLC ;
reg  QLD ;
reg  QLE ;
reg  QLF ;
reg  QLG ;
reg  QLH ;
reg  qma ;
reg  qmb ;
reg  qmc ;
reg  qmd ;
reg  raa ;
reg  rab ;
reg  rac ;
reg  rad ;
reg  rae ;
reg  raf ;
reg  rag ;
reg  rah ;
reg  rai ;
reg  raj ;
reg  rak ;
reg  ral ;
reg  ram ;
reg  ran ;
reg  rao ;
reg  rap ;
reg  rba ;
reg  rbb ;
reg  rbc ;
reg  rbd ;
reg  rbe ;
reg  rbf ;
reg  rbg ;
reg  rbh ;
reg  rbi ;
reg  rbj ;
reg  rbk ;
reg  rbl ;
reg  rbm ;
reg  rbn ;
reg  rbo ;
reg  rbp ;
reg  rca ;
reg  rcb ;
reg  rcc ;
reg  rcd ;
reg  rce ;
reg  rcf ;
reg  rcg ;
reg  rch ;
reg  rci ;
reg  rcj ;
reg  rck ;
reg  rcl ;
reg  rcm ;
reg  rcn ;
reg  rco ;
reg  rcp ;
reg  rda ;
reg  rdb ;
reg  rdc ;
reg  rdd ;
reg  rde ;
reg  rdf ;
reg  rdg ;
reg  rdh ;
reg  rdi ;
reg  rdj ;
reg  rdk ;
reg  rdl ;
reg  rdm ;
reg  rdn ;
reg  rdo ;
reg  TBA ;
reg  TBB ;
reg  TBC ;
reg  TBD ;
reg  TBE ;
reg  TBF ;
reg  TBG ;
reg  TBH ;
reg  TDA ;
reg  TDB ;
reg  TDC ;
reg  TDD ;
reg  WAA ;
reg  WAB ;
reg  WAC ;
reg  WAD ;
reg  WAE ;
reg  WAF ;
reg  WAG ;
reg  WAH ;
reg  WBA ;
wire  aaa ;
wire  aab ;
wire  aac ;
wire  aad ;
wire  aae ;
wire  aaf ;
wire  aag ;
wire  aah ;
wire  aai ;
wire  aaj ;
wire  aak ;
wire  aal ;
wire  aam ;
wire  aan ;
wire  aao ;
wire  aap ;
wire  aba ;
wire  abb ;
wire  abc ;
wire  abd ;
wire  abe ;
wire  abf ;
wire  abg ;
wire  abh ;
wire  abi ;
wire  abj ;
wire  abk ;
wire  abl ;
wire  abm ;
wire  abn ;
wire  abo ;
wire  abp ;
wire  aca ;
wire  acb ;
wire  acc ;
wire  acd ;
wire  ace ;
wire  acf ;
wire  acg ;
wire  ach ;
wire  aci ;
wire  acj ;
wire  ack ;
wire  acl ;
wire  acm ;
wire  acn ;
wire  aco ;
wire  acp ;
wire  ada ;
wire  adb ;
wire  adc ;
wire  add ;
wire  ade ;
wire  adf ;
wire  adg ;
wire  adh ;
wire  adi ;
wire  adj ;
wire  adk ;
wire  adl ;
wire  adm ;
wire  adn ;
wire  ado ;
wire  adp ;
wire  aea ;
wire  aeb ;
wire  aec ;
wire  aed ;
wire  aee ;
wire  aef ;
wire  aeg ;
wire  aeh ;
wire  aei ;
wire  aej ;
wire  aek ;
wire  ael ;
wire  aem ;
wire  aen ;
wire  aeo ;
wire  aep ;
wire  afa ;
wire  afb ;
wire  afc ;
wire  afd ;
wire  afe ;
wire  aff ;
wire  afg ;
wire  afh ;
wire  afi ;
wire  afj ;
wire  afk ;
wire  afl ;
wire  afm ;
wire  afn ;
wire  afo ;
wire  afp ;
wire  baa ;
wire  bab ;
wire  bac ;
wire  bad ;
wire  bae ;
wire  baf ;
wire  bag ;
wire  bah ;
wire  bai ;
wire  baj ;
wire  bak ;
wire  bal ;
wire  bam ;
wire  ban ;
wire  bao ;
wire  bap ;
wire  bba ;
wire  bbb ;
wire  bbc ;
wire  bbd ;
wire  bbe ;
wire  bbf ;
wire  bbg ;
wire  bbh ;
wire  bbi ;
wire  bbj ;
wire  bbk ;
wire  bbl ;
wire  bbm ;
wire  bbn ;
wire  bbo ;
wire  bbp ;
wire  bca ;
wire  bcb ;
wire  bcc ;
wire  bcd ;
wire  bce ;
wire  bcf ;
wire  bcg ;
wire  bch ;
wire  bci ;
wire  bcj ;
wire  bck ;
wire  bcl ;
wire  bcm ;
wire  bcn ;
wire  bco ;
wire  bcp ;
wire  bda ;
wire  bdb ;
wire  bdc ;
wire  bdd ;
wire  bde ;
wire  bdf ;
wire  bdg ;
wire  bdh ;
wire  bdi ;
wire  bdj ;
wire  bdk ;
wire  bdl ;
wire  bdm ;
wire  bdn ;
wire  bdo ;
wire  bdp ;
wire  bea ;
wire  beb ;
wire  bec ;
wire  bed ;
wire  bee ;
wire  bef ;
wire  beg ;
wire  beh ;
wire  bei ;
wire  bej ;
wire  bek ;
wire  bel ;
wire  bem ;
wire  ben ;
wire  beo ;
wire  bep ;
wire  bfa ;
wire  bfb ;
wire  bfc ;
wire  bfd ;
wire  bfe ;
wire  bff ;
wire  bfg ;
wire  bfh ;
wire  bfi ;
wire  bfj ;
wire  bfk ;
wire  bfl ;
wire  bfm ;
wire  bfn ;
wire  bfo ;
wire  bfp ;
wire  bga ;
wire  bgb ;
wire  bgc ;
wire  bgd ;
wire  bge ;
wire  bgf ;
wire  bgg ;
wire  bgh ;
wire  bgi ;
wire  bgj ;
wire  bgk ;
wire  bgl ;
wire  bgm ;
wire  bgn ;
wire  bgo ;
wire  bgp ;
wire  bha ;
wire  bhb ;
wire  bhc ;
wire  bhd ;
wire  bhe ;
wire  bhf ;
wire  bhg ;
wire  bhh ;
wire  bhi ;
wire  bhj ;
wire  bhk ;
wire  bhl ;
wire  bhm ;
wire  bhn ;
wire  bho ;
wire  bhp ;
wire  caa ;
wire  cab ;
wire  cac ;
wire  cad ;
wire  cae ;
wire  caf ;
wire  cag ;
wire  cah ;
wire  cai ;
wire  caj ;
wire  cak ;
wire  cal ;
wire  cam ;
wire  can ;
wire  cao ;
wire  cap ;
wire  cba ;
wire  cbb ;
wire  cbc ;
wire  cbd ;
wire  cbe ;
wire  cbf ;
wire  cbg ;
wire  cbh ;
wire  cbi ;
wire  cbj ;
wire  cbk ;
wire  cbl ;
wire  cbm ;
wire  cbn ;
wire  cbo ;
wire  cbp ;
wire  cca ;
wire  ccb ;
wire  ccc ;
wire  ccd ;
wire  cce ;
wire  ccf ;
wire  ccg ;
wire  cch ;
wire  cci ;
wire  ccj ;
wire  cck ;
wire  ccl ;
wire  ccm ;
wire  ccn ;
wire  cco ;
wire  ccp ;
wire  cda ;
wire  cdb ;
wire  cdc ;
wire  cdd ;
wire  cde ;
wire  cdf ;
wire  cdg ;
wire  cdh ;
wire  cdi ;
wire  cdj ;
wire  cdk ;
wire  cdl ;
wire  cdm ;
wire  cdn ;
wire  cdo ;
wire  cdp ;
wire  daa ;
wire  DAA ;
wire  dab ;
wire  DAB ;
wire  dac ;
wire  DAC ;
wire  dad ;
wire  DAD ;
wire  dae ;
wire  DAE ;
wire  daf ;
wire  DAF ;
wire  dag ;
wire  DAG ;
wire  dah ;
wire  DAH ;
wire  dai ;
wire  DAI ;
wire  daj ;
wire  DAJ ;
wire  dak ;
wire  DAK ;
wire  dal ;
wire  DAL ;
wire  dam ;
wire  DAM ;
wire  dan ;
wire  DAN ;
wire  dao ;
wire  DAO ;
wire  dap ;
wire  DAP ;
wire  dba ;
wire  DBA ;
wire  dbb ;
wire  DBB ;
wire  dbc ;
wire  DBC ;
wire  dbd ;
wire  DBD ;
wire  dbe ;
wire  DBE ;
wire  dbf ;
wire  DBF ;
wire  dbg ;
wire  DBG ;
wire  dbh ;
wire  DBH ;
wire  dbi ;
wire  DBI ;
wire  dbj ;
wire  DBJ ;
wire  dbk ;
wire  DBK ;
wire  dbl ;
wire  DBL ;
wire  dbm ;
wire  DBM ;
wire  dbn ;
wire  DBN ;
wire  dbo ;
wire  DBO ;
wire  dbp ;
wire  DBP ;
wire  eaa ;
wire  eab ;
wire  eac ;
wire  ead ;
wire  eae ;
wire  eaf ;
wire  eag ;
wire  eah ;
wire  eai ;
wire  eaj ;
wire  eak ;
wire  eal ;
wire  eba ;
wire  EBA ;
wire  ebb ;
wire  EBB ;
wire  ebc ;
wire  EBC ;
wire  ebd ;
wire  EBD ;
wire  ebe ;
wire  EBE ;
wire  ebf ;
wire  EBF ;
wire  ebg ;
wire  EBG ;
wire  ebh ;
wire  EBH ;
wire  ebi ;
wire  EBI ;
wire  ebj ;
wire  EBJ ;
wire  ebk ;
wire  EBK ;
wire  ebl ;
wire  EBL ;
wire  faa ;
wire  FAA ;
wire  fab ;
wire  FAB ;
wire  fac ;
wire  FAC ;
wire  fad ;
wire  FAD ;
wire  fae ;
wire  FAE ;
wire  faf ;
wire  FAF ;
wire  fag ;
wire  FAG ;
wire  fah ;
wire  FAH ;
wire  fba ;
wire  FBA ;
wire  fbb ;
wire  FBB ;
wire  fbc ;
wire  FBC ;
wire  fbd ;
wire  FBD ;
wire  fbe ;
wire  FBE ;
wire  fbf ;
wire  FBF ;
wire  fbg ;
wire  FBG ;
wire  fbh ;
wire  FBH ;
wire  fca ;
wire  FCA ;
wire  fcb ;
wire  FCB ;
wire  fcc ;
wire  FCC ;
wire  fcd ;
wire  FCD ;
wire  fce ;
wire  FCE ;
wire  fcf ;
wire  FCF ;
wire  fcg ;
wire  FCG ;
wire  fch ;
wire  FCH ;
wire  fda ;
wire  FDA ;
wire  fdb ;
wire  FDB ;
wire  fdc ;
wire  FDC ;
wire  fdd ;
wire  FDD ;
wire  fde ;
wire  FDE ;
wire  fdf ;
wire  FDF ;
wire  fdg ;
wire  FDG ;
wire  fdh ;
wire  FDH ;
wire  fea ;
wire  FEA ;
wire  feb ;
wire  FEB ;
wire  fec ;
wire  FEC ;
wire  fed ;
wire  FED ;
wire  fee ;
wire  FEE ;
wire  fef ;
wire  FEF ;
wire  feg ;
wire  FEG ;
wire  feh ;
wire  FEH ;
wire  ffa ;
wire  FFA ;
wire  ffb ;
wire  FFB ;
wire  ffc ;
wire  FFC ;
wire  ffd ;
wire  FFD ;
wire  ffe ;
wire  FFE ;
wire  fff ;
wire  FFF ;
wire  ffg ;
wire  FFG ;
wire  ffh ;
wire  FFH ;
wire  fga ;
wire  FGA ;
wire  fgb ;
wire  FGB ;
wire  fgc ;
wire  FGC ;
wire  fgd ;
wire  FGD ;
wire  fge ;
wire  FGE ;
wire  fgf ;
wire  FGF ;
wire  fgg ;
wire  FGG ;
wire  fgh ;
wire  FGH ;
wire  fha ;
wire  FHA ;
wire  fhb ;
wire  FHB ;
wire  fhc ;
wire  FHC ;
wire  fhd ;
wire  FHD ;
wire  fhe ;
wire  FHE ;
wire  fhf ;
wire  FHF ;
wire  fhg ;
wire  FHG ;
wire  fhh ;
wire  FHH ;
wire  fia ;
wire  FIA ;
wire  fib ;
wire  FIB ;
wire  fic ;
wire  FIC ;
wire  fid ;
wire  FID ;
wire  fie ;
wire  FIE ;
wire  fif ;
wire  FIF ;
wire  fig ;
wire  FIG ;
wire  fih ;
wire  FIH ;
wire  fja ;
wire  FJA ;
wire  fjb ;
wire  FJB ;
wire  fjc ;
wire  FJC ;
wire  fjd ;
wire  FJD ;
wire  fje ;
wire  FJE ;
wire  fjf ;
wire  FJF ;
wire  fjg ;
wire  FJG ;
wire  fjh ;
wire  FJH ;
wire  fka ;
wire  FKA ;
wire  fkb ;
wire  FKB ;
wire  fkc ;
wire  FKC ;
wire  fkd ;
wire  FKD ;
wire  fke ;
wire  FKE ;
wire  fkf ;
wire  FKF ;
wire  fkg ;
wire  FKG ;
wire  fkh ;
wire  FKH ;
wire  fla ;
wire  FLA ;
wire  flb ;
wire  FLB ;
wire  flc ;
wire  FLC ;
wire  fld ;
wire  FLD ;
wire  fle ;
wire  FLE ;
wire  flf ;
wire  FLF ;
wire  flg ;
wire  FLG ;
wire  flh ;
wire  FLH ;
wire  fma ;
wire  FMA ;
wire  fmb ;
wire  FMB ;
wire  fmc ;
wire  FMC ;
wire  fmd ;
wire  FMD ;
wire  fme ;
wire  FME ;
wire  fmf ;
wire  FMF ;
wire  fmg ;
wire  FMG ;
wire  fmh ;
wire  FMH ;
wire  fmi ;
wire  FMI ;
wire  fmj ;
wire  FMJ ;
wire  fmk ;
wire  FMK ;
wire  fml ;
wire  FML ;
wire  GAA ;
wire  GAB ;
wire  GAC ;
wire  GAD ;
wire  GAE ;
wire  GAF ;
wire  GAG ;
wire  GAH ;
wire  GAI ;
wire  GAJ ;
wire  GAK ;
wire  GAL ;
wire  GBA ;
wire  GBB ;
wire  GBC ;
wire  GBD ;
wire  GBE ;
wire  GBF ;
wire  GBG ;
wire  GBH ;
wire  GBI ;
wire  GBJ ;
wire  GBK ;
wire  GBL ;
wire  haa ;
wire  hab ;
wire  hac ;
wire  HAD ;
wire  HAE ;
wire  HAF ;
wire  HAG ;
wire  hba ;
wire  hbb ;
wire  hbc ;
wire  iaa ;
wire  iab ;
wire  iac ;
wire  iad ;
wire  iae ;
wire  iaf ;
wire  iag ;
wire  iah ;
wire  iai ;
wire  iaj ;
wire  iak ;
wire  ial ;
wire  iam ;
wire  ian ;
wire  iao ;
wire  iap ;
wire  iaq ;
wire  ias ;
wire  iat ;
wire  iba ;
wire  ibb ;
wire  ibc ;
wire  ibd ;
wire  ibe ;
wire  ibf ;
wire  ibg ;
wire  ibh ;
wire  ibi ;
wire  ibj ;
wire  ibk ;
wire  ibl ;
wire  ibm ;
wire  ibn ;
wire  ibo ;
wire  ibp ;
wire  ibq ;
wire  ibs ;
wire  ibt ;
wire  ica ;
wire  icb ;
wire  icc ;
wire  icd ;
wire  ice ;
wire  icf ;
wire  icg ;
wire  ich ;
wire  ici ;
wire  icj ;
wire  ick ;
wire  icl ;
wire  icm ;
wire  icn ;
wire  ico ;
wire  icp ;
wire  icq ;
wire  ics ;
wire  ict ;
wire  ida ;
wire  idb ;
wire  idc ;
wire  idd ;
wire  ide ;
wire  idf ;
wire  idg ;
wire  idh ;
wire  idi ;
wire  idj ;
wire  idk ;
wire  idl ;
wire  idm ;
wire  idn ;
wire  ido ;
wire  idp ;
wire  idq ;
wire  ids ;
wire  idt ;
wire  iea ;
wire  ieb ;
wire  iec ;
wire  ied ;
wire  iee ;
wire  ief ;
wire  ieg ;
wire  ieh ;
wire  iei ;
wire  iej ;
wire  iek ;
wire  iel ;
wire  iem ;
wire  ien ;
wire  ieo ;
wire  iep ;
wire  ifa ;
wire  ifb ;
wire  ifc ;
wire  ifd ;
wire  ife ;
wire  ifff  ;
wire  ifg ;
wire  ifh ;
wire  ifi ;
wire  ifj ;
wire  ifk ;
wire  ifl ;
wire  ifm ;
wire  ifn ;
wire  ifo ;
wire  ifp ;
wire  iga ;
wire  igb ;
wire  igc ;
wire  igd ;
wire  ige ;
wire  igf ;
wire  igg ;
wire  igh ;
wire  igi ;
wire  igj ;
wire  igk ;
wire  igl ;
wire  iha ;
wire  ihb ;
wire  ihc ;
wire  ihd ;
wire  ihe ;
wire  ihf ;
wire  ihg ;
wire  ihh ;
wire  ihi ;
wire  ihj ;
wire  ihk ;
wire  ihl ;
wire  jab ;
wire  JAB ;
wire  jac ;
wire  JAC ;
wire  jad ;
wire  JAD ;
wire  jae ;
wire  JAE ;
wire  jaf ;
wire  JAF ;
wire  jag ;
wire  JAG ;
wire  jah ;
wire  JAH ;
wire  jai ;
wire  JAI ;
wire  jaj ;
wire  JAJ ;
wire  jak ;
wire  JAK ;
wire  jal ;
wire  JAL ;
wire  jam ;
wire  JAM ;
wire  jan ;
wire  JAN ;
wire  jao ;
wire  JAO ;
wire  jap ;
wire  JAP ;
wire  jaq ;
wire  JAQ ;
wire  jar ;
wire  JAR ;
wire  jas ;
wire  JAS ;
wire  jat ;
wire  JAT ;
wire  jba ;
wire  JBA ;
wire  jbb ;
wire  JBB ;
wire  jbc ;
wire  JBC ;
wire  jbd ;
wire  JBD ;
wire  jbe ;
wire  JBE ;
wire  jbf ;
wire  JBF ;
wire  jbg ;
wire  JBG ;
wire  jbh ;
wire  JBH ;
wire  jbi ;
wire  JBI ;
wire  jbj ;
wire  JBJ ;
wire  jbk ;
wire  JBK ;
wire  jbl ;
wire  JBL ;
wire  jbm ;
wire  JBM ;
wire  jbn ;
wire  JBN ;
wire  jbo ;
wire  JBO ;
wire  jbp ;
wire  JBP ;
wire  jbq ;
wire  JBQ ;
wire  jbr ;
wire  JBR ;
wire  jbs ;
wire  JBS ;
wire  jca ;
wire  JCA ;
wire  jcb ;
wire  JCB ;
wire  jcc ;
wire  JCC ;
wire  jcd ;
wire  JCD ;
wire  jce ;
wire  JCE ;
wire  kaa ;
wire  KAA ;
wire  kab ;
wire  KAB ;
wire  kac ;
wire  KAC ;
wire  kad ;
wire  KAD ;
wire  kae ;
wire  KAE ;
wire  kaf ;
wire  KAF ;
wire  kag ;
wire  KAG ;
wire  kah ;
wire  KAH ;
wire  kai ;
wire  KAI ;
wire  kaj ;
wire  KAJ ;
wire  kak ;
wire  KAK ;
wire  kal ;
wire  KAL ;
wire  kam ;
wire  KAM ;
wire  kan ;
wire  KAN ;
wire  kao ;
wire  KAO ;
wire  kap ;
wire  KAP ;
wire  kba ;
wire  kbb ;
wire  kbc ;
wire  kbd ;
wire  kbe ;
wire  kbf ;
wire  kbg ;
wire  kbh ;
wire  kca ;
wire  KCA ;
wire  kcb ;
wire  KCB ;
wire  kcc ;
wire  KCC ;
wire  kda ;
wire  laa ;
wire  LAA ;
wire  lab ;
wire  LAB ;
wire  lac ;
wire  LAC ;
wire  lad ;
wire  LAD ;
wire  lae ;
wire  LAE ;
wire  laf ;
wire  LAF ;
wire  lag ;
wire  LAG ;
wire  lah ;
wire  LAH ;
wire  lai ;
wire  LAI ;
wire  laj ;
wire  LAJ ;
wire  lak ;
wire  LAK ;
wire  lal ;
wire  LAL ;
wire  lam ;
wire  LAM ;
wire  lan ;
wire  LAN ;
wire  lao ;
wire  LAO ;
wire  lap ;
wire  LAP ;
wire  lba ;
wire  lbb ;
wire  lbc ;
wire  lbd ;
wire  lbe ;
wire  lbf ;
wire  lbg ;
wire  lbh ;
wire  lca ;
wire  LCA ;
wire  lcb ;
wire  LCB ;
wire  lcc ;
wire  LCC ;
wire  lda ;
wire  lea ;
wire  LEA ;
wire  oaa ;
wire  oab ;
wire  oac ;
wire  oad ;
wire  oae ;
wire  oaf ;
wire  oag ;
wire  oah ;
wire  oai ;
wire  oaj ;
wire  oak ;
wire  oal ;
wire  oam ;
wire  oan ;
wire  oao ;
wire  oap ;
wire  OAQ ;
wire  OAR ;
wire  OAS ;
wire  OAT ;
wire  oba ;
wire  obb ;
wire  obc ;
wire  obd ;
wire  obe ;
wire  obf ;
wire  obg ;
wire  obh ;
wire  obi ;
wire  obj ;
wire  obk ;
wire  obl ;
wire  obm ;
wire  obn ;
wire  obo ;
wire  obp ;
wire  OBQ ;
wire  OBR ;
wire  OBS ;
wire  OBT ;
wire  oca ;
wire  ocb ;
wire  occ ;
wire  ocd ;
wire  oce ;
wire  ocf ;
wire  ocg ;
wire  och ;
wire  oci ;
wire  ocj ;
wire  ock ;
wire  ocl ;
wire  ocm ;
wire  ocn ;
wire  oco ;
wire  ocp ;
wire  OCQ ;
wire  OCR ;
wire  OCS ;
wire  OCT ;
wire  oda ;
wire  odb ;
wire  odc ;
wire  odd ;
wire  ode ;
wire  odf ;
wire  odg ;
wire  odh ;
wire  odi ;
wire  odj ;
wire  odk ;
wire  odl ;
wire  odm ;
wire  odn ;
wire  odo ;
wire  odp ;
wire  ODQ ;
wire  ODR ;
wire  ODS ;
wire  ODT ;
wire  oea ;
wire  oeb ;
wire  oec ;
wire  oed ;
wire  oee ;
wire  oef ;
wire  oeg ;
wire  oeh ;
wire  oei ;
wire  oej ;
wire  oek ;
wire  oel ;
wire  oem ;
wire  oen ;
wire  oeo ;
wire  oep ;
wire  ofa ;
wire  ofb ;
wire  ofc ;
wire  ofd ;
wire  ofe ;
wire  off ;
wire  ofg ;
wire  ofh ;
wire  ofi ;
wire  ofj ;
wire  ofk ;
wire  ofl ;
wire  ofm ;
wire  ofn ;
wire  ofo ;
wire  ofp ;
wire  oga ;
wire  ogb ;
wire  ogc ;
wire  ogd ;
wire  oha ;
wire  paa ;
wire  pab ;
wire  pac ;
wire  pad ;
wire  pae ;
wire  paf ;
wire  pag ;
wire  pah ;
wire  pai ;
wire  paj ;
wire  pak ;
wire  pal ;
wire  pam ;
wire  pan ;
wire  pao ;
wire  pap ;
wire  pba ;
wire  pbb ;
wire  pbc ;
wire  pbd ;
wire  pbe ;
wire  pbf ;
wire  pbg ;
wire  pbh ;
wire  pbi ;
wire  pbj ;
wire  pbk ;
wire  pbl ;
wire  pbm ;
wire  pbn ;
wire  pbo ;
wire  pbp ;
wire  pbq ;
wire  qaa ;
wire  qab ;
wire  qae ;
wire  qaf ;
wire  qag ;
wire  qah ;
wire  qai ;
wire  qaj ;
wire  qak ;
wire  qal ;
wire  QBA ;
wire  QBB ;
wire  QBC ;
wire  QBD ;
wire  QBE ;
wire  QBF ;
wire  QBG ;
wire  QBH ;
wire  qca ;
wire  qcb ;
wire  QCC ;
wire  QCD ;
wire  QCE ;
wire  QCF ;
wire  qcg ;
wire  qch ;
wire  QDA ;
wire  QDB ;
wire  QDC ;
wire  QDD ;
wire  qea ;
wire  qeb ;
wire  qec ;
wire  qed ;
wire  QEE ;
wire  QEF ;
wire  QEG ;
wire  QEH ;
wire  qfa ;
wire  qfb ;
wire  qfc ;
wire  qfd ;
wire  QFE ;
wire  QFF ;
wire  QFG ;
wire  QFH ;
wire  qga ;
wire  qgb ;
wire  qgc ;
wire  qgd ;
wire  QGE ;
wire  QGF ;
wire  QGG ;
wire  QGH ;
wire  qha ;
wire  qhb ;
wire  qhc ;
wire  qhd ;
wire  QHE ;
wire  QHF ;
wire  QHG ;
wire  QHH ;
wire  qia ;
wire  qib ;
wire  qic ;
wire  qid ;
wire  qie ;
wire  qif ;
wire  qig ;
wire  qih ;
wire  qja ;
wire  qjb ;
wire  qjc ;
wire  qjd ;
wire  qje ;
wire  qjf ;
wire  qjg ;
wire  qjh ;
wire  qka ;
wire  qkb ;
wire  qkc ;
wire  qkd ;
wire  qke ;
wire  qkf ;
wire  qkg ;
wire  qkh ;
wire  qla ;
wire  qlb ;
wire  qlc ;
wire  qld ;
wire  qle ;
wire  qlf ;
wire  qlg ;
wire  qlh ;
wire  QMA ;
wire  QMB ;
wire  QMC ;
wire  QMD ;
wire  RAA ;
wire  RAB ;
wire  RAC ;
wire  RAD ;
wire  RAE ;
wire  RAF ;
wire  RAG ;
wire  RAH ;
wire  RAI ;
wire  RAJ ;
wire  RAK ;
wire  RAL ;
wire  RAM ;
wire  RAN ;
wire  RAO ;
wire  RAP ;
wire  RBA ;
wire  RBB ;
wire  RBC ;
wire  RBD ;
wire  RBE ;
wire  RBF ;
wire  RBG ;
wire  RBH ;
wire  RBI ;
wire  RBJ ;
wire  RBK ;
wire  RBL ;
wire  RBM ;
wire  RBN ;
wire  RBO ;
wire  RBP ;
wire  RCA ;
wire  RCB ;
wire  RCC ;
wire  RCD ;
wire  RCE ;
wire  RCF ;
wire  RCG ;
wire  RCH ;
wire  RCI ;
wire  RCJ ;
wire  RCK ;
wire  RCL ;
wire  RCM ;
wire  RCN ;
wire  RCO ;
wire  RCP ;
wire  RDA ;
wire  RDB ;
wire  RDC ;
wire  RDD ;
wire  RDE ;
wire  RDF ;
wire  RDG ;
wire  RDH ;
wire  RDI ;
wire  RDJ ;
wire  RDK ;
wire  RDL ;
wire  RDM ;
wire  RDN ;
wire  RDO ;
wire  taa ;
wire  TAA ;
wire  tab ;
wire  TAB ;
wire  tac ;
wire  TAC ;
wire  tad ;
wire  TAD ;
wire  tba ;
wire  tbb ;
wire  tbc ;
wire  tbd ;
wire  tbe ;
wire  tbf ;
wire  tbg ;
wire  tbh ;
wire  tca ;
wire  TCA ;
wire  tcb ;
wire  TCB ;
wire  tcc ;
wire  TCC ;
wire  tcd ;
wire  TCD ;
wire  tce ;
wire  TCE ;
wire  tcf ;
wire  TCF ;
wire  tcg ;
wire  TCG ;
wire  tch ;
wire  TCH ;
wire  tci ;
wire  TCI ;
wire  tcj ;
wire  TCJ ;
wire  tck ;
wire  TCK ;
wire  tcl ;
wire  TCL ;
wire  tcm ;
wire  TCM ;
wire  tcn ;
wire  TCN ;
wire  tco ;
wire  TCO ;
wire  tcp ;
wire  TCP ;
wire  tcq ;
wire  TCQ ;
wire  tcr ;
wire  TCR ;
wire  tcs ;
wire  TCS ;
wire  tct ;
wire  TCT ;
wire  tcu ;
wire  TCU ;
wire  tcv ;
wire  TCV ;
wire  tcw ;
wire  TCW ;
wire  tcx ;
wire  TCX ;
wire  tda ;
wire  tdb ;
wire  tdc ;
wire  tdd ;
wire  tde ;
wire  TDE ;
wire  tdf ;
wire  TDF ;
wire  tdg ;
wire  TDG ;
wire  tdh ;
wire  TDH ;
wire  tdi ;
wire  TDI ;
wire  tdj ;
wire  TDJ ;
wire  tdk ;
wire  TDK ;
wire  tdl ;
wire  TDL ;
wire  tea ;
wire  TEA ;
wire  teb ;
wire  TEB ;
wire  tec ;
wire  TEC ;
wire  waa ;
wire  wab ;
wire  wac ;
wire  wad ;
wire  wae ;
wire  waf ;
wire  wag ;
wire  wah ;
wire  wba ;
wire  ZZI ;
wire  ZZO ;
assign ZZI = 1'b1;
assign ZZO = 1'b0;
assign FAA = EAA; 
assign faa = ~FAA; //complement 
assign FBA = EAB; 
assign fba = ~FBA;  //complement 
assign FCA = EAC; 
assign fca = ~FCA;  //complement 
assign FDA = EAD; 
assign fda = ~FDA;  //complement 
assign FEA = EAE; 
assign fea = ~FEA; //complement 
assign FFA = EAF; 
assign ffa = ~FFA;  //complement 
assign FGA = EAG; 
assign fga = ~FGA;  //complement 
assign FHA = EAH; 
assign fha = ~FHA;  //complement 
assign FIA = EAI; 
assign fia = ~FIA; //complement 
assign FJA = EAJ; 
assign fja = ~FJA;  //complement 
assign FKA = EAK; 
assign fka = ~FKA;  //complement 
assign FLA = EAL; 
assign fla = ~FLA;  //complement 
assign waa = ~WAA;  //complement 
assign GAA = ~gaa;  //complement 
assign GAB = ~gab;  //complement 
assign GAC = ~gac;  //complement 
assign GAD = ~gad;  //complement 
assign GBA = ~gba;  //complement 
assign GBB = ~gbb;  //complement 
assign GBC = ~gbc;  //complement 
assign GBD = ~gbd;  //complement 
assign GAE = ~gae;  //complement 
assign GAF = ~gaf;  //complement 
assign GAG = ~gag;  //complement 
assign GAH = ~gah;  //complement 
assign GBE = ~gbe;  //complement 
assign GBF = ~gbf;  //complement 
assign GBG = ~gbg;  //complement 
assign GBH = ~gbh;  //complement 
assign JAI =  HAB  ; 
assign jai = ~JAI;  //complement  
assign GAI = ~gai;  //complement 
assign GAJ = ~gaj;  //complement 
assign GAK = ~gak;  //complement 
assign GAL = ~gal;  //complement 
assign GBI = ~gbi;  //complement 
assign GBJ = ~gbj;  //complement 
assign GBK = ~gbk;  //complement 
assign GBL = ~gbl;  //complement 
assign kba = ~KBA;  //complement 
assign FMA =  GBA  ; 
assign fma = ~FMA;  //complement 
assign FMB =  GBB  ; 
assign fmb = ~FMB;  //complement 
assign FMC =  GBC  ; 
assign fmc = ~FMC;  //complement 
assign FMD =  GBD  ; 
assign fmd = ~FMD;  //complement 
assign lba = ~LBA;  //complement 
assign FME =  GBE  ; 
assign fme = ~FME;  //complement 
assign FMF =  GBF  ; 
assign fmf = ~FMF;  //complement 
assign FMG =  GBG  ; 
assign fmg = ~FMG;  //complement 
assign FMH =  GBH  ; 
assign fmh = ~FMH;  //complement 
assign JBA =  HAD  ; 
assign jba = ~JBA;  //complement  
assign wba = ~WBA;  //complement 
assign FMI =  GBI  ; 
assign fmi = ~FMI;  //complement 
assign FMJ =  GBJ  ; 
assign fmj = ~FMJ;  //complement 
assign FMK =  GBK  ; 
assign fmk = ~FMK;  //complement 
assign FML =  GBL  ; 
assign fml = ~FML;  //complement 
assign JBI =  HAF & HBB  ; 
assign jbi = ~JBI;  //complement  
assign RAA = ~raa;  //complement 
assign RCA = ~rca;  //complement 
assign oea = ~OEA;  //complement 
assign paa = ~PAA;  //complement 
assign DAA =  BAA & QEA  |  BCA & QFA  |  BEA & QGA  |  BGA & QHA  ; 
assign daa = ~DAA;  //complement 
assign aaa = ~AAA;  //complement 
assign aca = ~ACA;  //complement 
assign aea = ~AEA;  //complement 
assign eba = eaa; 
assign EBA = ~eba; //complement 
assign ebi = eai; 
assign EBI = ~ebi;  //complement 
assign TAA = QAL; 
assign taa = ~TAA;  //complement 
assign TAB = QAL; 
assign tab = ~TAB;  //complement 
assign RAI = ~rai;  //complement 
assign RCI = ~rci;  //complement 
assign oei = ~OEI;  //complement 
assign pai = ~PAI;  //complement 
assign DAI =  BAI & QEC  |  BCI & QFC  |  BEI & QGC  |  BGI & QHC  ; 
assign dai = ~DAI;  //complement 
assign KAA =  AEA & aei  |  aea & AEI  |  aea & aei  |  AEA & AEI  ; 
assign kaa = ~KAA; //complement 
assign KAI =  AFA & afi  |  afa & AFI  |  afa & afi  |  AFA & AFI  ; 
assign kai = ~KAI; //complement 
assign aai = ~AAI;  //complement 
assign aci = ~ACI;  //complement 
assign aei = ~AEI;  //complement 
assign qal = ~QAL;  //complement 
assign LAA =  PAA & pai  |  paa & PAI  |  paa & pai  |  PAA & PAI  ; 
assign laa = ~LAA; //complement 
assign LAI =  PBA & pbi  |  pba & PBI  |  pba & pbi  |  PBA & PBI  ; 
assign lai = ~LAI; //complement 
assign aba = ~ABA;  //complement 
assign ada = ~ADA;  //complement 
assign afa = ~AFA;  //complement 
assign RBA = ~rba;  //complement 
assign RDA = ~rda;  //complement 
assign ofa = ~OFA;  //complement 
assign pba = ~PBA;  //complement 
assign DBA =  BBA & QEE  |  BDA & QFE  |  BFA & QGE  |  BHA & QHE  ; 
assign dba = ~DBA;  //complement 
assign abi = ~ABI;  //complement 
assign adi = ~ADI;  //complement 
assign afi = ~AFI;  //complement 
assign tac = qal; 
assign TAC = ~tac; //complement 
assign tad = qal; 
assign TAD = ~tad;  //complement 
assign RBI = ~rbi;  //complement 
assign RDI = ~rdi;  //complement 
assign ofi = ~OFI;  //complement 
assign pbi = ~PBI;  //complement 
assign DBI =  BBI & QEG  |  BDI & QFG  |  BFI & QGG  |  BHI & QHG  ; 
assign dbi = ~DBI;  //complement 
assign baa = ~BAA;  //complement 
assign bai = ~BAI;  //complement 
assign bba = ~BBA;  //complement 
assign bbi = ~BBI;  //complement 
assign caa = ~CAA;  //complement 
assign oaa = ~OAA;  //complement 
assign cai = ~CAI;  //complement 
assign oai = ~OAI;  //complement 
assign eaa = ~EAA;  //complement 
assign eai = ~EAI;  //complement 
assign tcc = qie & qic ; 
assign TCC = ~tcc ; //complement 
assign tcd = qie & qic ; 
assign TCD = ~tcd ;  //complement 
assign tce = qif & qid ; 
assign TCE = ~tce ;  //complement 
assign tcf = qif & qid; 
assign TCF = ~tcf; 
assign tca = QIB; 
assign TCA = ~tca; //complement 
assign tcb = QIB; 
assign TCB = ~tcb;  //complement 
assign bca = ~BCA;  //complement 
assign bci = ~BCI;  //complement 
assign bda = ~BDA;  //complement 
assign bdi = ~BDI;  //complement 
assign cba = ~CBA;  //complement 
assign oba = ~OBA;  //complement 
assign cbi = ~CBI;  //complement 
assign obi = ~OBI;  //complement 
assign qic = ~QIC;  //complement 
assign qid = ~QID;  //complement 
assign qie = ~QIE;  //complement 
assign qif = ~QIF;  //complement 
assign qia = ~QIA;  //complement 
assign QBA = ~qba;  //complement 
assign QBE = ~qbe;  //complement 
assign QMA = ~qma;  //complement 
assign OAS = ~oas;  //complement 
assign qib = ~QIB;  //complement 
assign OAQ = ~oaq;  //complement 
assign OAR = ~oar;  //complement 
assign OAT = ~oat;  //complement 
assign bea = ~BEA;  //complement 
assign bei = ~BEI;  //complement 
assign bfa = ~BFA;  //complement 
assign bfi = ~BFI;  //complement 
assign cca = ~CCA;  //complement 
assign oca = ~OCA;  //complement 
assign cci = ~CCI;  //complement 
assign oci = ~OCI;  //complement 
assign bga = ~BGA;  //complement 
assign bgi = ~BGI;  //complement 
assign bha = ~BHA;  //complement 
assign bhi = ~BHI;  //complement 
assign cda = ~CDA;  //complement 
assign oda = ~ODA;  //complement 
assign cdi = ~CDI;  //complement 
assign odi = ~ODI;  //complement 
assign FAB = EAA; 
assign fab = ~FAB; //complement 
assign FBB = EAB; 
assign fbb = ~FBB;  //complement 
assign FCB = EAC; 
assign fcb = ~FCB;  //complement 
assign FDB = EAD; 
assign fdb = ~FDB;  //complement 
assign FEB = EAE; 
assign feb = ~FEB; //complement 
assign FFB = EAF; 
assign ffb = ~FFB;  //complement 
assign FGB = EAG; 
assign fgb = ~FGB;  //complement 
assign FHB = EAH; 
assign fhb = ~FHB;  //complement 
assign FIB = EAI; 
assign fib = ~FIB; //complement 
assign FJB = EAJ; 
assign fjb = ~FJB;  //complement 
assign FKB = EAK; 
assign fkb = ~FKB;  //complement 
assign FLB = EAL; 
assign flb = ~FLB;  //complement 
assign JAB =  RCA  ; 
assign jab = ~JAB;  //complement  
assign wab = ~WAB;  //complement 
assign JAJ =  HAB & RCI  ; 
assign jaj = ~JAJ;  //complement  
assign kbb = ~KBB;  //complement 
assign lbb = ~LBB;  //complement 
assign JBB =  HAD & RDA  ; 
assign jbb = ~JBB;  //complement  
assign JBJ =  HAF & HBB & RDI  ; 
assign jbj = ~JBJ;  //complement  
assign RAB = ~rab;  //complement 
assign RCB = ~rcb;  //complement 
assign oeb = ~OEB;  //complement 
assign pab = ~PAB;  //complement 
assign DAB =  BAB & QEA  |  BCB & QFA  |  BEB & QGA  |  BGB & QHA  ; 
assign dab = ~DAB;  //complement 
assign aab = ~AAB;  //complement 
assign acb = ~ACB;  //complement 
assign aeb = ~AEB;  //complement 
assign ebb = eab; 
assign EBB = ~ebb; //complement 
assign ebj = eaj; 
assign EBJ = ~ebj;  //complement 
assign RAJ = ~raj;  //complement 
assign RCJ = ~rcj;  //complement 
assign oej = ~OEJ;  //complement 
assign paj = ~PAJ;  //complement 
assign DAJ =  BAJ & QEC  |  BCJ & QFC  |  BEJ & QGC  |  BGJ & QHC  ; 
assign daj = ~DAJ;  //complement 
assign KAB =  AEB & aej  |  aeb & AEJ  |  aeb & aej  |  AEB & AEJ  ; 
assign kab = ~KAB; //complement 
assign KAJ =  AFB & afj  |  afb & AFJ  |  afb & afj  |  AFB & AFJ  ; 
assign kaj = ~KAJ; //complement 
assign aaj = ~AAJ;  //complement 
assign acj = ~ACJ;  //complement 
assign aej = ~AEJ;  //complement 
assign LAB =  PAB & paj  |  pab & PAJ  |  pab & paj  |  PAB & PAJ  ; 
assign lab = ~LAB; //complement 
assign LAJ =  PBB & pbj  |  pbb & PBJ  |  pbb & pbj  |  PBB & PBJ  ; 
assign laj = ~LAJ; //complement 
assign abb = ~ABB;  //complement 
assign adb = ~ADB;  //complement 
assign afb = ~AFB;  //complement 
assign RBB = ~rbb;  //complement 
assign RDB = ~rdb;  //complement 
assign ofb = ~OFB;  //complement 
assign pbb = ~PBB;  //complement 
assign DBB =  BBB & QEE  |  BDB & QFE  |  BFB & QGE  |  BHB & QHE  ; 
assign dbb = ~DBB;  //complement 
assign abj = ~ABJ;  //complement 
assign adj = ~ADJ;  //complement 
assign afj = ~AFJ;  //complement 
assign RBJ = ~rbj;  //complement 
assign RDJ = ~rdj;  //complement 
assign ofj = ~OFJ;  //complement 
assign pbj = ~PBJ;  //complement 
assign DBJ =  BBJ & QEG  |  BDJ & QFG  |  BFJ & QGG  |  BHJ & QHG  ; 
assign dbj = ~DBJ;  //complement 
assign bab = ~BAB;  //complement 
assign baj = ~BAJ;  //complement 
assign bbb = ~BBB;  //complement 
assign bbj = ~BBJ;  //complement 
assign cab = ~CAB;  //complement 
assign oab = ~OAB;  //complement 
assign caj = ~CAJ;  //complement 
assign oaj = ~OAJ;  //complement 
assign eab = ~EAB;  //complement 
assign eaj = ~EAJ;  //complement 
assign tci = qje & qjc ; 
assign TCI = ~tci ; //complement 
assign tcj = qje & qjc ; 
assign TCJ = ~tcj ;  //complement 
assign tck = qjf & qjd ; 
assign TCK = ~tck ;  //complement 
assign tcl = qjf & qjd; 
assign TCL = ~tcl; 
assign tcg = QJB; 
assign TCG = ~tcg; //complement 
assign tch = QJB; 
assign TCH = ~tch;  //complement 
assign bcb = ~BCB;  //complement 
assign bcj = ~BCJ;  //complement 
assign bdb = ~BDB;  //complement 
assign bdj = ~BDJ;  //complement 
assign cbb = ~CBB;  //complement 
assign obb = ~OBB;  //complement 
assign cbj = ~CBJ;  //complement 
assign obj = ~OBJ;  //complement 
assign qjc = ~QJC;  //complement 
assign qjd = ~QJD;  //complement 
assign qje = ~QJE;  //complement 
assign qjf = ~QJF;  //complement 
assign qja = ~QJA;  //complement 
assign QBB = ~qbb;  //complement 
assign QBF = ~qbf;  //complement 
assign QMB = ~qmb;  //complement 
assign OBS = ~obs;  //complement 
assign qjb = ~QJB;  //complement 
assign OBQ = ~obq;  //complement 
assign OBR = ~obr;  //complement 
assign OBT = ~obt;  //complement 
assign beb = ~BEB;  //complement 
assign bej = ~BEJ;  //complement 
assign bfb = ~BFB;  //complement 
assign bfj = ~BFJ;  //complement 
assign ccb = ~CCB;  //complement 
assign ocb = ~OCB;  //complement 
assign ccj = ~CCJ;  //complement 
assign ocj = ~OCJ;  //complement 
assign bgb = ~BGB;  //complement 
assign bgj = ~BGJ;  //complement 
assign bhb = ~BHB;  //complement 
assign bhj = ~BHJ;  //complement 
assign cdb = ~CDB;  //complement 
assign odb = ~ODB;  //complement 
assign cdj = ~CDJ;  //complement 
assign odj = ~ODJ;  //complement 
assign FAC = EAA; 
assign fac = ~FAC; //complement 
assign FBC = EAB; 
assign fbc = ~FBC;  //complement 
assign FCC = EAC; 
assign fcc = ~FCC;  //complement 
assign FDC = EAD; 
assign fdc = ~FDC;  //complement 
assign FEC = EAE; 
assign fec = ~FEC; //complement 
assign FFC = EAF; 
assign ffc = ~FFC;  //complement 
assign FGC = EAG; 
assign fgc = ~FGC;  //complement 
assign FHC = EAH; 
assign fhc = ~FHC;  //complement 
assign FIC = EAI; 
assign fic = ~FIC; //complement 
assign FJC = EAJ; 
assign fjc = ~FJC;  //complement 
assign FKC = EAK; 
assign fkc = ~FKC;  //complement 
assign FLC = EAL; 
assign flc = ~FLC;  //complement 
assign JAC =  RCA & RCB  ; 
assign jac = ~JAC;  //complement  
assign wac = ~WAC;  //complement 
assign JAK =  HAB & RCI & RCJ  ; 
assign jak = ~JAK;  //complement  
assign kbc = ~KBC;  //complement 
assign lbc = ~LBC;  //complement 
assign JBC =  HAD & RDA & RDB  ; 
assign jbc = ~JBC;  //complement  
assign HAD = ~had;  //complement 
assign HAE = ~hae;  //complement 
assign JBK =  HAF & HBB & RDI & RDJ  ; 
assign jbk = ~JBK;  //complement  
assign RAC = ~rac;  //complement 
assign RCC = ~rcc;  //complement 
assign oec = ~OEC;  //complement 
assign pac = ~PAC;  //complement 
assign DAC =  BAC & QEA  |  BCC & QFA  |  BEC & QGA  |  BGC & QHA  ; 
assign dac = ~DAC;  //complement 
assign aac = ~AAC;  //complement 
assign acc = ~ACC;  //complement 
assign aec = ~AEC;  //complement 
assign ebc = eac; 
assign EBC = ~ebc; //complement 
assign ebk = eak; 
assign EBK = ~ebk;  //complement 
assign RAK = ~rak;  //complement 
assign RCK = ~rck;  //complement 
assign oek = ~OEK;  //complement 
assign pak = ~PAK;  //complement 
assign DAK =  BAK & QEC  |  BCK & QFC  |  BEK & QGC  |  BGK & QHC  ; 
assign dak = ~DAK;  //complement 
assign KAC =  AEC & aek  |  aec & AEK  |  aec & aek  |  AEC & AEK  ; 
assign kac = ~KAC; //complement 
assign KAK =  AFC & afk  |  afc & AFK  |  afc & afk  |  AFC & AFK  ; 
assign kak = ~KAK; //complement 
assign aak = ~AAK;  //complement 
assign ack = ~ACK;  //complement 
assign aek = ~AEK;  //complement 
assign LAC =  PAC & pak  |  pac & PAK  |  pac & pak  |  PAC & PAK  ; 
assign lac = ~LAC; //complement 
assign LAK =  PBC & pbk  |  pbc & PBK  |  pbc & pbk  |  PBC & PBK  ; 
assign lak = ~LAK; //complement 
assign abc = ~ABC;  //complement 
assign adc = ~ADC;  //complement 
assign afc = ~AFC;  //complement 
assign RBC = ~rbc;  //complement 
assign RDC = ~rdc;  //complement 
assign ofc = ~OFC;  //complement 
assign pbc = ~PBC;  //complement 
assign DBC =  BBC & QEE  |  BDC & QFE  |  BFC & QGE  |  BHC & QHE  ; 
assign dbc = ~DBC;  //complement 
assign abk = ~ABK;  //complement 
assign adk = ~ADK;  //complement 
assign afk = ~AFK;  //complement 
assign RBK = ~rbk;  //complement 
assign RDK = ~rdk;  //complement 
assign ofk = ~OFK;  //complement 
assign pbk = ~PBK;  //complement 
assign DBK =  BBK & QEG  |  BDK & QFG  |  BFK & QGG  |  BHK & QHG  ; 
assign dbk = ~DBK;  //complement 
assign bac = ~BAC;  //complement 
assign bak = ~BAK;  //complement 
assign bbc = ~BBC;  //complement 
assign bbk = ~BBK;  //complement 
assign cac = ~CAC;  //complement 
assign oac = ~OAC;  //complement 
assign cak = ~CAK;  //complement 
assign oak = ~OAK;  //complement 
assign eac = ~EAC;  //complement 
assign eak = ~EAK;  //complement 
assign bcc = ~BCC;  //complement 
assign bck = ~BCK;  //complement 
assign bdc = ~BDC;  //complement 
assign bdk = ~BDK;  //complement 
assign cbc = ~CBC;  //complement 
assign obc = ~OBC;  //complement 
assign cbk = ~CBK;  //complement 
assign obk = ~OBK;  //complement 
assign qkc = ~QKC;  //complement 
assign qkd = ~QKD;  //complement 
assign qke = ~QKE;  //complement 
assign qkf = ~QKF;  //complement 
assign qka = ~QKA;  //complement 
assign QBC = ~qbc;  //complement 
assign QBG = ~qbg;  //complement 
assign QMC = ~qmc;  //complement 
assign OCS = ~ocs;  //complement 
assign qkb = ~QKB;  //complement 
assign OCQ = ~ocq;  //complement 
assign OCR = ~ocr;  //complement 
assign OCT = ~oct;  //complement 
assign bec = ~BEC;  //complement 
assign bek = ~BEK;  //complement 
assign bfc = ~BFC;  //complement 
assign bfk = ~BFK;  //complement 
assign ccc = ~CCC;  //complement 
assign occ = ~OCC;  //complement 
assign cck = ~CCK;  //complement 
assign ock = ~OCK;  //complement 
assign tco = qke & qkc ; 
assign TCO = ~tco ; //complement 
assign tcp = qke & qkc ; 
assign TCP = ~tcp ;  //complement 
assign tcq = qkf & qkd ; 
assign TCQ = ~tcq ;  //complement 
assign tcr = qkf & qkd; 
assign TCR = ~tcr; 
assign tcm = QKB; 
assign TCM = ~tcm; //complement 
assign tcn = QKB; 
assign TCN = ~tcn;  //complement 
assign bgc = ~BGC;  //complement 
assign bgk = ~BGK;  //complement 
assign bhc = ~BHC;  //complement 
assign bhk = ~BHK;  //complement 
assign cdc = ~CDC;  //complement 
assign odc = ~ODC;  //complement 
assign cdk = ~CDK;  //complement 
assign odk = ~ODK;  //complement 
assign FAD = EAA; 
assign fad = ~FAD; //complement 
assign FBD = EAB; 
assign fbd = ~FBD;  //complement 
assign FCD = EAC; 
assign fcd = ~FCD;  //complement 
assign FDD = EAD; 
assign fdd = ~FDD;  //complement 
assign FED = EAE; 
assign fed = ~FED; //complement 
assign FFD = EAF; 
assign ffd = ~FFD;  //complement 
assign FGD = EAG; 
assign fgd = ~FGD;  //complement 
assign FHD = EAH; 
assign fhd = ~FHD;  //complement 
assign FID = EAI; 
assign fid = ~FID; //complement 
assign FJD = EAJ; 
assign fjd = ~FJD;  //complement 
assign FKD = EAK; 
assign fkd = ~FKD;  //complement 
assign FLD = EAL; 
assign fld = ~FLD;  //complement 
assign JAQ =  rca & RCB & RCC & RCD  ; 
assign jaq = ~JAQ;  //complement  
assign JAD =  RCA & RCB & RCC  ; 
assign jad = ~JAD;  //complement 
assign wad = ~WAD;  //complement 
assign kda = ~KDA;  //complement 
assign JAS =  RCI & RCJ & RCK & RCL  ; 
assign jas = ~JAS;  //complement  
assign JAL =  HAB & RCI & RCJ & RCK  ; 
assign jal = ~JAL;  //complement 
assign KCB =  KBD & kbe  |  kbd & KBE  |  kbd & kbe  |  KBD & KBE  ; 
assign kcb = ~KCB; //complement 
assign KCA =  KBA & kbb & kbc  |  kba & KBB & kbc  |  kba & kbb & KBC  |  KBA & KBB & KBC  ; 
assign kca = ~KCA; //complement 
assign kbd = ~KBD;  //complement 
assign LCA =  LBA & lbb & lbc  |  lba & LBB & lbc  |  lba & lbb & LBC  |  LBA & LBB & LBC  ; 
assign lca = ~LCA; //complement 
assign lbd = ~LBD;  //complement 
assign JBQ =  RDA & RDB & RDC & RDD  ; 
assign jbq = ~JBQ;  //complement  
assign JBD =  HAD & RDA & RDB & RDC  ; 
assign jbd = ~JBD;  //complement 
assign HAF = ~haf;  //complement 
assign HAG = ~hag;  //complement 
assign JBL =  HAF & HBB & RDI & RDJ & RDK  ; 
assign jbl = ~JBL;  //complement  
assign JBS =  RDI & RDJ & RDK & RDL  ; 
assign jbs = ~JBS;  //complement 
assign RAD = ~rad;  //complement 
assign RCD = ~rcd;  //complement 
assign pad = ~PAD;  //complement 
assign oed = ~OED;  //complement 
assign DAD =  BAD & QEA  |  BCD & QFA  |  BED & QGA  |  BGD & QHA  ; 
assign dad = ~DAD;  //complement 
assign aad = ~AAD;  //complement 
assign acd = ~ACD;  //complement 
assign aed = ~AED;  //complement 
assign qea = ~QEA;  //complement 
assign qfa = ~QFA;  //complement 
assign qga = ~QGA;  //complement 
assign qha = ~QHA;  //complement 
assign RAL = ~ral;  //complement 
assign RCL = ~rcl;  //complement 
assign pal = ~PAL;  //complement 
assign oel = ~OEL;  //complement 
assign DAL =  BAL & QEC  |  BCL & QFC  |  BEL & QGC  |  BGL & QHC  ; 
assign dal = ~DAL;  //complement 
assign KAD =  AED & ael  |  aed & AEL  |  aed & ael  |  AED & AEL  ; 
assign kad = ~KAD; //complement 
assign KAL =  AFD & afl  |  afd & AFL  |  afd & afl  |  AFD & AFL  ; 
assign kal = ~KAL; //complement 
assign aal = ~AAL;  //complement 
assign acl = ~ACL;  //complement 
assign ael = ~AEL;  //complement 
assign qec = ~QEC;  //complement 
assign qfc = ~QFC;  //complement 
assign qgc = ~QGC;  //complement 
assign qhc = ~QHC;  //complement 
assign LAD =  PAD & pal  |  pad & PAL  |  pad & pal  |  PAD & PAL  ; 
assign lad = ~LAD; //complement 
assign LAL =  PBD & pbl  |  pbd & PBL  |  pbd & pbl  |  PBD & PBL  ; 
assign lal = ~LAL; //complement 
assign abd = ~ABD;  //complement 
assign add = ~ADD;  //complement 
assign afd = ~AFD;  //complement 
assign QEE = ~qee;  //complement 
assign QFE = ~qfe;  //complement 
assign QGE = ~qge;  //complement 
assign QHE = ~qhe;  //complement 
assign RBD = ~rbd;  //complement 
assign RDD = ~rdd;  //complement 
assign ofd = ~OFD;  //complement 
assign pbd = ~PBD;  //complement 
assign DBD =  BBD & QEE  |  BDD & QFE  |  BFD & QGE  |  BHD & QHE  ; 
assign dbd = ~DBD;  //complement 
assign abl = ~ABL;  //complement 
assign adl = ~ADL;  //complement 
assign afl = ~AFL;  //complement 
assign QEG = ~qeg;  //complement 
assign QFG = ~qfg;  //complement 
assign QGG = ~qgg;  //complement 
assign QHG = ~qhg;  //complement 
assign RBL = ~rbl;  //complement 
assign RDL = ~rdl;  //complement 
assign ofl = ~OFL;  //complement 
assign pbl = ~PBL;  //complement 
assign DBL =  BBL & QEG  |  BDL & QFG  |  BFL & QGG  |  BHL & QHG  ; 
assign dbl = ~DBL;  //complement 
assign bad = ~BAD;  //complement 
assign bal = ~BAL;  //complement 
assign bbd = ~BBD;  //complement 
assign bbl = ~BBL;  //complement 
assign cad = ~CAD;  //complement 
assign oad = ~OAD;  //complement 
assign cal = ~CAL;  //complement 
assign oal = ~OAL;  //complement 
assign ead = ~EAD;  //complement 
assign eal = ~EAL;  //complement 
assign ebd = ead; 
assign EBD = ~ebd; //complement 
assign ebl = eal; 
assign EBL = ~ebl;  //complement 
assign bcd = ~BCD;  //complement 
assign bcl = ~BCL;  //complement 
assign bdd = ~BDD;  //complement 
assign bdl = ~BDL;  //complement 
assign cbd = ~CBD;  //complement 
assign obd = ~OBD;  //complement 
assign cbl = ~CBL;  //complement 
assign obl = ~OBL;  //complement 
assign qlc = ~QLC;  //complement 
assign qld = ~QLD;  //complement 
assign qle = ~QLE;  //complement 
assign qlf = ~QLF;  //complement 
assign qla = ~QLA;  //complement 
assign QBD = ~qbd;  //complement 
assign QBH = ~qbh;  //complement 
assign QMD = ~qmd;  //complement 
assign ODS = ~ods;  //complement 
assign qlb = ~QLB;  //complement 
assign ODQ = ~odq;  //complement 
assign ODR = ~odr;  //complement 
assign ODT = ~odt;  //complement 
assign bed = ~BED;  //complement 
assign bel = ~BEL;  //complement 
assign bfd = ~BFD;  //complement 
assign bfl = ~BFL;  //complement 
assign ccd = ~CCD;  //complement 
assign ocd = ~OCD;  //complement 
assign ccl = ~CCL;  //complement 
assign ocl = ~OCL;  //complement 
assign tcu = qle & qlc ; 
assign TCU = ~tcu ; //complement 
assign tcv = qle & qlc ; 
assign TCV = ~tcv ;  //complement 
assign tcw = qlf & qld ; 
assign TCW = ~tcw ;  //complement 
assign tcx = qlf & qld; 
assign TCX = ~tcx; 
assign tcs = QLB; 
assign TCS = ~tcs; //complement 
assign tct = QLB; 
assign TCT = ~tct;  //complement 
assign bgd = ~BGD;  //complement 
assign bgl = ~BGL;  //complement 
assign bhd = ~BHD;  //complement 
assign bhl = ~BHL;  //complement 
assign cdd = ~CDD;  //complement 
assign odd = ~ODD;  //complement 
assign cdl = ~CDL;  //complement 
assign odl = ~ODL;  //complement 
assign FAE = EAA; 
assign fae = ~FAE; //complement 
assign FBE = EAB; 
assign fbe = ~FBE;  //complement 
assign FCE = EAC; 
assign fce = ~FCE;  //complement 
assign FDE = EAD; 
assign fde = ~FDE;  //complement 
assign FEE = EAE; 
assign fee = ~FEE; //complement 
assign FFE = EAF; 
assign ffe = ~FFE;  //complement 
assign FGE = EAG; 
assign fge = ~FGE;  //complement 
assign FHE = EAH; 
assign fhe = ~FHE;  //complement 
assign FIE = EAI; 
assign fie = ~FIE; //complement 
assign FJE = EAJ; 
assign fje = ~FJE;  //complement 
assign FKE = EAK; 
assign fke = ~FKE;  //complement 
assign FLE = EAL; 
assign fle = ~FLE;  //complement 
assign JAE =  HAA  ; 
assign jae = ~JAE;  //complement  
assign wae = ~WAE;  //complement 
assign haa = ~HAA;  //complement 
assign JAM =  HAC  ; 
assign jam = ~JAM;  //complement  
assign LCB =  LBD & lbe  |  lbd & LBE  |  lbd & lbe  |  LBD & LBE  ; 
assign lcb = ~LCB; //complement 
assign KCC =  KBF & kbg & kbh  |  kbf & KBG & kbh  |  kbf & kbg & KBH  |  KBF & KBG & KBH  ; 
assign kcc = ~KCC; //complement 
assign kbe = ~KBE;  //complement 
assign lda = ~LDA;  //complement 
assign LCC =  LBF & lbg & lbh  |  lbf & LBG & lbh  |  lbf & lbg & LBH  |  LBF & LBG & LBH  ; 
assign lcc = ~LCC; //complement 
assign lbe = ~LBE;  //complement 
assign JBE =  HAE & HBA  ; 
assign jbe = ~JBE;  //complement  
assign hba = ~HBA;  //complement 
assign JBM =  HAG & HBC  ; 
assign jbm = ~JBM;  //complement  
assign RAE = ~rae;  //complement 
assign RCE = ~rce;  //complement 
assign oee = ~OEE;  //complement 
assign pae = ~PAE;  //complement 
assign DAE =  BAE & QEB  |  BCE & QFB  |  BEE & QGB  |  BGE & QHB  ; 
assign dae = ~DAE;  //complement 
assign aae = ~AAE;  //complement 
assign ace = ~ACE;  //complement 
assign aee = ~AEE;  //complement 
assign qeb = ~QEB;  //complement 
assign qfb = ~QFB;  //complement 
assign qgb = ~QGB;  //complement 
assign qhb = ~QHB;  //complement 
assign RAM = ~ram;  //complement 
assign RCM = ~rcm;  //complement 
assign oem = ~OEM;  //complement 
assign pam = ~PAM;  //complement 
assign DAM =  BAM & QED  |  BCM & QFD  |  BEM & QGD  |  BGM & QHD  ; 
assign dam = ~DAM;  //complement 
assign KAE =  AEE & aem  |  aee & AEM  |  aee & aem  |  AEE & AEM  ; 
assign kae = ~KAE; //complement 
assign KAM =  AFE & afm  |  afe & AFM  |  afe & afm  |  AFE & AFM  ; 
assign kam = ~KAM; //complement 
assign aam = ~AAM;  //complement 
assign acm = ~ACM;  //complement 
assign aem = ~AEM;  //complement 
assign qed = ~QED;  //complement 
assign qfd = ~QFD;  //complement 
assign qgd = ~QGD;  //complement 
assign qhd = ~QHD;  //complement 
assign LAE =  PAE & pam  |  pae & PAM  |  pae & pam  |  PAE & PAM  ; 
assign lae = ~LAE; //complement 
assign LAM =  PBE & pbm  |  pbe & PBM  |  pbe & pbm  |  PBE & PBM  ; 
assign lam = ~LAM; //complement 
assign abe = ~ABE;  //complement 
assign ade = ~ADE;  //complement 
assign afe = ~AFE;  //complement 
assign QEF = ~qef;  //complement 
assign QFF = ~qff;  //complement 
assign QGF = ~qgf;  //complement 
assign QHF = ~qhf;  //complement 
assign RBE = ~rbe;  //complement 
assign RDE = ~rde;  //complement 
assign ofe = ~OFE;  //complement 
assign pbe = ~PBE;  //complement 
assign DBE =  BBE & QEF  |  BDE & QFF  |  BFE & QGF  |  BHE & QHF  ; 
assign dbe = ~DBE;  //complement 
assign abm = ~ABM;  //complement 
assign adm = ~ADM;  //complement 
assign afm = ~AFM;  //complement 
assign QGH = ~qgh;  //complement 
assign QHH = ~qhh;  //complement 
assign QEH = ~qeh;  //complement 
assign QFH = ~qfh;  //complement 
assign RBM = ~rbm;  //complement 
assign RDM = ~rdm;  //complement 
assign ofm = ~OFM;  //complement 
assign pbm = ~PBM;  //complement 
assign DBM =  BBM & QEH  |  BDM & QFH  |  BFM & QGH  |  BHM & QHH  ; 
assign dbm = ~DBM;  //complement 
assign bae = ~BAE;  //complement 
assign bam = ~BAM;  //complement 
assign bbe = ~BBE;  //complement 
assign bbm = ~BBM;  //complement 
assign cae = ~CAE;  //complement 
assign oae = ~OAE;  //complement 
assign cam = ~CAM;  //complement 
assign oam = ~OAM;  //complement 
assign eae = ~EAE;  //complement 
assign ebe = eae; 
assign EBE = ~ebe; //complement 
assign bce = ~BCE;  //complement 
assign bcm = ~BCM;  //complement 
assign bde = ~BDE;  //complement 
assign bdm = ~BDM;  //complement 
assign cbe = ~CBE;  //complement 
assign obe = ~OBE;  //complement 
assign cbm = ~CBM;  //complement 
assign obm = ~OBM;  //complement 
assign JCA =  QAE & qab & qaa  ; 
assign jca = ~JCA;  //complement 
assign JCB =  QAE & qab & QAA  ; 
assign jcb = ~JCB;  //complement 
assign JCE =  QAE & QAA  ; 
assign jce = ~JCE;  //complement 
assign JCC =  QAE & QAB & qaa  ; 
assign jcc = ~JCC;  //complement 
assign JCD =  QAE & QAB & QAA  ; 
assign jcd = ~JCD;  //complement 
assign qaa = ~QAA;  //complement 
assign qab = ~QAB;  //complement 
assign qae = ~QAE;  //complement 
assign bee = ~BEE;  //complement 
assign bem = ~BEM;  //complement 
assign bfe = ~BFE;  //complement 
assign bfm = ~BFM;  //complement 
assign cce = ~CCE;  //complement 
assign oce = ~OCE;  //complement 
assign ccm = ~CCM;  //complement 
assign ocm = ~OCM;  //complement 
assign bge = ~BGE;  //complement 
assign bgm = ~BGM;  //complement 
assign bhe = ~BHE;  //complement 
assign bhm = ~BHM;  //complement 
assign cde = ~CDE;  //complement 
assign ode = ~ODE;  //complement 
assign cdm = ~CDM;  //complement 
assign odm = ~ODM;  //complement 
assign FAF = EAA; 
assign faf = ~FAF; //complement 
assign FBF = EAB; 
assign fbf = ~FBF;  //complement 
assign FCF = EAC; 
assign fcf = ~FCF;  //complement 
assign FDF = EAD; 
assign fdf = ~FDF;  //complement 
assign FEF = EAE; 
assign fef = ~FEF; //complement 
assign FFF = EAF; 
assign fff = ~FFF;  //complement 
assign FGF = EAG; 
assign fgf = ~FGF;  //complement 
assign FHF = EAH; 
assign fhf = ~FHF;  //complement 
assign FIF = EAI; 
assign fif = ~FIF; //complement 
assign FJF = EAJ; 
assign fjf = ~FJF;  //complement 
assign FKF = EAK; 
assign fkf = ~FKF;  //complement 
assign FLF = EAL; 
assign flf = ~FLF;  //complement 
assign JAF =  HAA & RCE  ; 
assign jaf = ~JAF;  //complement  
assign waf = ~WAF;  //complement 
assign qca = ~QCA;  //complement 
assign qcb = ~QCB;  //complement 
assign hab = ~HAB;  //complement 
assign QCC = ~qcc;  //complement 
assign QCD = ~qcd;  //complement 
assign QCE = ~qce;  //complement 
assign QCF = ~qcf;  //complement 
assign JAN =  HAC & RCM  ; 
assign jan = ~JAN;  //complement  
assign kbf = ~KBF;  //complement 
assign lbf = ~LBF;  //complement 
assign JBF =  HAE & HBA & RDE  ; 
assign jbf = ~JBF;  //complement  
assign qcg = ~QCG;  //complement 
assign qch = ~QCH;  //complement 
assign hbb = ~HBB;  //complement 
assign pbq = ~PBQ;  //complement 
assign LEA =  LDA & pbq  |  lda & PBQ  ; 
assign lea = ~LEA; //complement 
assign JBN =  HAG & HBC & RDM  ; 
assign jbn = ~JBN;  //complement  
assign RAF = ~raf;  //complement 
assign RCF = ~rcf;  //complement 
assign paf = ~PAF;  //complement 
assign oef = ~OEF;  //complement 
assign DAF =  BAF & QEB  |  BCF & QFB  |  BEF & QGB  |  BGF & QHB  ; 
assign daf = ~DAF;  //complement 
assign QDA = ~qda;  //complement 
assign QDB = ~qdb;  //complement 
assign aaf = ~AAF;  //complement 
assign acf = ~ACF;  //complement 
assign aef = ~AEF;  //complement 
assign ebf = aea; 
assign EBF = ~ebf; //complement 
assign TDI = QAG; 
assign tdi = ~TDI;  //complement 
assign TDJ = QAG; 
assign tdj = ~TDJ;  //complement 
assign RAN = ~ran;  //complement 
assign RCN = ~rcn;  //complement 
assign pan = ~PAN;  //complement 
assign oen = ~OEN;  //complement 
assign DAN =  BAN & QED  |  BCN & QFD  |  BEN & QGD  |  BGN & QHD  ; 
assign dan = ~DAN;  //complement 
assign KAF =  AEF & aen  |  aef & AEN  |  aef & aen  |  AEF & AEN  ; 
assign kaf = ~KAF; //complement 
assign KAN =  AFF & afn  |  aff & AFN  |  aff & afn  |  AFF & AFN  ; 
assign kan = ~KAN; //complement 
assign aan = ~AAN;  //complement 
assign acn = ~ACN;  //complement 
assign aen = ~AEN;  //complement 
assign qag = ~QAG;  //complement 
assign qah = ~QAH;  //complement 
assign LAF =  PAF & pan  |  paf & PAN  |  paf & pan  |  PAF & PAN  ; 
assign laf = ~LAF; //complement 
assign LAN =  PBF & pbn  |  pbf & PBN  |  pbf & pbn  |  PBF & PBN  ; 
assign lan = ~LAN; //complement 
assign abf = ~ABF;  //complement 
assign adf = ~ADF;  //complement 
assign aff = ~AFF;  //complement 
assign RBF = ~rbf;  //complement 
assign RDF = ~rdf;  //complement 
assign pbf = ~PBF;  //complement 
assign off = ~OFF;  //complement 
assign DBF =  BBF & QEF  |  BDF & QFF  |  BFF & QGF  |  BHF & QHF  ; 
assign dbf = ~DBF;  //complement 
assign QDC = ~qdc;  //complement 
assign QDD = ~qdd;  //complement 
assign abn = ~ABN;  //complement 
assign adn = ~ADN;  //complement 
assign afn = ~AFN;  //complement 
assign tdk = qag; 
assign TDK = ~tdk; //complement 
assign tdl = qag; 
assign TDL = ~tdl;  //complement 
assign RBN = ~rbn;  //complement 
assign RDN = ~rdn;  //complement 
assign pbn = ~PBN;  //complement 
assign ofn = ~OFN;  //complement 
assign DBN =  BBN & QEH  |  BDN & QFH  |  BFN & QGH  |  BHN & QHH  ; 
assign dbn = ~DBN;  //complement 
assign baf = ~BAF;  //complement 
assign ban = ~BAN;  //complement 
assign bbf = ~BBF;  //complement 
assign bbn = ~BBN;  //complement 
assign caf = ~CAF;  //complement 
assign oaf = ~OAF;  //complement 
assign can = ~CAN;  //complement 
assign oan = ~OAN;  //complement 
assign eaf = ~EAF;  //complement 
assign TEA = qai & qaj ; 
assign tea = ~TEA ; //complement 
assign teb = qai & qai ; 
assign TEB = ~teb ;  //complement 
assign tec = qaj; 
assign TEC = ~tec;  //complement 
assign bcf = ~BCF;  //complement 
assign bcn = ~BCN;  //complement 
assign bdf = ~BDF;  //complement 
assign bdn = ~BDN;  //complement 
assign cbf = ~CBF;  //complement 
assign obf = ~OBF;  //complement 
assign cbn = ~CBN;  //complement 
assign obn = ~OBN;  //complement 
assign qai = ~QAI;  //complement 
assign qaj = ~QAJ;  //complement 
assign oha = ~OHA;  //complement 
assign qak = ~QAK;  //complement 
assign bef = ~BEF;  //complement 
assign ben = ~BEN;  //complement 
assign bff = ~BFF;  //complement 
assign bfn = ~BFN;  //complement 
assign ccf = ~CCF;  //complement 
assign ocf = ~OCF;  //complement 
assign ccn = ~CCN;  //complement 
assign ocn = ~OCN;  //complement 
assign bgf = ~BGF;  //complement 
assign bgn = ~BGN;  //complement 
assign bhf = ~BHF;  //complement 
assign bhn = ~BHN;  //complement 
assign cdf = ~CDF;  //complement 
assign odf = ~ODF;  //complement 
assign cdn = ~CDN;  //complement 
assign odn = ~ODN;  //complement 
assign FAG = EAA; 
assign fag = ~FAG; //complement 
assign FBG = EAB; 
assign fbg = ~FBG;  //complement 
assign FCG = EAC; 
assign fcg = ~FCG;  //complement 
assign FDG = EAD; 
assign fdg = ~FDG;  //complement 
assign FEG = EAE; 
assign feg = ~FEG; //complement 
assign FFG = EAF; 
assign ffg = ~FFG;  //complement 
assign FGG = EAG; 
assign fgg = ~FGG;  //complement 
assign FHG = EAH; 
assign fhg = ~FHG;  //complement 
assign FIG = EAI; 
assign fig = ~FIG; //complement 
assign FJG = EAJ; 
assign fjg = ~FJG;  //complement 
assign FKG = EAK; 
assign fkg = ~FKG;  //complement 
assign FLG = EAL; 
assign flg = ~FLG;  //complement 
assign JAG =  HAA & RCE & RCF  ; 
assign jag = ~JAG;  //complement  
assign wag = ~WAG;  //complement 
assign hac = ~HAC;  //complement 
assign JAO =  HAC & RCM & RCN  ; 
assign jao = ~JAO;  //complement  
assign kbg = ~KBG;  //complement 
assign lbg = ~LBG;  //complement 
assign JBG =  HAE & HBA & RDE & RDF  ; 
assign jbg = ~JBG;  //complement  
assign hbc = ~HBC;  //complement 
assign JBO =  HAG & HBC & RDM & RDN  ; 
assign jbo = ~JBO;  //complement  
assign RAG = ~rag;  //complement 
assign RCG = ~rcg;  //complement 
assign oeg = ~OEG;  //complement 
assign pag = ~PAG;  //complement 
assign DAG =  BAG & QEB  |  BCG & QFB  |  BEG & QGB  |  BGG & QHB  ; 
assign dag = ~DAG;  //complement 
assign aag = ~AAG;  //complement 
assign acg = ~ACG;  //complement 
assign aeg = ~AEG;  //complement 
assign ebg = eag; 
assign EBG = ~ebg; //complement 
assign TDE = QAF; 
assign tde = ~TDE;  //complement 
assign TDF = QAF; 
assign tdf = ~TDF;  //complement 
assign RAO = ~rao;  //complement 
assign RCO = ~rco;  //complement 
assign oeo = ~OEO;  //complement 
assign pao = ~PAO;  //complement 
assign DAO =  BAO & QED  |  BCO & QFD  |  BEO & QGD  |  BGO & QHD  ; 
assign dao = ~DAO;  //complement 
assign KAG =  AEG & aeo  |  aeg & AEO  |  aeg & aeo  |  AEG & AEO  ; 
assign kag = ~KAG; //complement 
assign KAO =  AFG & afo  |  afg & AFO  |  afg & afo  |  AFG & AFO  ; 
assign kao = ~KAO; //complement 
assign aao = ~AAO;  //complement 
assign aco = ~ACO;  //complement 
assign aeo = ~AEO;  //complement 
assign qaf = ~QAF;  //complement 
assign LAG =  PAG & pao  |  pag & PAO  |  pag & pao  |  PAG & PAO  ; 
assign lag = ~LAG; //complement 
assign LAO =  PBG & pbo  |  pbg & PBO  |  pbg & pbo  |  PBG & PBO  ; 
assign lao = ~LAO; //complement 
assign abg = ~ABG;  //complement 
assign adg = ~ADG;  //complement 
assign afg = ~AFG;  //complement 
assign RBG = ~rbg;  //complement 
assign RDG = ~rdg;  //complement 
assign ofg = ~OFG;  //complement 
assign pbg = ~PBG;  //complement 
assign DBG =  BBG & QEF  |  BDG & QFF  |  BFG & QGF  |  BHG & QHF  ; 
assign dbg = ~DBG;  //complement 
assign abo = ~ABO;  //complement 
assign ado = ~ADO;  //complement 
assign afo = ~AFO;  //complement 
assign tdg = qaf; 
assign TDG = ~tdg; //complement 
assign tdh = qaf; 
assign TDH = ~tdh;  //complement 
assign RBO = ~rbo;  //complement 
assign RDO = ~rdo;  //complement 
assign ofo = ~OFO;  //complement 
assign pbo = ~PBO;  //complement 
assign DBO =  BBO & QEH  |  BDO & QFH  |  BFO & QGH  |  BHO & QHH  ; 
assign dbo = ~DBO;  //complement 
assign bag = ~BAG;  //complement 
assign bao = ~BAO;  //complement 
assign bbg = ~BBG;  //complement 
assign bbo = ~BBO;  //complement 
assign cag = ~CAG;  //complement 
assign oag = ~OAG;  //complement 
assign cao = ~CAO;  //complement 
assign oao = ~OAO;  //complement 
assign eag = ~EAG;  //complement 
assign tba = ~TBA;  //complement 
assign tbb = ~TBB;  //complement 
assign tbc = ~TBC;  //complement 
assign tbd = ~TBD;  //complement 
assign bcg = ~BCG;  //complement 
assign bco = ~BCO;  //complement 
assign bdg = ~BDG;  //complement 
assign bdo = ~BDO;  //complement 
assign cbg = ~CBG;  //complement 
assign obg = ~OBG;  //complement 
assign cbo = ~CBO;  //complement 
assign obo = ~OBO;  //complement 
assign qih = ~QIH;  //complement 
assign qjh = ~QJH;  //complement 
assign oga = ~OGA;  //complement 
assign qig = ~QIG;  //complement 
assign ogb = ~OGB;  //complement 
assign qjg = ~QJG;  //complement 
assign beg = ~BEG;  //complement 
assign beo = ~BEO;  //complement 
assign bfg = ~BFG;  //complement 
assign bfo = ~BFO;  //complement 
assign ccg = ~CCG;  //complement 
assign ocg = ~OCG;  //complement 
assign cco = ~CCO;  //complement 
assign oco = ~OCO;  //complement 
assign bgg = ~BGG;  //complement 
assign bgo = ~BGO;  //complement 
assign bhg = ~BHG;  //complement 
assign bho = ~BHO;  //complement 
assign cdg = ~CDG;  //complement 
assign odg = ~ODG;  //complement 
assign cdo = ~CDO;  //complement 
assign odo = ~ODO;  //complement 
assign FAH = EAA; 
assign fah = ~FAH; //complement 
assign FBH = EAB; 
assign fbh = ~FBH;  //complement 
assign FCH = EAC; 
assign fch = ~FCH;  //complement 
assign FDH = EAD; 
assign fdh = ~FDH;  //complement 
assign FEH = EAE; 
assign feh = ~FEH; //complement 
assign FFH = EAF; 
assign ffh = ~FFH;  //complement 
assign FGH = EAG; 
assign fgh = ~FGH;  //complement 
assign FHH = EAH; 
assign fhh = ~FHH;  //complement 
assign FIH = EAI; 
assign fih = ~FIH; //complement 
assign FJH = EAJ; 
assign fjh = ~FJH;  //complement 
assign FKH = EAK; 
assign fkh = ~FKH;  //complement 
assign FLH = EAL; 
assign flh = ~FLH;  //complement 
assign JAR =  RCE & RCF & RCG & RCH  ; 
assign jar = ~JAR;  //complement  
assign JAH =  HAA & RCE & RCF & RCG  ; 
assign jah = ~JAH;  //complement 
assign wah = ~WAH;  //complement 
assign JAT =  RCM & RCN & RCO & RCP  ; 
assign jat = ~JAT;  //complement  
assign JAP =  HAC & RCM & RCN & RCO  ; 
assign jap = ~JAP;  //complement 
assign kbh = ~KBH;  //complement 
assign lbh = ~LBH;  //complement 
assign JBH =  HAE & HBA & RDE & RDF & RDG  ; 
assign jbh = ~JBH;  //complement  
assign JBR =  RDE & RDF & RDG & RDH  ; 
assign jbr = ~JBR;  //complement 
assign JBP =  HAG & HBC & RDM & RDN & RDO  ; 
assign jbp = ~JBP;  //complement  
assign RAH = ~rah;  //complement 
assign RCH = ~rch;  //complement 
assign oeh = ~OEH;  //complement 
assign pah = ~PAH;  //complement 
assign DAH =  BAH & QEB  |  BCH & QFB  |  BEH & QGB  |  BGH & QHB  ; 
assign dah = ~DAH;  //complement 
assign aah = ~AAH;  //complement 
assign ach = ~ACH;  //complement 
assign aeh = ~AEH;  //complement 
assign ebh = eah; 
assign EBH = ~ebh; //complement 
assign RAP = ~rap;  //complement 
assign RCP = ~rcp;  //complement 
assign oep = ~OEP;  //complement 
assign pap = ~PAP;  //complement 
assign DAP =  BAP & QED  |  BCP & QFD  |  BEP & QGD  |  BGP & QHD  ; 
assign dap = ~DAP;  //complement 
assign KAH =  AEH & aep  |  aeh & AEP  |  aeh & aep  |  AEH & AEP  ; 
assign kah = ~KAH; //complement 
assign KAP =  AFH & afp  |  afh & AFP  |  afh & afp  |  AFH & AFP  ; 
assign kap = ~KAP; //complement 
assign aap = ~AAP;  //complement 
assign acp = ~ACP;  //complement 
assign aep = ~AEP;  //complement 
assign tda = ~TDA;  //complement 
assign tdb = ~TDB;  //complement 
assign tdc = ~TDC;  //complement 
assign tdd = ~TDD;  //complement 
assign LAH =  PAH & pap  |  pah & PAP  |  pah & pap  |  PAH & PAP  ; 
assign lah = ~LAH; //complement 
assign LAP =  PBH & pbp  |  pbn & PBP  |  pbn & pbp  |  PBH & PBP  ; 
assign lap = ~LAP; //complement 
assign abh = ~ABH;  //complement 
assign adh = ~ADH;  //complement 
assign afh = ~AFH;  //complement 
assign RBH = ~rbh;  //complement 
assign RDH = ~rdh;  //complement 
assign ofh = ~OFH;  //complement 
assign pbh = ~PBH;  //complement 
assign DBH =  BBH & QEF  |  BDH & QFF  |  BFH & QGG  |  BHH & QHF  ; 
assign dbh = ~DBH;  //complement 
assign abp = ~ABP;  //complement 
assign adp = ~ADP;  //complement 
assign afp = ~AFP;  //complement 
assign RBP = ~rbp;  //complement 
assign ofp = ~OFP;  //complement 
assign pbp = ~PBP;  //complement 
assign DBP =  BBP & QEH  |  BDP & QFH  |  BFP & QGH  |  BHP & QHH  ; 
assign dbp = ~DBP;  //complement 
assign bah = ~BAH;  //complement 
assign bap = ~BAP;  //complement 
assign bbh = ~BBH;  //complement 
assign bbp = ~BBP;  //complement 
assign cah = ~CAH;  //complement 
assign oah = ~OAH;  //complement 
assign cap = ~CAP;  //complement 
assign oap = ~OAP;  //complement 
assign eah = ~EAH;  //complement 
assign bch = ~BCH;  //complement 
assign bcp = ~BCP;  //complement 
assign bdh = ~BDH;  //complement 
assign bdp = ~BDP;  //complement 
assign cbh = ~CBH;  //complement 
assign obh = ~OBH;  //complement 
assign cbp = ~CBP;  //complement 
assign obp = ~OBP;  //complement 
assign qkh = ~QKH;  //complement 
assign qlh = ~QLH;  //complement 
assign ogc = ~OGC;  //complement 
assign qkg = ~QKG;  //complement 
assign ogd = ~OGD;  //complement 
assign qlg = ~QLG;  //complement 
assign beh = ~BEH;  //complement 
assign bep = ~BEP;  //complement 
assign bfh = ~BFH;  //complement 
assign bfp = ~BFP;  //complement 
assign cch = ~CCH;  //complement 
assign och = ~OCH;  //complement 
assign ccp = ~CCP;  //complement 
assign ocp = ~OCP;  //complement 
assign tbe = ~TBE;  //complement 
assign tbf = ~TBF;  //complement 
assign tbh = ~TBH;  //complement 
assign tbg = ~TBG;  //complement 
assign bgh = ~BGH;  //complement 
assign bgp = ~BGP;  //complement 
assign bhh = ~BHH;  //complement 
assign bhp = ~BHP;  //complement 
assign cdh = ~CDH;  //complement 
assign odh = ~ODH;  //complement 
assign cdp = ~CDP;  //complement 
assign odp = ~ODP;  //complement 
assign iaa = ~IAA; //complement 
assign iab = ~IAB; //complement 
assign iac = ~IAC; //complement 
assign iad = ~IAD; //complement 
assign iae = ~IAE; //complement 
assign iaf = ~IAF; //complement 
assign iag = ~IAG; //complement 
assign iah = ~IAH; //complement 
assign iai = ~IAI; //complement 
assign iaj = ~IAJ; //complement 
assign iak = ~IAK; //complement 
assign ial = ~IAL; //complement 
assign iam = ~IAM; //complement 
assign ian = ~IAN; //complement 
assign iao = ~IAO; //complement 
assign iap = ~IAP; //complement 
assign iaq = ~IAQ; //complement 
assign ias = ~IAS; //complement 
assign iat = ~IAT; //complement 
assign iba = ~IBA; //complement 
assign ibb = ~IBB; //complement 
assign ibc = ~IBC; //complement 
assign ibd = ~IBD; //complement 
assign ibe = ~IBE; //complement 
assign ibf = ~IBF; //complement 
assign ibg = ~IBG; //complement 
assign ibh = ~IBH; //complement 
assign ibi = ~IBI; //complement 
assign ibj = ~IBJ; //complement 
assign ibk = ~IBK; //complement 
assign ibl = ~IBL; //complement 
assign ibm = ~IBM; //complement 
assign ibn = ~IBN; //complement 
assign ibo = ~IBO; //complement 
assign ibp = ~IBP; //complement 
assign ibq = ~IBQ; //complement 
assign ibs = ~IBS; //complement 
assign ibt = ~IBT; //complement 
assign ica = ~ICA; //complement 
assign icb = ~ICB; //complement 
assign icc = ~ICC; //complement 
assign icd = ~ICD; //complement 
assign ice = ~ICE; //complement 
assign icf = ~ICF; //complement 
assign icg = ~ICG; //complement 
assign ich = ~ICH; //complement 
assign ici = ~ICI; //complement 
assign icj = ~ICJ; //complement 
assign ick = ~ICK; //complement 
assign icl = ~ICL; //complement 
assign icm = ~ICM; //complement 
assign icn = ~ICN; //complement 
assign ico = ~ICO; //complement 
assign icp = ~ICP; //complement 
assign icq = ~ICQ; //complement 
assign ics = ~ICS; //complement 
assign ict = ~ICT; //complement 
assign ida = ~IDA; //complement 
assign idb = ~IDB; //complement 
assign idc = ~IDC; //complement 
assign idd = ~IDD; //complement 
assign ide = ~IDE; //complement 
assign idf = ~IDF; //complement 
assign idg = ~IDG; //complement 
assign idh = ~IDH; //complement 
assign idi = ~IDI; //complement 
assign idj = ~IDJ; //complement 
assign idk = ~IDK; //complement 
assign idl = ~IDL; //complement 
assign idm = ~IDM; //complement 
assign idn = ~IDN; //complement 
assign ido = ~IDO; //complement 
assign idp = ~IDP; //complement 
assign idq = ~IDQ; //complement 
assign ids = ~IDS; //complement 
assign idt = ~IDT; //complement 
assign iea = ~IEA; //complement 
assign ieb = ~IEB; //complement 
assign iec = ~IEC; //complement 
assign ied = ~IED; //complement 
assign iee = ~IEE; //complement 
assign ief = ~IEF; //complement 
assign ieg = ~IEG; //complement 
assign ieh = ~IEH; //complement 
assign iei = ~IEI; //complement 
assign iej = ~IEJ; //complement 
assign iek = ~IEK; //complement 
assign iel = ~IEL; //complement 
assign iem = ~IEM; //complement 
assign ien = ~IEN; //complement 
assign ieo = ~IEO; //complement 
assign iep = ~IEP; //complement 
assign ifa = ~IFA; //complement 
assign ifb = ~IFB; //complement 
assign ifc = ~IFC; //complement 
assign ifd = ~IFD; //complement 
assign ife = ~IFE; //complement 
assign ifff  = ~IFFF ; //complement 
assign ifg = ~IFG; //complement 
assign ifh = ~IFH; //complement 
assign ifi = ~IFI; //complement 
assign ifj = ~IFJ; //complement 
assign ifk = ~IFK; //complement 
assign ifl = ~IFL; //complement 
assign ifm = ~IFM; //complement 
assign ifn = ~IFN; //complement 
assign ifo = ~IFO; //complement 
assign ifp = ~IFP; //complement 
assign iga = ~IGA; //complement 
assign igb = ~IGB; //complement 
assign igc = ~IGC; //complement 
assign igd = ~IGD; //complement 
assign ige = ~IGE; //complement 
assign igf = ~IGF; //complement 
assign igg = ~IGG; //complement 
assign igh = ~IGH; //complement 
assign igi = ~IGI; //complement 
assign igj = ~IGJ; //complement 
assign igk = ~IGK; //complement 
assign igl = ~IGL; //complement 
assign iha = ~IHA; //complement 
assign ihb = ~IHB; //complement 
assign ihc = ~IHC; //complement 
assign ihd = ~IHD; //complement 
assign ihe = ~IHE; //complement 
assign ihf = ~IHF; //complement 
assign ihg = ~IHG; //complement 
assign ihh = ~IHH; //complement 
assign ihi = ~IHI; //complement 
assign ihj = ~IHJ; //complement 
assign ihk = ~IHK; //complement 
assign ihl = ~IHL; //complement 
always@(posedge IZZ )
   begin 
 WAA <= QCB ; 
 gaa <= eba ; 
 gab <= ebb ; 
 gac <= ebc ; 
 gad <= ebd ; 
 gba <= gaa ; 
 gbb <= gab ; 
 gbc <= gac ; 
 gbd <= gad ; 
 gae <= ebe ; 
 gaf <= ebf ; 
 gag <= ebg ; 
 gah <= ebh ; 
 gbe <= gae ; 
 gbf <= gaf ; 
 gbg <= gag ; 
 gbh <= gah ; 
 gai <= ebi ; 
 gaj <= ebj ; 
 gak <= ebk ; 
 gal <= ebl ; 
 gbi <= gai ; 
 gbj <= gaj ; 
 gbk <= gak ; 
 gbl <= gal ; 
 KBA <=  KAA & kai  |  kaa & KAI  |  kaa & kai  |  KAA & KAI  ;
 LBA <=  LAA & lai  |  laa & LAI  |  laa & lai  |  LAA & LAI  ;
 WBA <= QCD ; 
 raa <=  RAA  |  QDA  ; 
 rca <=  RAA  |  QDA  ; 
 OEA <=  DAA & TDA  |  RAA & TDE  |  MAA & TDI  ; 
 PAA <=  DAA & TDA  |  RAA & TDE  |  MAA & TDI  ; 
 AAA <=  AAA & taa  |  IEA & TAA  ; 
 ACA <=  AAA & taa  |  IEA & TAA  ; 
 AEA <=  AAA & taa  |  IEA & TAA  ; 
 rai <=  rai & jai  |  RAI & JAI  |  QDB  ; 
 rci <=  rai & jai  |  RAI & JAI  |  QDB  ; 
 OEI <=  DAI & TDB  |  RAI & TDF  |  MAI & TDJ  ; 
 PAI <=  DAI & TDB  |  RAI & TDF  |  MAI & TDJ  ; 
 AAI <=  AAI & tab  |  IEI & TAB  ; 
 ACI <=  AAI & tab  |  IEI & TAB  ; 
 AEI <=  AAI & tab  |  IEI & TAB  ; 
 QAL <= IHL ; 
 ABA <=  ABA & tac  |  IFA & TAC  ; 
 ADA <=  ABA & tac  |  IFA & TAC  ; 
 AFA <=  ABA & tac  |  IFA & TAC  ; 
 rba <=  rba & jba  |  RBA & JBA  |  QDC  ; 
 rda <=  rba & jba  |  RBA & JBA  |  QDC  ; 
 OFA <=  DBA & TDC  |  RBA & TDG  |  MBA & TDK  ; 
 PBA <=  DBA & TDC  |  RBA & TDG  |  MBA & TDK  ; 
 ABI <=  ABI & tad  |  IFI & TAD  ; 
 ADI <=  ABI & tad  |  IFI & TAD  ; 
 AFI <=  ABI & tad  |  IFI & TAD  ; 
 rbi <=  rbi & jbi  |  RBI & JBI  |  QDD  ; 
 rdi <=  rbi & jbi  |  RBI & JBI  |  QDD  ; 
 OFI <=  DBI & TDD  |  RBI & TDH  |  MBI & TDL  ; 
 PBI <=  DBI & TDD  |  RBI & TDH  |  MBI & TDL  ; 
 BAA <=  BAA & tba  |  CAA & TBA  ; 
 BAI <=  BAI & tba  |  CAI & TBA  ; 
 BBA <=  BBA & tbb  |  CAA & TBB  ; 
 BBI <=  BBI & tbb  |  CAI & TBB  ; 
 CAA <=  IAA & TCA  |  ABA & TCC  |  AAA & TCE  ; 
 OAA <=  IAA & TCA  |  ABA & TCC  |  AAA & TCE  ; 
 CAI <=  IAI & TCB  |  ABI & TCD  |  AAI & TCF  ; 
 OAI <=  IAI & TCB  |  ABI & TCD  |  AAI & TCF  ; 
 EAA <=  EBA & TEA  |  IGA & TEB  |  AAA & TEC  ; 
 EAI <=  EBI & TEA  |  IGI & TEB  |  AAI & TEC  ; 
 BCA <=  BCA & tbc  |  CBA & TBC  ; 
 BCI <=  BCI & tbc  |  CBI & TBC  ; 
 BDA <=  BDA & tbd  |  CBA & TBD  ; 
 BDI <=  BDI & tbd  |  CBI & TBD  ; 
 CBA <=  IBA & TCG  |  ABA & TCI  |  AAA & TCK  ; 
 OBA <=  IBA & TCG  |  ABA & TCI  |  AAA & TCK  ; 
 CBI <=  IBI & TCH  |  ABI & TCJ  |  AAI & TCL  ; 
 OBI <=  IBI & TCH  |  ABI & TCJ  |  AAI & TCL  ; 
 QIC <= QBE ; 
 QID <= QIC ; 
 QIE <= QID ; 
 QIF <= QIE ; 
 QIA <=  QBA  |  QBE  |  QIC  |  QID  ; 
 qba <=  ihc  |  IHB  |  IHA  ; 
 qbe <=  ihd  |  IHB  |  IHA  ; 
 qma <=  qma & qba  |  QAK  |  QBE  ; 
 oas <=  ias  |  QAK  |  QMA  ; 
 QIB <=  QBA  |  QBE  |  QIA  ; 
 oaq <= qba ; 
 oar <= qbe ; 
 oat <= ZZI ; 
 BEA <=  BEA & tbe  |  CCA & TBE  ; 
 BEI <=  BEI & tbe  |  CCI & TBE  ; 
 BFA <=  BFA & tbf  |  CCA & TBF  ; 
 BFI <=  BFI & tbf  |  CCI & TBF  ; 
 CCA <=  ICA & TCM  |  ABA & TCO  |  AAA & TCQ  ; 
 OCA <=  ICA & TCM  |  ABA & TCO  |  AAA & TCQ  ; 
 CCI <=  ICI & TCN  |  ABI & TCP  |  AAI & TCR  ; 
 OCI <=  ICI & TCN  |  ABI & TCP  |  AAI & TCR  ; 
 BGA <=  BGA & tbg  |  CDA & TBG  ; 
 BGI <=  BGI & tbg  |  CDI & TBG  ; 
 BHA <=  BHA & tbh  |  CDA & TBH  ; 
 BHI <=  BHI & tbh  |  CDI & TBH  ; 
 CDA <=  IDA & TCS  |  ABA & TCU  |  AAA & TCW  ; 
 ODA <=  IDA & TCS  |  ABA & TCU  |  AAA & TCW  ; 
 CDI <=  IDI & TCT  |  ABI & TCV  |  AAI & TCX  ; 
 ODI <=  IDI & TCT  |  ABI & TCV  |  AAI & TCX  ; 
 WAB <= QCB ; 
 KBB <=  KAB & kaj  |  kab & KAJ  |  kab & kaj  |  KAB & KAJ  ;
 LBB <=  LAB & laj  |  lab & LAJ  |  lab & laj  |  LAB & LAJ  ;
 rab <=  rab & jab  |  RAB & JAB  |  QDA  ; 
 rcb <=  rab & jab  |  RAB & JAB  |  QDA  ; 
 OEB <=  DAB & TDA  |  RAB & TDE  |  MAB & TDI  ; 
 PAB <=  DAB & TDA  |  RAB & TDE  |  MAB & TDI  ; 
 AAB <=  AAB & taa  |  IEB & TAA  ; 
 ACB <=  AAB & taa  |  IEB & TAA  ; 
 AEB <=  AAB & taa  |  IEB & TAA  ; 
 raj <=  raj & jaj  |  RAJ & JAJ  |  QDB  ; 
 rcj <=  raj & jaj  |  RAJ & JAJ  |  QDB  ; 
 OEJ <=  DAJ & TDB  |  RAJ & TDF  |  MAJ & TDJ  ; 
 PAJ <=  DAJ & TDB  |  RAJ & TDF  |  MAJ & TDJ  ; 
 AAJ <=  AAJ & tab  |  IEJ & TAB  ; 
 ACJ <=  AAJ & tab  |  IEJ & TAB  ; 
 AEJ <=  AAJ & tab  |  IEJ & TAB  ; 
 ABB <=  ABB & tac  |  IFB & TAC  ; 
 ADB <=  ABB & tac  |  IFB & TAC  ; 
 AFB <=  ABB & tac  |  IFB & TAC  ; 
 rbb <=  rbb & jbb  |  RBB & JBB  |  QDC  ; 
 rdb <=  rbb & jbb  |  RBB & JBB  |  QDC  ; 
 OFB <=  DBB & TDC  |  RBB & TDG  |  MBB & TDK  ; 
 PBB <=  DBB & TDC  |  RBB & TDG  |  MBB & TDK  ; 
 ABJ <=  ABJ & tad  |  IFJ & TAD  ; 
 ADJ <=  ABJ & tad  |  IFJ & TAD  ; 
 AFJ <=  ABJ & tad  |  IFJ & TAD  ; 
 rbj <=  rbj & jbj  |  RBJ & JBJ  |  QDD  ; 
 rdj <=  rbj & jbj  |  RBJ & JBJ  |  QDD  ; 
 OFJ <=  DBJ & TDD  |  RBJ & TDH  |  MBJ & TDL  ; 
 PBJ <=  DBJ & TDD  |  RBJ & TDH  |  MBJ & TDL  ; 
 BAB <=  BAB & tba  |  CAB & TBA  ; 
 BAJ <=  BAJ & tba  |  CAJ & TBA  ; 
 BBB <=  BBB & tbb  |  CAB & TBB  ; 
 BBJ <=  BBJ & tbb  |  CAJ & TBB  ; 
 CAB <=  IAB & TCA  |  ABB & TCC  |  AAB & TCE  ; 
 OAB <=  IAB & TCA  |  ABB & TCC  |  AAB & TCE  ; 
 CAJ <=  IAJ & TCB  |  ABJ & TCD  |  AAJ & TCF  ; 
 OAJ <=  IAJ & TCB  |  ABJ & TCD  |  AAJ & TCF  ; 
 EAB <=  EBB & TEA  |  IGB & TEB  |  AAB & TEC  ; 
 EAJ <=  EBJ & TEA  |  IGJ & TEB  |  AAJ & TEC  ; 
 BCB <=  BCB & tbc  |  CBB & TBC  ; 
 BCJ <=  BCJ & tbc  |  CBJ & TBC  ; 
 BDB <=  BDB & tbd  |  CBB & TBD  ; 
 BDJ <=  BDJ & tbd  |  CBJ & TBD  ; 
 CBB <=  IBB & TCG  |  ABB & TCI  |  AAB & TCK  ; 
 OBB <=  IBB & TCG  |  ABB & TCI  |  AAB & TCK  ; 
 CBJ <=  IBJ & TCH  |  ABJ & TCJ  |  AAJ & TCL  ; 
 OBJ <=  IBJ & TCH  |  ABJ & TCJ  |  AAJ & TCL  ; 
 QJC <= QBF ; 
 QJD <= QJC ; 
 QJE <= QJD ; 
 QJF <= QJE ; 
 QJA <=  QBB  |  QBF  |  QJC  |  QJD  ; 
 qbb <=  ihc  |  IHB  |  iha  ; 
 qbf <=  ihd  |  IHB  |  iha  ; 
 qmb <=  qmb & qbb  |  QAK  |  QBF  ; 
 obs <=  ibs  |  QAK  |  QMB  ; 
 QJB <=  QBB  |  QBF  |  QJA  ; 
 obq <= qbb ; 
 obr <= qbf ; 
 obt <= ZZI ; 
 BEB <=  BEB & tbe  |  CCB & TBE  ; 
 BEJ <=  BEJ & tbe  |  CCJ & TBE  ; 
 BFB <=  BFB & tbf  |  CCB & TBF  ; 
 BFJ <=  BFJ & tbf  |  CCJ & TBF  ; 
 CCB <=  ICB & TCM  |  ABB & TCO  |  AAB & TCQ  ; 
 OCB <=  ICB & TCM  |  ABB & TCO  |  AAB & TCQ  ; 
 CCJ <=  ICJ & TCN  |  ABJ & TCP  |  AAJ & TCR  ; 
 OCJ <=  ICJ & TCN  |  ABJ & TCP  |  AAJ & TCR  ; 
 BGB <=  BGB & tbg  |  CDB & TBG  ; 
 BGJ <=  BGJ & tbg  |  CDJ & TBG  ; 
 BHB <=  BHB & tbh  |  CDB & TBH  ; 
 BHJ <=  BHJ & tbh  |  CDJ & TBH  ; 
 CDB <=  IDB & TCS  |  ABB & TCU  |  AAB & TCW  ; 
 ODB <=  IDB & TCS  |  ABB & TCU  |  AAB & TCW  ; 
 CDJ <=  IDJ & TCT  |  ABJ & TCV  |  AAJ & TCX  ; 
 ODJ <=  IDJ & TCT  |  ABJ & TCV  |  AAJ & TCX  ; 
 WAC <= QCB ; 
 KBC <=  KAC & kak  |  kac & KAK  |  kac & kak  |  KAC & KAK  ;
 LBC <=  LAC & lak  |  lac & LAK  |  lac & lak  |  LAC & LAK  ;
 had <=  jaq  |  jar  |  jas  |  jat  ; 
 hae <=  jaq  |  jar  |  jas  |  jat  ; 
 rac <=  rac & jac  |  RAC & JAC  |  QDA  ; 
 rcc <=  rac & jac  |  RAC & JAC  |  QDA  ; 
 OEC <=  DAC & TDA  |  RAC & TDE  |  MAC & TDI  ; 
 PAC <=  DAC & TDA  |  RAC & TDE  |  MAC & TDI  ; 
 AAC <=  AAC & taa  |  IEC & TAA  ; 
 ACC <=  AAC & taa  |  IEC & TAA  ; 
 AEC <=  AAC & taa  |  IEC & TAA  ; 
 rak <=  rak & jak  |  RAK & JAK  |  QDB  ; 
 rck <=  rak & jak  |  RAK & JAK  |  QDB  ; 
 OEK <=  DAK & TDB  |  RAK & TDF  |  MAK & TDJ  ; 
 PAK <=  DAK & TDB  |  RAK & TDF  |  MAK & TDJ  ; 
 AAK <=  AAK & tab  |  IEK & TAB  ; 
 ACK <=  AAK & tab  |  IEK & TAB  ; 
 AEK <=  AAK & tab  |  IEK & TAB  ; 
 ABC <=  ABC & tac  |  IFC & TAC  ; 
 ADC <=  ABC & tac  |  IFC & TAC  ; 
 AFC <=  ABC & tac  |  IFC & TAC  ; 
 rbc <=  rbc & jbc  |  RBC & JBC  |  QDC  ; 
 rdc <=  rbc & jbc  |  RBC & JBC  |  QDC  ; 
 OFC <=  DBC & TDC  |  RBC & TDG  |  MBC & TDK  ; 
 PBC <=  DBC & TDC  |  RBC & TDG  |  MBC & TDK  ; 
 ABK <=  ABK & tad  |  IFK & TAD  ; 
 ADK <=  ABK & tad  |  IFK & TAD  ; 
 AFK <=  ABK & tad  |  IFK & TAD  ; 
 rbk <=  rbk & jbk  |  RBK & JBK  |  QDD  ; 
 rdk <=  rbk & jbk  |  RBK & JBK  |  QDD  ; 
 OFK <=  DBK & TDD  |  RBK & TDH  |  MBK & TDL  ; 
 PBK <=  DBK & TDD  |  RBK & TDH  |  MBK & TDL  ; 
 BAC <=  BAC & tba  |  CAC & TBA  ; 
 BAK <=  BAK & tba  |  CAK & TBA  ; 
 BBC <=  BBC & tbb  |  CAC & TBB  ; 
 BBK <=  BBK & tbb  |  CAK & TBB  ; 
 CAC <=  IAC & TCA  |  ABC & TCC  |  AAC & TCE  ; 
 OAC <=  IAC & TCA  |  ABC & TCC  |  AAC & TCE  ; 
 CAK <=  IAK & TCB  |  ABK & TCD  |  AAK & TCF  ; 
 OAK <=  IAK & TCB  |  ABK & TCD  |  AAK & TCF  ; 
 EAC <=  EBC & TEA  |  IGC & TEB  |  AAC & TEC  ; 
 EAK <=  EBK & TEA  |  IGK & TEB  |  AAK & TEC  ; 
 BCC <=  BCC & tbc  |  CBC & TBC  ; 
 BCK <=  BCK & tbc  |  CBK & TBC  ; 
 BDC <=  BDC & tbd  |  CBC & TBD  ; 
 BDK <=  BDK & tbd  |  CBK & TBD  ; 
 CBC <=  IBC & TCG  |  ABC & TCI  |  AAC & TCK  ; 
 OBC <=  IBC & TCG  |  ABC & TCI  |  AAC & TCK  ; 
 CBK <=  IBK & TCH  |  ABK & TCJ  |  AAK & TCL  ; 
 OBK <=  IBK & TCH  |  ABK & TCJ  |  AAK & TCL  ; 
 QKC <= QBG ; 
 QKD <= QKC ; 
 QKE <= QKD ; 
 QKF <= QKE ; 
 QKA <=  QBC  |  QBG  |  QKC  |  QKD  ; 
 qbc <=  ihc  |  ihb  |  IHA  ; 
 qbg <=  ihd  |  ihb  |  IHA  ; 
 qmc <=  qmc & qbc  |  QAK  |  QBG  ; 
 ocs <=  ics  |  QAK  |  QMC  ; 
 QKB <=  QBC  |  QBG  |  QKA  ; 
 ocq <= qbc ; 
 ocr <= qbg ; 
 oct <= ZZI ; 
 BEC <=  BEC & tbe  |  CCC & TBE  ; 
 BEK <=  BEK & tbe  |  CCK & TBE  ; 
 BFC <=  BFC & tbf  |  CCC & TBF  ; 
 BFK <=  BFK & tbf  |  CCK & TBF  ; 
 CCC <=  ICC & TCM  |  ABC & TCO  |  AAC & TCQ  ; 
 OCC <=  ICC & TCM  |  ABC & TCO  |  AAC & TCQ  ; 
 CCK <=  ICK & TCN  |  ABK & TCP  |  AAK & TCR  ; 
 OCK <=  ICK & TCN  |  ABK & TCP  |  AAK & TCR  ; 
 BGC <=  BGC & tbg  |  CDC & TBG  ; 
 BGK <=  BGK & tbg  |  CDK & TBG  ; 
 BHC <=  BHC & tbh  |  CDC & TBH  ; 
 BHK <=  BHK & tbh  |  CDK & TBH  ; 
 CDC <=  IDC & TCS  |  ABC & TCU  |  AAC & TCW  ; 
 ODC <=  IDC & TCS  |  ABC & TCU  |  AAC & TCW  ; 
 CDK <=  IDK & TCT  |  ABK & TCV  |  AAK & TCX  ; 
 ODK <=  IDK & TCT  |  ABK & TCV  |  AAK & TCX  ; 
 WAD <= QCB ; 
 KDA <=  KCA & kcb & kcc  |  kca & KCB & kcc  |  kca & kcb & KCC  |  KCA & KCB & KCC  ;
 KBD <=  KAD & kal  |  kad & KAL  |  kad & kal  |  KAD & KAL  ;
 LBD <=  LAD & lal  |  lad & LAL  |  lad & lal  |  LAD & LAL  ;
 haf <=  jaq  |  jar  |  jas  |  jat  ; 
 hag <=  jaq  |  jar  |  jas  |  jat  ; 
 rad <=  rad & jad  |  RAD & JAD  |  QDA  ; 
 rcd <=  rad & jad  |  RAD & JAD  |  QDA  ; 
 PAD <=  DAD & TDA  |  RAD & TDE  |  MAD & TDI  ; 
 OED <=  DAD & TDA  |  RAD & TDE  |  MAD & TDI  ; 
 AAD <=  AAD & taa  |  IED & TAA  ; 
 ACD <=  AAD & taa  |  IED & TAA  ; 
 AED <=  AAD & taa  |  IED & TAA  ; 
 QEA <= JCA ; 
 QFA <= JCB ; 
 QGA <= JCC ; 
 QHA <= JCD ; 
 ral <=  ral & jal  |  RAL & JAL  |  QDB  ; 
 rcl <=  ral & jal  |  RAL & JAL  |  QDB  ; 
 PAL <=  DAL & TDB  |  RAL & TDF  |  MAL & TDJ  ; 
 OEL <=  DAL & TDB  |  RAL & TDF  |  MAL & TDJ  ; 
 AAL <=  AAL & tab  |  IEL & TAB  ; 
 ACL <=  AAL & tab  |  IEL & TAB  ; 
 AEL <=  AAL & tab  |  IEL & TAB  ; 
 QEC <= JCA ; 
 QFC <= JCB ; 
 QGC <= JCC ; 
 QHC <= JCD ; 
 ABD <=  ABD & tac  |  IFD & TAC  ; 
 ADD <=  ABD & tac  |  IFD & TAC  ; 
 AFD <=  ABD & tac  |  IFD & TAC  ; 
 qee <= jca ; 
 qfe <= jcb ; 
 qge <= jcc ; 
 qhe <= jcd ; 
 rbd <=  rbd & jbd  |  RBD & JBD  |  QDC  ; 
 rdd <=  rbd & jbd  |  RBD & JBD  |  QDC  ; 
 OFD <=  DBD & TDC  |  RBD & TDG  |  MBD & TDK  ; 
 PBD <=  DBD & TDC  |  RBD & TDG  |  MBD & TDK  ; 
 ABL <=  ABL & tad  |  IFL & TAD  ; 
 ADL <=  ABL & tad  |  IFL & TAD  ; 
 AFL <=  ABL & tad  |  IFL & TAD  ; 
 qeg <= jca ; 
 qfg <= jcb ; 
 qgg <= jcc ; 
 qhg <= jcd ; 
 rbl <=  rbl & jbl  |  RBL & JBL  |  QDD  ; 
 rdl <=  rbl & jbl  |  RBL & JBL  |  QDD  ; 
 OFL <=  DBL & TDD  |  RBL & TDH  |  MBL & TDL  ; 
 PBL <=  DBL & TDD  |  RBL & TDH  |  MBL & TDL  ; 
 BAD <=  BAD & tba  |  CAD & TBA  ; 
 BAL <=  BAL & tba  |  CAL & TBA  ; 
 BBD <=  BBD & tbb  |  CAD & TBB  ; 
 BBL <=  BBL & tbb  |  CAL & TBB  ; 
 CAD <=  IAD & TCA  |  ABD & TCC  |  AAD & TCE  ; 
 OAD <=  IAD & TCA  |  ABD & TCC  |  AAD & TCE  ; 
 CAL <=  IAL & TCB  |  ABL & TCD  |  AAL & TCF  ; 
 OAL <=  IAL & TCB  |  ABL & TCD  |  AAL & TCF  ; 
 EAD <=  EBD & TEA  |  IGD & TEB  |  AAD & TEC  ; 
 EAL <=  EBL & TEA  |  IGL & TEB  |  AAL & TEC  ; 
 BCD <=  BCD & tbc  |  CBD & TBC  ; 
 BCL <=  BCL & tbc  |  CBL & TBC  ; 
 BDD <=  BDD & tbd  |  CBD & TBD  ; 
 BDL <=  BDL & tbd  |  CBL & TBD  ; 
 CBD <=  IBD & TCG  |  ABD & TCI  |  AAD & TCK  ; 
 OBD <=  IBD & TCG  |  ABD & TCI  |  AAD & TCK  ; 
 CBL <=  IBL & TCH  |  ABL & TCJ  |  AAL & TCL  ; 
 OBL <=  IBL & TCH  |  ABL & TCJ  |  AAL & TCL  ; 
 QLC <= QBH ; 
 QLD <= QLC ; 
 QLE <= QLD ; 
 QLF <= QLE ; 
 QLA <=  QBD  |  QBH  |  QLC  |  QLD  ; 
 qbd <=  ihc  |  ihb  |  iha  ; 
 qbh <=  ihd  |  ihb  |  iha  ; 
 qmd <=  qmd & qbd  |  QAK  |  QBH  ; 
 ods <=  ids  |  QAK  |  QMD  ; 
 QLB <=  QBD  |  QBH  |  QLA  ; 
 odq <= qbd ; 
 odr <= qbh ; 
 odt <= ZZI ; 
 BED <=  BED & tbe  |  CCD & TBE  ; 
 BEL <=  BEL & tbe  |  CCL & TBE  ; 
 BFD <=  BFD & tbf  |  CCD & TBF  ; 
 BFL <=  BFL & tbf  |  CCL & TBF  ; 
 CCD <=  ICD & TCM  |  ABD & TCO  |  AAD & TCQ  ; 
 OCD <=  ICD & TCM  |  ABD & TCO  |  AAD & TCQ  ; 
 CCL <=  ICL & TCN  |  ABL & TCP  |  AAL & TCR  ; 
 OCL <=  ICL & TCN  |  ABL & TCP  |  AAL & TCR  ; 
 BGD <=  BGD & tbg  |  CDD & TBG  ; 
 BGL <=  BGL & tbg  |  CDL & TBG  ; 
 BHD <=  BHD & tbh  |  CDD & TBH  ; 
 BHL <=  BHL & tbh  |  CDL & TBH  ; 
 CDD <=  IDD & TCS  |  ABD & TCU  |  AAD & TCW  ; 
 ODD <=  IDD & TCS  |  ABD & TCU  |  AAD & TCW  ; 
 CDL <=  IDL & TCT  |  ABL & TCV  |  AAL & TCX  ; 
 ODL <=  IDL & TCT  |  ABL & TCV  |  AAL & TCX  ; 
 WAE <= QCB ; 
 HAA <=  JAQ  ; 
 KBE <=  KAE & kam  |  kae & KAM  |  kae & kam  |  KAE & KAM  ;
 LDA <=  LCA & lcb & lcc  |  lca & LCB & lcc  |  lca & lcb & LCC  |  LCA & LCB & LCC  ;
 LBE <=  LAE & lam  |  lae & LAM  |  lae & lam  |  LAE & LAM  ;
 HBA <=  JBQ  ; 
 rae <=  rae & jae  |  RAE & JAE  |  QDA  ; 
 rce <=  rae & jae  |  RAE & JAE  |  QDA  ; 
 OEE <=  DAE & TDA  |  RAE & TDE  |  MAE & TDI  ; 
 PAE <=  DAE & TDA  |  RAE & TDE  |  MAE & TDI  ; 
 AAE <=  AAE & taa  |  IEE & TAA  ; 
 ACE <=  AAE & taa  |  IEE & TAA  ; 
 AEE <=  AAE & taa  |  IEE & TAA  ; 
 QEB <= JCA ; 
 QFB <= JCB ; 
 QGB <= JCC ; 
 QHB <= JCD ; 
 ram <=  ram & jam  |  RAM & JAM  |  QDB  ; 
 rcm <=  ram & jam  |  RAM & JAM  |  QDB  ; 
 OEM <=  DAM & TDB  |  RAM & TDF  |  MAM & TDJ  ; 
 PAM <=  DAM & TDB  |  RAM & TDF  |  MAM & TDJ  ; 
 AAM <=  AAM & tab  |  IEM & TAB  ; 
 ACM <=  AAM & tab  |  IEM & TAB  ; 
 AEM <=  AAM & tab  |  IEM & TAB  ; 
 QED <= JCA ; 
 QFD <= JCB ; 
 QGD <= JCC ; 
 QHD <= JCD ; 
 ABE <=  ABE & tac  |  IFE & TAC  ; 
 ADE <=  ABE & tac  |  IFE & TAC  ; 
 AFE <=  ABE & tac  |  IFE & TAC  ; 
 qef <= jca ; 
 qff <= jcb ; 
 qgf <= jcc ; 
 qhf <= jcd ; 
 rbe <=  rbe & jbe  |  RBE & JBE  |  QDC  ; 
 rde <=  rbe & jbe  |  RBE & JBE  |  QDC  ; 
 OFE <=  DBE & TDC  |  RBE & TDG  |  MBE & TDK  ; 
 PBE <=  DBE & TDC  |  RBE & TDG  |  MBE & TDK  ; 
 ABM <=  ABM & tad  |  IFM & TAD  ; 
 ADM <=  ABM & tad  |  IFM & TAD  ; 
 AFM <=  ABM & tad  |  IFM & TAD  ; 
 qgh <= jcc ; 
 qhh <= jcd ; 
 qeh <= jca ; 
 qfh <= jcb ; 
 rbm <=  rbm & jbm  |  RBM & JBM  |  QDD  ; 
 rdm <=  rbm & jbm  |  RBM & JBM  |  QDD  ; 
 OFM <=  DBM & TDD  |  RBM & TDH  |  MBM & TDL  ; 
 PBM <=  DBM & TDD  |  RBM & TDH  |  MBM & TDL  ; 
 BAE <=  BAE & tba  |  CAE & TBA  ; 
 BAM <=  BAM & tba  |  CAM & TBA  ; 
 BBE <=  BBE & tbb  |  CAE & TBB  ; 
 BBM <=  BBM & tbb  |  CAM & TBB  ; 
 CAE <=  IAE & TCA  |  ABE & TCC  |  AAE & TCE  ; 
 OAE <=  IAE & TCA  |  ABE & TCC  |  AAE & TCE  ; 
 CAM <=  IAM & TCB  |  ABM & TCD  |  AAM & TCF  ; 
 OAM <=  IAM & TCB  |  ABM & TCD  |  AAM & TCF  ; 
 EAE <=  EBE & TEA  |  IGE & TEB  |  AAE & TEC  ; 
 BCE <=  BCE & tbc  |  CBE & TBC  ; 
 BCM <=  BCM & tbc  |  CBM & TBC  ; 
 BDE <=  BDE & tbd  |  CBE & TBD  ; 
 BDM <=  BDM & tbd  |  CBM & TBD  ; 
 CBE <=  IBE & TCG  |  ABE & TCI  |  AAE & TCK  ; 
 OBE <=  IBE & TCG  |  ABE & TCI  |  AAE & TCK  ; 
 CBM <=  IBM & TCH  |  ABM & TCJ  |  AAM & TCL  ; 
 OBM <=  IBM & TCH  |  ABM & TCJ  |  AAM & TCL  ; 
 QAA <= IHA ; 
 QAB <= IHB ; 
 QAE <= IHE ; 
 BEE <=  BEE & tbe  |  CCE & TBE  ; 
 BEM <=  BEM & tbe  |  CCM & TBE  ; 
 BFE <=  BFE & tbf  |  CCE & TBF  ; 
 BFM <=  BFM & tbf  |  CCM & TBF  ; 
 CCE <=  ICE & TCM  |  ABE & TCO  |  AAE & TCQ  ; 
 OCE <=  ICE & TCM  |  ABE & TCO  |  AAE & TCQ  ; 
 CCM <=  ICM & TCN  |  ABM & TCP  |  AAM & TCR  ; 
 OCM <=  ICM & TCN  |  ABM & TCP  |  AAM & TCR  ; 
 BGE <=  BGE & tbg  |  CDE & TBG  ; 
 BGM <=  BGM & tbg  |  CDM & TBG  ; 
 BHE <=  BHE & tbh  |  CDE & TBH  ; 
 BHM <=  BHM & tbh  |  CDM & TBH  ; 
 CDE <=  IDE & TCS  |  ABE & TCU  |  AAE & TCW  ; 
 ODE <=  IDE & TCS  |  ABE & TCU  |  AAE & TCW  ; 
 CDM <=  IDM & TCT  |  ABM & TCV  |  AAM & TCX  ; 
 ODM <=  IDM & TCT  |  ABM & TCV  |  AAM & TCX  ; 
 WAF <= QCB ; 
 QCA <=  QAH  ; 
 QCB <=  QAH  |  QCA  ; 
 HAB <=  JAQ & JAR  ; 
 qcc <= qcb ; 
 qcd <= qcc ; 
 qce <= tdi ; 
 qcf <= qce ; 
 KBF <=  KAF & kan  |  kaf & KAN  |  kaf & kan  |  KAF & KAN  ;
 LBF <=  LAF & lan  |  laf & LAN  |  laf & lan  |  LAF & LAN  ;
 QCG <= QCF ; 
 QCH <=  LEA & QCG  ; 
 HBB <=  JBQ & JBR  ; 
 PBQ <=  MBQ & QCF  ; 
 raf <=  raf & jaf  |  RAF & JAF  |  QDA  ; 
 rcf <=  raf & jaf  |  RAF & JAF  |  QDA  ; 
 PAF <=  DAF & TDA  |  RAF & TDE  |  MAF & TDI  ; 
 OEF <=  DAF & TDA  |  RAF & TDE  |  MAF & TDI  ; 
 qda <= qak ; 
 qdb <= qak ; 
 AAF <=  AAF & taa  |  IEF & TAA  ; 
 ACF <=  AAF & taa  |  IEF & TAA  ; 
 AEF <=  AAF & taa  |  IEF & TAA  ; 
 ran <=  ran & jan  |  RAN & JAN  |  QDB  ; 
 rcn <=  ran & jan  |  RAN & JAN  |  QDB  ; 
 PAN <=  DAN & TDB  |  RAN & TDF  |  MAN & TDJ  ; 
 OEN <=  DAN & TDB  |  RAN & TDF  |  MAN & TDJ  ; 
 AAN <=  AAN & tab  |  IEN & TAB  ; 
 ACN <=  AAN & tab  |  IEN & TAB  ; 
 AEN <=  AAN & tab  |  IEN & TAB  ; 
 QAG <= qcb & IHG ; 
 QAH <= qcb & IHH ; 
 ABF <=  ABF & tac  |  IFFF  & TAC  ; 
 ADF <=  ABF & tac  |  IFFF  & TAC  ; 
 AFF <=  ABF & tac  |  IFFF  & TAC  ; 
 rbf <=  rbf & jbf  |  RBF & JBF  |  QDC  ; 
 rdf <=  rbf & jbf  |  RBF & JBF  |  QDC  ; 
 PBF <=  DBF & TDC  |  RBF & TDG  |  MBF & TDK  ; 
 OFF <=  DBF & TDC  |  RBF & TDG  |  MBF & TDK  ; 
 qdc <= qak ; 
 qdd <= qak ; 
 ABN <=  ABN & tad  |  IFN & TAD  ; 
 ADN <=  ABN & tad  |  IFN & TAD  ; 
 AFN <=  ABN & tad  |  IFN & TAD  ; 
 rbn <=  rbn & jbn  |  RBN & JBN  |  QDD  ; 
 rdn <=  rbn & jbn  |  RBN & JBN  |  QDD  ; 
 PBN <=  DBN & TDD  |  RBN & TDH  |  MBN & TDL  ; 
 OFN <=  DBN & TDD  |  RBN & TDH  |  MBN & TDL  ; 
 BAF <=  BAF & tba  |  CAF & TBA  ; 
 BAN <=  BAN & tba  |  CAN & TBA  ; 
 BBF <=  BBF & tbb  |  CAF & TBB  ; 
 BBN <=  BBN & tbb  |  CAN & TBB  ; 
 CAF <=  IAF & TCA  |  ABF & TCC  |  AAF & TCE  ; 
 OAF <=  IAF & TCA  |  ABF & TCC  |  AAF & TCE  ; 
 CAN <=  IAN & TCB  |  ABN & TCD  |  AAN & TCF  ; 
 OAN <=  IAN & TCB  |  ABN & TCD  |  AAN & TCF  ; 
 EAF <=  EBF & TEA  |  IGF & TEB  |  AAF & TEC  ; 
 BCF <=  BCF & tbc  |  CBF & TBC  ; 
 BCN <=  BCN & tbc  |  CBN & TBC  ; 
 BDF <=  BDF & tbd  |  CBF & TBD  ; 
 BDN <=  BDN & tbd  |  CBN & TBD  ; 
 CBF <=  IBF & TCG  |  ABF & TCI  |  AAF & TCK  ; 
 OBF <=  IBF & TCG  |  ABF & TCI  |  AAF & TCK  ; 
 CBN <=  IBN & TCH  |  ABN & TCJ  |  AAN & TCL  ; 
 OBN <=  IBN & TCH  |  ABN & TCJ  |  AAN & TCL  ; 
 QAI <= IHI ; 
 QAJ <= IHJ ; 
 OHA <= QCH ; 
 QAK <= IHK ; 
 BEF <=  BEF & tbe  |  CCF & TBE  ; 
 BEN <=  BEN & tbe  |  CCN & TBE  ; 
 BFF <=  BFF & tbf  |  CCF & TBF  ; 
 BFN <=  BFN & tbf  |  CCN & TBF  ; 
 CCF <=  ICF & TCM  |  ABF & TCO  |  AAF & TCQ  ; 
 OCF <=  ICF & TCM  |  ABF & TCO  |  AAF & TCQ  ; 
 CCN <=  ICN & TCN  |  ABN & TCP  |  AAN & TCR  ; 
 OCN <=  ICN & TCN  |  ABN & TCP  |  AAN & TCR  ; 
 BGF <=  BGF & tbg  |  CDF & TBG  ; 
 BGN <=  BGN & tbg  |  CDN & TBG  ; 
 BHF <=  BHF & tbh  |  CDF & TBH  ; 
 BHN <=  BHN & tbh  |  CDN & TBH  ; 
 CDF <=  IDF & TCS  |  ABF & TCU  |  AAF & TCW  ; 
 ODF <=  IDF & TCS  |  ABF & TCU  |  AAF & TCW  ; 
 CDN <=  IDN & TCT  |  ABN & TCV  |  AAN & TCX  ; 
 ODN <=  IDN & TCT  |  ABN & TCV  |  AAN & TCX  ; 
 WAG <= QCB ; 
 HAC <=  JAQ & JAR & JAS  ; 
 KBG <=  KAG & kao  |  kag & KAO  |  kag & kao  |  KAG & KAO  ;
 LBG <=  LAG & lao  |  lag & LAO  |  lag & lao  |  LAG & LAO  ;
 HBC <=  JBQ & JBR & JBS  ; 
 rag <=  rag & jag  |  RAG & JAG  |  QDA  ; 
 rcg <=  rag & jag  |  RAG & JAG  |  QDA  ; 
 OEG <=  DAG & TDA  |  RAG & TDE  |  MAG & TDI  ; 
 PAG <=  DAG & TDA  |  RAG & TDE  |  MAG & TDI  ; 
 AAG <=  AAG & taa  |  IEG & TAA  ; 
 ACG <=  AAG & taa  |  IEG & TAA  ; 
 AEG <=  AAG & taa  |  IEG & TAA  ; 
 rao <=  rao & jao  |  RAO & JAO  |  QDB  ; 
 rco <=  rao & jao  |  RAO & JAO  |  QDB  ; 
 OEO <=  DAO & TDB  |  RAO & TDF  |  MAO & TDJ  ; 
 PAO <=  DAO & TDB  |  RAO & TDF  |  MAO & TDJ  ; 
 AAO <=  AAO & tab  |  IEO & TAB  ; 
 ACO <=  AAO & tab  |  IEO & TAB  ; 
 AEO <=  AAO & tab  |  IEO & TAB  ; 
 QAF <= IHF ; 
 ABG <=  ABG & tac  |  IFG & TAC  ; 
 ADG <=  ABG & tac  |  IFG & TAC  ; 
 AFG <=  ABG & tac  |  IFG & TAC  ; 
 rbg <=  rbg & jbg  |  RBG & JBG  |  QDC  ; 
 rdg <=  rbg & jbg  |  RBG & JBG  |  QDC  ; 
 OFG <=  DBG & TDC  |  RBG & TDG  |  MBG & TDK  ; 
 PBG <=  DBG & TDC  |  RBG & TDG  |  MBG & TDK  ; 
 ABO <=  ABO & tad  |  IFO & TAD  ; 
 ADO <=  ABO & tad  |  IFO & TAD  ; 
 AFO <=  ABO & tad  |  IFO & TAD  ; 
 rbo <=  rbo & jbo  |  RBO & JBO  |  QDD  ; 
 rdo <=  rbo & jbo  |  RBO & JBO  |  QDD  ; 
 OFO <=  DBO & TDD  |  RBO & TDH  |  MBO & TDL  ; 
 PBO <=  DBO & TDD  |  RBO & TDH  |  MBO & TDL  ; 
 BAG <=  BAG & tba  |  CAG & TBA  ; 
 BAO <=  BAO & tba  |  CAO & TBA  ; 
 BBG <=  BBG & tbb  |  CAG & TBB  ; 
 BBO <=  BBO & tbb  |  CAO & TBB  ; 
 CAG <=  IAG & TCA  |  ABG & TCC  |  AAG & TCE  ; 
 OAG <=  IAG & TCA  |  ABG & TCC  |  AAG & TCE  ; 
 CAO <=  IAO & TCB  |  ABO & TCD  |  AAO & TCF  ; 
 OAO <=  IAO & TCB  |  ABO & TCD  |  AAO & TCF  ; 
 EAG <=  EBG & TEA  |  IGG & TEB  |  AAG & TEC  ; 
 TBA <= QIH ; 
 TBB <= QIG ; 
 TBC <= QJH ; 
 TBD <= QJG ; 
 BCG <=  BCG & tbc  |  CBG & TBC  ; 
 BCO <=  BCO & tbc  |  CBO & TBC  ; 
 BDG <=  BDG & tbd  |  CBG & TBD  ; 
 BDO <=  BDO & tbd  |  CBO & TBD  ; 
 CBG <=  IBG & TCG  |  ABG & TCI  |  AAG & TCK  ; 
 OBG <=  IBG & TCG  |  ABG & TCI  |  AAG & TCK  ; 
 CBO <=  IBO & TCH  |  ABO & TCJ  |  AAO & TCL  ; 
 OBO <=  IBO & TCH  |  ABO & TCJ  |  AAO & TCL  ; 
 QIH <= QIG ; 
 QJH <= QJG ; 
 OGA <=  IAQ  |  IAT  ; 
 QIG <=  IAQ  |  IAT  ; 
 OGB <=  IBQ  |  IBT  ; 
 QJG <=  IBQ  |  IBT  ; 
 BEG <=  BEG & tbe  |  CCG & TBE  ; 
 BEO <=  BEO & tbe  |  CCO & TBE  ; 
 BFG <=  BFG & tbf  |  CCG & TBF  ; 
 BFO <=  BFO & tbf  |  CCO & TBF  ; 
 CCG <=  ICG & TCM  |  ABG & TCO  |  AAG & TCQ  ; 
 OCG <=  ICG & TCM  |  ABG & TCO  |  AAG & TCQ  ; 
 CCO <=  ICO & TCN  |  ABO & TCP  |  AAO & TCR  ; 
 OCO <=  ICO & TCN  |  ABO & TCP  |  AAO & TCR  ; 
 BGG <=  BGG & tbg  |  CDG & TBG  ; 
 BGO <=  BGO & tbg  |  CDO & TBG  ; 
 BHG <=  BHG & tbh  |  CDG & TBH  ; 
 BHO <=  BHO & tbh  |  CDO & TBH  ; 
 CDG <=  IDG & TCS  |  ABG & TCU  |  AAG & TCW  ; 
 ODG <=  IDG & TCS  |  ABG & TCU  |  AAG & TCW  ; 
 CDO <=  IDO & TCT  |  ABO & TCV  |  AAO & TCX  ; 
 ODO <=  IDO & TCT  |  ABO & TCV  |  AAO & TCX  ; 
 WAH <= QCB ; 
 KBH <=  KAH & kap  |  kah & KAP  |  kah & kap  |  KAH & KAP  ;
 LBH <=  LAH & lap  |  lah & LAP  |  lah & lap  |  LAH & LAP  ;
 rah <=  rah & jah  |  RAH & JAH  |  QDA  ; 
 rch <=  rah & jah  |  RAH & JAH  |  QDA  ; 
 OEH <=  DAH & TDA  |  RAH & TDE  |  MAH & TDI  ; 
 PAH <=  DAH & TDA  |  RAH & TDE  |  MAH & TDI  ; 
 AAH <=  AAH & taa  |  IEH & TAA  ; 
 ACH <=  AAH & taa  |  IEH & TAA  ; 
 AEH <=  AAH & taa  |  IEH & TAA  ; 
 rap <=  rap & jap  |  RAP & JAP  |  QDB  ; 
 rcp <=  rap & jap  |  RAP & JAP  |  QDB  ; 
 OEP <=  DAP & TDB  |  RAP & TDF  |  MAP & TDJ  ; 
 PAP <=  DAP & TDB  |  RAP & TDF  |  MAP & TDJ  ; 
 AAP <=  AAP & tab  |  IEP & TAB  ; 
 ACP <=  AAP & tab  |  IEP & TAB  ; 
 AEP <=  AAP & tab  |  IEP & TAB  ; 
 TDA <= JCE ; 
 TDB <= JCE ; 
 TDC <= JCE ; 
 TDD <= JCE ; 
 ABH <=  ABH & tac  |  IFH & TAC  ; 
 ADH <=  ABH & tac  |  IFH & TAC  ; 
 AFH <=  ABH & tac  |  IFH & TAC  ; 
 rbh <=  rbh & jbh  |  RBH & JBH  |  QDC  ; 
 rdh <=  rbh & jbh  |  RBH & JBH  |  QDC  ; 
 OFH <=  DBH & TDC  |  RBH & TDG  |  MBH & TDK  ; 
 PBH <=  DBH & TDC  |  RBH & TDG  |  MBH & TDK  ; 
 ABP <=  ABP & tad  |  IFP & TAD  ; 
 ADP <=  ABP & tad  |  IFP & TAD  ; 
 AFP <=  ABP & tad  |  IFP & TAD  ; 
 rbp <=  rbp & jbp  |  RBP & JAP  |  QDD  ; 
 OFP <=  DBP & TDD  |  RBP & TDH  |  MBP & TDL  ; 
 PBP <=  DBP & TDD  |  RBP & TDH  |  MBP & TDL  ; 
 BAH <=  BAH & tba  |  CAH & TBA  ; 
 BAP <=  BAP & tba  |  CAP & TBA  ; 
 BBH <=  BBH & tbb  |  CAH & TBB  ; 
 BBP <=  BBP & tbb  |  CAP & TBB  ; 
 CAH <=  IAH & TCA  |  ABH & TCC  |  AAH & TCE  ; 
 OAH <=  IAH & TCA  |  ABH & TCC  |  AAH & TCE  ; 
 CAP <=  IAP & TCB  |  ABP & TCD  |  AAP & TCF  ; 
 OAP <=  IAP & TCB  |  ABP & TCD  |  AAP & TCF  ; 
 EAH <=  EBH & TEA  |  IGH & TEB  |  AAH & TEC  ; 
 BCH <=  BCH & tbc  |  CBH & TBC  ; 
 BCP <=  BCP & tbc  |  CBP & TBC  ; 
 BDH <=  BDH & tbd  |  CBH & TBD  ; 
 BDP <=  BDP & tbd  |  CBP & TBD  ; 
 CBH <=  IBH & TCG  |  ABH & TCI  |  AAH & TCK  ; 
 OBH <=  IBH & TCG  |  ABH & TCI  |  AAH & TCK  ; 
 CBP <=  IBP & TCH  |  ABP & TCJ  |  AAP & TCL  ; 
 OBP <=  IBP & TCH  |  ABP & TCJ  |  AAP & TCL  ; 
 QKH <= QKG ; 
 QLH <= QLG ; 
 OGC <=  ICQ  |  ICT  ; 
 QKG <=  ICQ  |  ICT  ; 
 OGD <=  IDQ  |  IDT  ; 
 QLG <=  IDQ  |  IDT  ; 
 BEH <=  BEH & tbe  |  CCH & TBE  ; 
 BEP <=  BEP & tbe  |  CCP & TBE  ; 
 BFH <=  BFH & tbf  |  CCH & TBF  ; 
 BFP <=  BFP & tbf  |  CCP & TBF  ; 
 CCH <=  ICH & TCM  |  ABH & TCO  |  AAH & TCQ  ; 
 OCH <=  ICH & TCM  |  ABH & TCO  |  AAH & TCQ  ; 
 CCP <=  ICP & TCN  |  ABP & TCP  |  AAP & TCR  ; 
 OCP <=  ICP & TCN  |  ABP & TCP  |  AAP & TCR  ; 
 TBE <= QKH ; 
 TBF <= QKG ; 
 TBH <= QLG ; 
 TBG <= QLH ; 
 BGH <=  BGH & tbg  |  CDH & TBG  ; 
 BGP <=  BGP & tbg  |  CDP & TBG  ; 
 BHH <=  BHH & tbh  |  CDH & TBH  ; 
 BHP <=  BHP & tbh  |  CDP & TBH  ; 
 CDH <=  IDH & TCS  |  ABH & TCU  |  AAH & TCW  ; 
 ODH <=  IDH & TCS  |  ABH & TCU  |  AAH & TCW  ; 
 CDP <=  IDP & TCT  |  ABP & TCV  |  AAP & TCX  ; 
 ODP <=  IDP & TCT  |  ABP & TCV  |  AAP & TCX  ; 
end
ram_4096x1 sinst_000(MAA,ACA,{FAA,FBA,FCA,FDA,FEA,FFA,FGA,FHA,FIA,FJA,FKA,FLA}, ZZI, WAA, IZZ); 
ram_4096x1 sinst_001(MAI,ACI,{FAA,FBA,FCA,FDA,FEA,FFA,FGA,FHA,FIA,FJA,FKA,FLA}, ZZI, WAA, IZZ); 
ram_4096x1 sinst_002(MBA,ADA,{FAA,FBA,FCA,FDA,FEA,FFA,FGA,FHA,FIA,FJA,FKA,FLA}, ZZI, WAA, IZZ); 
ram_4096x1 sinst_003(MBI,ADI,{FAA,FBA,FCA,FDA,FEA,FFA,FGA,FHA,FIA,FJA,FKA,FLA}, ZZI, WAA, IZZ); 
ram_4096x1 sinst_004(MBQ,KDA,{FMA,FMB,FMC,FMD,FME,FMF,FMG,FMH,FMI,FMJ,FMK,FML}, ZZI, WBA, IZZ); 
ram_4096x1 sinst_005(MAB,ACB,{FAB,FBB,FCB,FDB,FEB,FFB,FGB,FHB,FIB,FJB,FKB,FLB}, ZZI, WAB, IZZ); 
ram_4096x1 sinst_006(MAJ,ACJ,{FAB,FBB,FCB,FDB,FEB,FFB,FGB,FHB,FIB,FJB,FKB,FLB}, ZZI, WAB, IZZ); 
ram_4096x1 sinst_007(MBB,ADB,{FAB,FBB,FCB,FDB,FEB,FFB,FGB,FHB,FIB,FJB,FKB,FLB}, ZZI, WAB, IZZ); 
ram_4096x1 sinst_008(MBJ,ADJ,{FAB,FBB,FCB,FDB,FEB,FFB,FGB,FHB,FIB,FJB,FKB,FLB}, ZZI, WAB, IZZ); 
ram_4096x1 sinst_009(MAC,ACC,{FAC,FBC,FCC,FDC,FEC,FFC,FGC,FHC,FIC,FJC,FKC,FLC}, ZZI, WAC, IZZ); 
ram_4096x1 sinst_010(MAK,ACK,{FAC,FBC,FCC,FDC,FEC,FFC,FGC,FHC,FIC,FJC,FKC,FLC}, ZZI, WAC, IZZ); 
ram_4096x1 sinst_011(MBC,ADC,{FAC,FBC,FCC,FDC,FEC,FFC,FGC,FHC,FIC,FJC,FKC,FLC}, ZZI, WAC, IZZ); 
ram_4096x1 sinst_012(MBK,ADK,{FAC,FBC,FCC,FDC,FEC,FFC,FGC,FHC,FIC,FJC,FKC,FLC}, ZZI, WAC, IZZ); 
ram_4096x1 sinst_013(MAD,ACD,{FAD,FBD,FCD,FDD,FED,FFD,FGD,FHD,FID,FJD,FKD,FLD}, ZZI, WAD, IZZ); 
ram_4096x1 sinst_014(MAL,ACL,{FAD,FBD,FCD,FDD,FED,FFD,FGD,FHD,FID,FJD,FKD,FLD}, ZZI, WAD, IZZ); 
ram_4096x1 sinst_015(MBD,ADD,{FAD,FBD,FCD,FDD,FED,FFD,FGD,FHD,FID,FJD,FKD,FLD}, ZZI, WAD, IZZ); 
ram_4096x1 sinst_016(MBL,ADL,{FAD,FBD,FCD,FDD,FED,FFD,FGD,FHD,FID,FJD,FKD,FLD}, ZZI, WAD, IZZ); 
ram_4096x1 sinst_017(MAE,ACE,{FAE,FBE,FCE,FDE,FEE,FFE,FGE,FHE,FIE,FJE,FKE,FLE}, ZZI, WAE, IZZ); 
ram_4096x1 sinst_018(MAM,ACM,{FAE,FBE,FCE,FDE,FEE,FFE,FGE,FHE,FIE,FJE,FKE,FLE}, ZZI, WAE, IZZ); 
ram_4096x1 sinst_019(MBE,ADE,{FAE,FBE,FCE,FDE,FEE,FFE,FGE,FHE,FIE,FJE,FKE,FLE}, ZZI, WAE, IZZ); 
ram_4096x1 sinst_020(MBM,ADM,{FAE,FBE,FCE,FDE,FEE,FFE,FGE,FHE,FIE,FJE,FKE,FLE}, ZZI, WAE, IZZ); 
ram_4096x1 sinst_021(MAF,ACF,{FAF,FBF,FCF,FDF,FEF,FFF,FGF,FHF,FIF,FJF,FKF,FLF}, ZZI, WAF, IZZ); 
ram_4096x1 sinst_022(MAN,ACN,{FAF,FBF,FCF,FDF,FEF,FFF,FGF,FHF,FIF,FJF,FKF,FLF}, ZZI, WAF, IZZ); 
ram_4096x1 sinst_023(MBF,ADF,{FAF,FBF,FCF,FDF,FEF,FFF,FGF,FHF,FIF,FJF,FKF,FLF}, ZZI, WAF, IZZ); 
ram_4096x1 sinst_024(MBN,ADN,{FAF,FBF,FCF,FDF,FEF,FFF,FGF,FHF,FIF,FJF,FKF,FLF}, ZZI, WAF, IZZ); 
ram_4096x1 sinst_025(MAG,ACG,{FAG,FBG,FCG,FDG,FEG,FFG,FGG,FHG,FIG,FJG,FKG,FLG}, ZZI, WAG, IZZ); 
ram_4096x1 sinst_026(MAO,ACO,{FAG,FBG,FCG,FDG,FEG,FFG,FGG,FHG,FIG,FJG,FKG,FLG}, ZZI, WAG, IZZ); 
ram_4096x1 sinst_027(MBG,ADG,{FAG,FBG,FCG,FDG,FEG,FFG,FGG,FHG,FIG,FJG,FKG,FLG}, ZZI, WAG, IZZ); 
ram_4096x1 sinst_028(MBO,ADO,{FAG,FBG,FCG,FDG,FEG,FFG,FGG,FHG,FIG,FJG,FKG,FLG}, ZZI, WAG, IZZ); 
ram_4096x1 sinst_029(MAH,ACH,{FAH,FBH,FCH,FDH,FEH,FFH,FGH,FHH,FIH,FJH,FKH,FLH}, ZZI, WAH, IZZ); 
ram_4096x1 sinst_030(MAP,ACP,{FAH,FBH,FCH,FDH,FEH,FFH,FGH,FHH,FIH,FJH,FKH,FLH}, ZZI, WAH, IZZ); 
ram_4096x1 sinst_031(MBH,ADH,{FAH,FBH,FCH,FDH,FEH,FFH,FGH,FHH,FIH,FJH,FKH,FLH}, ZZI, WAH, IZZ); 
ram_4096x1 sinst_032(MBP,ADP,{FAH,FBH,FCH,FDH,FEH,FFH,FGH,FHH,FIH,FJH,FKH,FLH}, ZZI, WAH, IZZ); 
endmodule;
