module ma( IZZ,
 IAA, 
 IAB, 
 IAC, 
 IAD, 
 IAE, 
 IAF, 
 IAG, 
 IAH, 
 IAI, 
 IAJ, 
 IAK, 
 IAL, 
 IAM, 
 IAN, 
 IAO, 
 IAP, 
 IBA, 
 IBB, 
 IBC, 
 IBD, 
 IBE, 
 IBF, 
 IBG, 
 IBH, 
 IBI, 
 IBJ, 
 IBK, 
 IBL, 
 IBM, 
 IBN, 
 IBO, 
 IBP, 
 ICA, 
 ICB, 
 ICC, 
 ICD, 
 ICE, 
 ICF, 
 ICG, 
 ICH, 
 ICI, 
 ICJ, 
 ICK, 
 ICL, 
 ICM, 
 ICN, 
 ICO, 
 ICP, 
 IDA, 
 IDB, 
 IDC, 
 IDD, 
 IDE, 
 IDF, 
 IDG, 
 IDH, 
 IDI, 
 IDJ, 
 IDK, 
 IDL, 
 IDM, 
 IDN, 
 IDO, 
 IDP, 
 IEA, 
 IEB, 
 IEC, 
 IED, 
 IEE, 
 IEF, 
 IEG, 
 IEH, 
 IEI, 
 IEJ, 
 IEK, 
 IEL, 
 IEM, 
 IEN, 
 IEO, 
 IEP, 
 IEQ, 
 IER, 
 IES, 
 IET, 
 IEU, 
 IEV, 
 IEW, 
 IEX, 
 IEY, 
 IEZ, 
 IFA, 
 IFB, 
 IFC, 
 IFD, 
 IFE, 
 IFFF , 
 IFG, 
 IFH, 
 IFI, 
 IFJ, 
 IFK, 
 IFL, 
 IFM, 
 IFN, 
 IFO, 
 IFP, 
 IGA, 
 IHA, 
 IKA, 
 IMM, 
 IMR, 
 IMS, 
 IRA, 
 ISA, 
 ITA, 
 OAA, 
 OAB, 
 OAC, 
 OAD, 
 OAE, 
 OAF, 
 OAG, 
 OAH, 
 OAI, 
 OAJ, 
 OAK, 
 OAL, 
 OAM, 
 OAN, 
 OAO, 
 OAP, 
 OBA, 
 OBB, 
 OBC, 
 OBD, 
 OBE, 
 OBF, 
 OBG, 
 OBH, 
 OBI, 
 OBJ, 
 OBK, 
 OBL, 
 OBM, 
 OBN, 
 OBO, 
 OBP, 
 OCG, 
 OCH, 
 OCI, 
 OCJ, 
 OCK, 
 OCL, 
 OCM, 
 OCN, 
 OCO, 
 OCP, 
 ODA, 
 ODB, 
 ODC, 
 ODD, 
 ODE, 
 ODF, 
 ODG, 
 ODH, 
 ODI, 
 ODJ, 
 ODK, 
 ODL, 
 ODM, 
 ODN, 
 ODO, 
 ODP, 
 OEA, 
 OEB, 
 OEC, 
 OED, 
 OEE, 
 OEF, 
 OEG, 
 OEH, 
 OEI, 
 OEJ, 
 OEK, 
 OEL, 
 OEM, 
 OEN, 
 OEO, 
 OEP, 
 OFG, 
 OFH, 
 OFI, 
 OFJ, 
 OFK, 
 OFL, 
 OFM, 
 OFN, 
 OFO, 
 OFP, 
 OGA, 
 OGB, 
 OGC, 
 OGD, 
 OGE, 
 OGF, 
 OGG, 
 OGH, 
 OGI, 
 OGJ, 
 OGK, 
 OGL, 
 OGM, 
 OGN, 
 OGO, 
 OGP, 
 OHA, 
 OHB, 
 OHC, 
 OHD, 
 OHE, 
 OHF, 
 OHG, 
 OHH, 
 OHI, 
 OHJ, 
 OHK, 
 OIH, 
 OII, 
 OIJ, 
 OKA, 
 OKB, 
 OKC, 
 OKD, 
 OKE, 
 OKF, 
 OLD, 
 OMA, 
 OMB, 
 ONB, 
 OPK, 
 OPM, 
 OPO, 
 OPQ, 
 OPR, 
 OQJ, 
 OQK, 
 OQM, 
 OQO, 
OQQ ); 
    
 input IZZ; 
 input IAA; 
 input IAB; 
 input IAC; 
 input IAD; 
 input IAE; 
 input IAF; 
 input IAG; 
 input IAH; 
 input IAI; 
 input IAJ; 
 input IAK; 
 input IAL; 
 input IAM; 
 input IAN; 
 input IAO; 
 input IAP; 
 input IBA; 
 input IBB; 
 input IBC; 
 input IBD; 
 input IBE; 
 input IBF; 
 input IBG; 
 input IBH; 
 input IBI; 
 input IBJ; 
 input IBK; 
 input IBL; 
 input IBM; 
 input IBN; 
 input IBO; 
 input IBP; 
 input ICA; 
 input ICB; 
 input ICC; 
 input ICD; 
 input ICE; 
 input ICF; 
 input ICG; 
 input ICH; 
 input ICI; 
 input ICJ; 
 input ICK; 
 input ICL; 
 input ICM; 
 input ICN; 
 input ICO; 
 input ICP; 
 input IDA; 
 input IDB; 
 input IDC; 
 input IDD; 
 input IDE; 
 input IDF; 
 input IDG; 
 input IDH; 
 input IDI; 
 input IDJ; 
 input IDK; 
 input IDL; 
 input IDM; 
 input IDN; 
 input IDO; 
 input IDP; 
 input IEA; 
 input IEB; 
 input IEC; 
 input IED; 
 input IEE; 
 input IEF; 
 input IEG; 
 input IEH; 
 input IEI; 
 input IEJ; 
 input IEK; 
 input IEL; 
 input IEM; 
 input IEN; 
 input IEO; 
 input IEP; 
 input IEQ; 
 input IER; 
 input IES; 
 input IET; 
 input IEU; 
 input IEV; 
 input IEW; 
 input IEX; 
 input IEY; 
 input IEZ; 
 input IFA; 
 input IFB; 
 input IFC; 
 input IFD; 
 input IFE; 
 input IFFF ; 
 input IFG; 
 input IFH; 
 input IFI; 
 input IFJ; 
 input IFK; 
 input IFL; 
 input IFM; 
 input IFN; 
 input IFO; 
 input IFP; 
 input IGA; 
 input IHA; 
 input IKA; 
 input IMM; 
 input IMR; 
 input IMS; 
 input IRA; 
 input ISA; 
 input ITA; 
 output OAA; 
 output OAB; 
 output OAC; 
 output OAD; 
 output OAE; 
 output OAF; 
 output OAG; 
 output OAH; 
 output OAI; 
 output OAJ; 
 output OAK; 
 output OAL; 
 output OAM; 
 output OAN; 
 output OAO; 
 output OAP; 
 output OBA; 
 output OBB; 
 output OBC; 
 output OBD; 
 output OBE; 
 output OBF; 
 output OBG; 
 output OBH; 
 output OBI; 
 output OBJ; 
 output OBK; 
 output OBL; 
 output OBM; 
 output OBN; 
 output OBO; 
 output OBP; 
 output OCG; 
 output OCH; 
 output OCI; 
 output OCJ; 
 output OCK; 
 output OCL; 
 output OCM; 
 output OCN; 
 output OCO; 
 output OCP; 
 output ODA; 
 output ODB; 
 output ODC; 
 output ODD; 
 output ODE; 
 output ODF; 
 output ODG; 
 output ODH; 
 output ODI; 
 output ODJ; 
 output ODK; 
 output ODL; 
 output ODM; 
 output ODN; 
 output ODO; 
 output ODP; 
 output OEA; 
 output OEB; 
 output OEC; 
 output OED; 
 output OEE; 
 output OEF; 
 output OEG; 
 output OEH; 
 output OEI; 
 output OEJ; 
 output OEK; 
 output OEL; 
 output OEM; 
 output OEN; 
 output OEO; 
 output OEP; 
 output OFG; 
 output OFH; 
 output OFI; 
 output OFJ; 
 output OFK; 
 output OFL; 
 output OFM; 
 output OFN; 
 output OFO; 
 output OFP; 
 output OGA; 
 output OGB; 
 output OGC; 
 output OGD; 
 output OGE; 
 output OGF; 
 output OGG; 
 output OGH; 
 output OGI; 
 output OGJ; 
 output OGK; 
 output OGL; 
 output OGM; 
 output OGN; 
 output OGO; 
 output OGP; 
 output OHA; 
 output OHB; 
 output OHC; 
 output OHD; 
 output OHE; 
 output OHF; 
 output OHG; 
 output OHH; 
 output OHI; 
 output OHJ; 
 output OHK; 
 output OIH; 
 output OII; 
 output OIJ; 
 output OKA; 
 output OKB; 
 output OKC; 
 output OKD; 
 output OKE; 
 output OKF; 
 output OLD; 
 output OMA; 
 output OMB; 
 output ONB; 
 output OPK; 
 output OPM; 
 output OPO; 
 output OPQ; 
 output OPR; 
 output OQJ; 
 output OQK; 
 output OQM; 
 output OQO; 
 output OQQ; 
  
  
reg  AAA ;
reg  AAB ;
reg  AAC ;
reg  AAD ;
reg  AAE ;
reg  AAF ;
reg  AAG ;
reg  AAH ;
reg  AAI ;
reg  AAJ ;
reg  AAK ;
reg  AAL ;
reg  AAM ;
reg  AAN ;
reg  AAO ;
reg  AAP ;
reg  BAA ;
reg  BAB ;
reg  BAC ;
reg  BAD ;
reg  BAE ;
reg  BAF ;
reg  BAG ;
reg  BAH ;
reg  BAI ;
reg  BAJ ;
reg  BAK ;
reg  BAL ;
reg  BAM ;
reg  BAN ;
reg  BAO ;
reg  BAP ;
reg  bba ;
reg  bbb ;
reg  bbc ;
reg  bbd ;
reg  bbe ;
reg  bbf ;
reg  bbg ;
reg  bbh ;
reg  bbi ;
reg  bbj ;
reg  bbk ;
reg  bbl ;
reg  bbm ;
reg  bbn ;
reg  bbo ;
reg  bbp ;
reg  BCA ;
reg  BCB ;
reg  BCC ;
reg  BCD ;
reg  BCE ;
reg  BCF ;
reg  BCG ;
reg  BCH ;
reg  BCI ;
reg  BCJ ;
reg  BCK ;
reg  BCL ;
reg  BCM ;
reg  BCN ;
reg  BCO ;
reg  BCP ;
reg  BDA ;
reg  BDB ;
reg  BDC ;
reg  BDD ;
reg  BDE ;
reg  BDF ;
reg  BDG ;
reg  BDH ;
reg  BDI ;
reg  BDJ ;
reg  BDK ;
reg  BDL ;
reg  BDM ;
reg  BDN ;
reg  BDO ;
reg  BDP ;
reg  BEA ;
reg  BEB ;
reg  BEC ;
reg  BED ;
reg  BEE ;
reg  BEF ;
reg  BEG ;
reg  BEH ;
reg  BEI ;
reg  BEJ ;
reg  BEK ;
reg  BEL ;
reg  BEM ;
reg  BEN ;
reg  BEO ;
reg  BEP ;
reg  caa ;
reg  CAB ;
reg  CAC ;
reg  CAD ;
reg  CAE ;
reg  CAF ;
reg  CAG ;
reg  CAH ;
reg  CAI ;
reg  CAJ ;
reg  CAK ;
reg  CAL ;
reg  CAM ;
reg  CAN ;
reg  CAO ;
reg  CAP ;
reg  CBA ;
reg  CBB ;
reg  CBC ;
reg  CBD ;
reg  CBE ;
reg  CBF ;
reg  CBG ;
reg  CBH ;
reg  CBI ;
reg  CBJ ;
reg  CBK ;
reg  CBL ;
reg  CBM ;
reg  CBN ;
reg  CBO ;
reg  CBP ;
reg  CCA ;
reg  CCB ;
reg  CCC ;
reg  CCD ;
reg  CCE ;
reg  CCF ;
reg  CCG ;
reg  CCH ;
reg  CCI ;
reg  CCJ ;
reg  CCK ;
reg  CCL ;
reg  CCM ;
reg  CCN ;
reg  CCO ;
reg  CCP ;
reg  cda ;
reg  CDB ;
reg  CDC ;
reg  CDD ;
reg  CDE ;
reg  CDF ;
reg  CDG ;
reg  CDH ;
reg  CDI ;
reg  CDJ ;
reg  CDK ;
reg  CDL ;
reg  CDM ;
reg  CDN ;
reg  CDO ;
reg  CDP ;
reg  CEA ;
reg  CEB ;
reg  CEC ;
reg  CED ;
reg  CEE ;
reg  CEF ;
reg  CEG ;
reg  CEH ;
reg  CEI ;
reg  CEJ ;
reg  CEK ;
reg  CEL ;
reg  CEM ;
reg  CEN ;
reg  CEO ;
reg  CEP ;
reg  CFA ;
reg  CFB ;
reg  CFC ;
reg  CFD ;
reg  CFE ;
reg  CFF ;
reg  CFG ;
reg  CFH ;
reg  CFI ;
reg  CFJ ;
reg  CFK ;
reg  CFL ;
reg  CFM ;
reg  DAF ;
reg  DAG ;
reg  DAH ;
reg  DAI ;
reg  DAJ ;
reg  DAK ;
reg  DAL ;
reg  DAM ;
reg  DAN ;
reg  DAO ;
reg  DAP ;
reg  DBA ;
reg  dbb ;
reg  dbc ;
reg  dbd ;
reg  dbe ;
reg  dbf ;
reg  dbg ;
reg  dbh ;
reg  dbi ;
reg  DBN ;
reg  DBO ;
reg  DBP ;
reg  DCA ;
reg  DCB ;
reg  DCC ;
reg  DCD ;
reg  DCE ;
reg  DCF ;
reg  DCG ;
reg  DCH ;
reg  DCI ;
reg  DCJ ;
reg  DCK ;
reg  DCL ;
reg  DCM ;
reg  DDA ;
reg  DDB ;
reg  DDC ;
reg  DDD ;
reg  DDE ;
reg  ddf ;
reg  ddg ;
reg  ddh ;
reg  ddi ;
reg  ddj ;
reg  ddk ;
reg  ddl ;
reg  ddm ;
reg  DEB ;
reg  DEC ;
reg  DED ;
reg  DEE ;
reg  DEF ;
reg  DEG ;
reg  DEH ;
reg  DEI ;
reg  DEJ ;
reg  DEK ;
reg  DEL ;
reg  DEM ;
reg  den ;
reg  deo ;
reg  dep ;
reg  dfa ;
reg  dfb ;
reg  dfc ;
reg  dfd ;
reg  dfe ;
reg  DGA ;
reg  DGB ;
reg  DGC ;
reg  DGD ;
reg  DGE ;
reg  dgf ;
reg  dgg ;
reg  dgh ;
reg  dgi ;
reg  DGK ;
reg  DGL ;
reg  DGM ;
reg  DGN ;
reg  DGO ;
reg  DGP ;
reg  DHA ;
reg  dhb ;
reg  dhc ;
reg  dhd ;
reg  dhe ;
reg  DHG ;
reg  DHH ;
reg  DHI ;
reg  DHJ ;
reg  DHK ;
reg  DHL ;
reg  DHM ;
reg  dhn ;
reg  dho ;
reg  dhp ;
reg  dia ;
reg  DIC ;
reg  DID ;
reg  DIE ;
reg  DIF ;
reg  DIG ;
reg  DIH ;
reg  DII ;
reg  DIJ ;
reg  DIK ;
reg  DIL ;
reg  DIM ;
reg  DIN ;
reg  DIO ;
reg  DIP ;
reg  FAA ;
reg  FAB ;
reg  FAC ;
reg  FAD ;
reg  FAE ;
reg  FAF ;
reg  FAG ;
reg  FAH ;
reg  FAI ;
reg  FAJ ;
reg  FAK ;
reg  FAL ;
reg  FAM ;
reg  FAN ;
reg  fba ;
reg  fbb ;
reg  fbc ;
reg  fbd ;
reg  fbe ;
reg  fbf ;
reg  fbg ;
reg  fbh ;
reg  fbi ;
reg  fbj ;
reg  fbk ;
reg  fbl ;
reg  fbm ;
reg  fbn ;
reg  FCA ;
reg  FCB ;
reg  FCC ;
reg  FCD ;
reg  FCE ;
reg  FCF ;
reg  FCG ;
reg  FCH ;
reg  FCI ;
reg  FCJ ;
reg  FCK ;
reg  FCL ;
reg  FCM ;
reg  FCN ;
reg  FCO ;
reg  fdb ;
reg  fdc ;
reg  fdd ;
reg  fde ;
reg  fdf ;
reg  fdg ;
reg  fdh ;
reg  fdi ;
reg  fdj ;
reg  fdk ;
reg  fdl ;
reg  fdm ;
reg  fdn ;
reg  fdo ;
reg  FEA ;
reg  FEB ;
reg  FEC ;
reg  FED ;
reg  FEE ;
reg  FEF ;
reg  FEG ;
reg  FEH ;
reg  FEI ;
reg  FEJ ;
reg  FEK ;
reg  FEL ;
reg  FEM ;
reg  FEN ;
reg  FEO ;
reg  FEP ;
reg  ffc ;
reg  ffd ;
reg  ffe ;
reg  fff ;
reg  ffg ;
reg  ffh ;
reg  ffi ;
reg  ffj ;
reg  ffk ;
reg  ffl ;
reg  ffm ;
reg  ffn ;
reg  ffo ;
reg  ffp ;
reg  FGA ;
reg  FGB ;
reg  FGC ;
reg  FGD ;
reg  FGE ;
reg  FGF ;
reg  FGG ;
reg  FGH ;
reg  FGI ;
reg  FGJ ;
reg  FGK ;
reg  FGL ;
reg  FGM ;
reg  FGN ;
reg  FGO ;
reg  fha ;
reg  fhb ;
reg  fhc ;
reg  fhd ;
reg  fhe ;
reg  fhf ;
reg  fhg ;
reg  fhh ;
reg  fhi ;
reg  fhj ;
reg  fhk ;
reg  fhl ;
reg  fhm ;
reg  fhn ;
reg  fho ;
reg  FIA ;
reg  FIB ;
reg  FIC ;
reg  FID ;
reg  FIE ;
reg  FIF ;
reg  FIG ;
reg  FIH ;
reg  FII ;
reg  FIJ ;
reg  FIK ;
reg  FIL ;
reg  FIM ;
reg  FIN ;
reg  FIO ;
reg  FIP ;
reg  fjb ;
reg  fjc ;
reg  fjd ;
reg  fje ;
reg  fjf ;
reg  fjg ;
reg  fjh ;
reg  fji ;
reg  fjj ;
reg  fjk ;
reg  fjl ;
reg  fjm ;
reg  fjn ;
reg  fjo ;
reg  fjp ;
reg  FKA ;
reg  FKB ;
reg  FKC ;
reg  FKD ;
reg  FKE ;
reg  FKF ;
reg  FKG ;
reg  FKH ;
reg  FKI ;
reg  FKJ ;
reg  FKK ;
reg  FKL ;
reg  FKM ;
reg  FKN ;
reg  FKO ;
reg  FKP ;
reg  FKQ ;
reg  flc ;
reg  fld ;
reg  fle ;
reg  flf ;
reg  flg ;
reg  flh ;
reg  fli ;
reg  flj ;
reg  flk ;
reg  fll ;
reg  flm ;
reg  fln ;
reg  flo ;
reg  flp ;
reg  flq ;
reg  FMA ;
reg  FMB ;
reg  FMC ;
reg  FMD ;
reg  FME ;
reg  FMF ;
reg  FMG ;
reg  FMH ;
reg  FMI ;
reg  FMJ ;
reg  FMK ;
reg  FML ;
reg  FMM ;
reg  FMN ;
reg  FMO ;
reg  FMP ;
reg  fna ;
reg  fnb ;
reg  fnc ;
reg  fnd ;
reg  fne ;
reg  fnf ;
reg  fng ;
reg  fnh ;
reg  fni ;
reg  fnj ;
reg  fnk ;
reg  fnl ;
reg  fnm ;
reg  fnn ;
reg  fno ;
reg  fnp ;
reg  FOA ;
reg  FOB ;
reg  FOC ;
reg  FOD ;
reg  FOE ;
reg  FOF ;
reg  FOG ;
reg  FOH ;
reg  FOI ;
reg  FOJ ;
reg  FOK ;
reg  FOL ;
reg  FOM ;
reg  FON ;
reg  FOO ;
reg  FOP ;
reg  FOQ ;
reg  fpb ;
reg  fpc ;
reg  fpd ;
reg  fpe ;
reg  fpf ;
reg  fpg ;
reg  fph ;
reg  fpi ;
reg  fpj ;
reg  fpk ;
reg  fpl ;
reg  fpm ;
reg  fpn ;
reg  fpo ;
reg  fpp ;
reg  fpq ;
reg  FQA ;
reg  FQB ;
reg  FQC ;
reg  FQD ;
reg  FQE ;
reg  FQF ;
reg  FQG ;
reg  FQH ;
reg  FQI ;
reg  FQJ ;
reg  FQK ;
reg  FQL ;
reg  FQM ;
reg  FQN ;
reg  FQO ;
reg  FQP ;
reg  HAA ;
reg  HAB ;
reg  hba ;
reg  hbb ;
reg  HCA ;
reg  HCB ;
reg  HCC ;
reg  HCD ;
reg  HCE ;
reg  hda ;
reg  hdb ;
reg  hdc ;
reg  hdd ;
reg  hde ;
reg  HEA ;
reg  HEB ;
reg  HEC ;
reg  HED ;
reg  HEE ;
reg  HEF ;
reg  HEG ;
reg  hfa ;
reg  hfb ;
reg  hfc ;
reg  hfd ;
reg  hfe ;
reg  hff ;
reg  HGA ;
reg  HGB ;
reg  HGC ;
reg  HGD ;
reg  HGE ;
reg  HGF ;
reg  HGG ;
reg  hha ;
reg  hhb ;
reg  hhc ;
reg  hhd ;
reg  hhe ;
reg  hhf ;
reg  hhg ;
reg  HIA ;
reg  HIB ;
reg  HIC ;
reg  HID ;
reg  HIE ;
reg  HIF ;
reg  HIG ;
reg  HIH ;
reg  hja ;
reg  hjb ;
reg  hjc ;
reg  hjd ;
reg  hje ;
reg  hjf ;
reg  HKA ;
reg  HKB ;
reg  HKC ;
reg  HKD ;
reg  HKE ;
reg  HKF ;
reg  HKG ;
reg  HKH ;
reg  hla ;
reg  hlb ;
reg  hlc ;
reg  hld ;
reg  hle ;
reg  hlf ;
reg  hlg ;
reg  HMA ;
reg  HMB ;
reg  HMC ;
reg  HMD ;
reg  HME ;
reg  HMF ;
reg  HMG ;
reg  hna ;
reg  hnb ;
reg  hnc ;
reg  hnd ;
reg  hne ;
reg  hnf ;
reg  hng ;
reg  HOA ;
reg  HOB ;
reg  HOC ;
reg  HOD ;
reg  HOE ;
reg  HOF ;
reg  HOG ;
reg  hpa ;
reg  hpb ;
reg  hpc ;
reg  hpd ;
reg  hpe ;
reg  hpf ;
reg  hpg ;
reg  HQA ;
reg  HQB ;
reg  HQC ;
reg  HQD ;
reg  HQE ;
reg  HQF ;
reg  HQG ;
reg  HQH ;
reg  HQI ;
reg  KCA ;
reg  KCB ;
reg  kda ;
reg  KEA ;
reg  KEB ;
reg  kfa ;
reg  kfb ;
reg  KGA ;
reg  KGB ;
reg  KGC ;
reg  kha ;
reg  khb ;
reg  khc ;
reg  KIA ;
reg  KIB ;
reg  KIC ;
reg  kja ;
reg  kjb ;
reg  kjc ;
reg  KKA ;
reg  KKB ;
reg  KKC ;
reg  KKD ;
reg  KKE ;
reg  kla ;
reg  klb ;
reg  klc ;
reg  KMA ;
reg  KMB ;
reg  KMC ;
reg  KMD ;
reg  kna ;
reg  knb ;
reg  knc ;
reg  KOA ;
reg  KOB ;
reg  KOC ;
reg  KOD ;
reg  kpa ;
reg  kpb ;
reg  kpc ;
reg  KQA ;
reg  KQB ;
reg  KQC ;
reg  KQD ;
reg  mfa ;
reg  MGA ;
reg  MGB ;
reg  mha ;
reg  MIA ;
reg  mja ;
reg  MKA ;
reg  MKB ;
reg  mla ;
reg  mlb ;
reg  MMA ;
reg  MMB ;
reg  MMC ;
reg  mna ;
reg  MOA ;
reg  MOB ;
reg  MOC ;
reg  mpa ;
reg  MQA ;
reg  MQB ;
reg  MQC ;
reg  OAA ;
reg  OAB ;
reg  OAC ;
reg  OAD ;
reg  OAE ;
reg  OAF ;
reg  OAG ;
reg  OAH ;
reg  OAI ;
reg  OAJ ;
reg  OAK ;
reg  OAL ;
reg  OAM ;
reg  OAN ;
reg  OAO ;
reg  OAP ;
reg  OBA ;
reg  OBB ;
reg  OBC ;
reg  OBD ;
reg  OBE ;
reg  OBF ;
reg  OBG ;
reg  OBH ;
reg  OBI ;
reg  OBJ ;
reg  OBK ;
reg  OBL ;
reg  OBM ;
reg  OBN ;
reg  OBO ;
reg  OBP ;
reg  OCG ;
reg  OCH ;
reg  OCI ;
reg  OCJ ;
reg  OCK ;
reg  OCL ;
reg  OCM ;
reg  OCN ;
reg  OCO ;
reg  OCP ;
reg  ODA ;
reg  ODB ;
reg  ODC ;
reg  ODD ;
reg  ODE ;
reg  ODF ;
reg  ODG ;
reg  ODH ;
reg  ODI ;
reg  ODJ ;
reg  ODK ;
reg  ODL ;
reg  ODM ;
reg  ODN ;
reg  ODO ;
reg  ODP ;
reg  OEA ;
reg  OEB ;
reg  OEC ;
reg  OED ;
reg  OEE ;
reg  OEF ;
reg  OEG ;
reg  OEH ;
reg  OEI ;
reg  OEJ ;
reg  OEK ;
reg  OEL ;
reg  OEM ;
reg  OEN ;
reg  OEO ;
reg  OEP ;
reg  OFG ;
reg  OFH ;
reg  OFI ;
reg  OFJ ;
reg  OFK ;
reg  OFL ;
reg  OFM ;
reg  OFN ;
reg  OFO ;
reg  OFP ;
reg  oga ;
reg  ogb ;
reg  ogc ;
reg  ogd ;
reg  oge ;
reg  ogf ;
reg  ogg ;
reg  ogh ;
reg  ogi ;
reg  ogj ;
reg  ogk ;
reg  ogl ;
reg  ogm ;
reg  ogn ;
reg  ogo ;
reg  ogp ;
reg  oha ;
reg  ohb ;
reg  ohc ;
reg  ohd ;
reg  ohe ;
reg  ohf ;
reg  ohg ;
reg  OHH ;
reg  OHI ;
reg  OHJ ;
reg  OHK ;
reg  oih ;
reg  oii ;
reg  oij ;
reg  oka ;
reg  okb ;
reg  okc ;
reg  OKD ;
reg  OKE ;
reg  OKF ;
reg  old ;
reg  oma ;
reg  OMB ;
reg  onb ;
reg  OPK ;
reg  OPM ;
reg  OPO ;
reg  OPQ ;
reg  OPR ;
reg  oqj ;
reg  oqk ;
reg  oqm ;
reg  oqo ;
reg  oqq ;
reg  QAA ;
reg  QAB ;
reg  QAC ;
reg  QAD ;
reg  QAE ;
reg  QAF ;
reg  QAG ;
reg  QAH ;
reg  QAI ;
reg  QGA ;
reg  QHA ;
reg  QKA ;
reg  QMM ;
reg  QMR ;
reg  QMS ;
reg  QRA ;
reg  QSA ;
reg  QTA ;
reg  TAM ;
reg  TAR ;
reg  TAS ;
reg  TGA ;
reg  tgb ;
reg  TGC ;
reg  tgd ;
reg  TGE ;
reg  tgf ;
reg  THA ;
reg  thb ;
reg  THC ;
reg  thd ;
reg  THE ;
reg  thf ;
reg  TKA ;
reg  tkb ;
reg  TKC ;
reg  tkd ;
reg  TKE ;
reg  tkf ;
reg  TRA ;
reg  TRB ;
reg  trc ;
reg  TSA ;
reg  tsb ;
reg  TSC ;
reg  tsd ;
reg  TSE ;
reg  tsf ;
reg  TTA ;
reg  ttb ;
reg  TTC ;
reg  ttd ;
reg  TTE ;
reg  ttf ;
wire  aaa ;
wire  aab ;
wire  aac ;
wire  aad ;
wire  aae ;
wire  aaf ;
wire  aag ;
wire  aah ;
wire  aai ;
wire  aaj ;
wire  aak ;
wire  aal ;
wire  aam ;
wire  aan ;
wire  aao ;
wire  aap ;
wire  baa ;
wire  bab ;
wire  bac ;
wire  bad ;
wire  bae ;
wire  baf ;
wire  bag ;
wire  bah ;
wire  bai ;
wire  baj ;
wire  bak ;
wire  bal ;
wire  bam ;
wire  ban ;
wire  bao ;
wire  bap ;
wire  BBA ;
wire  BBB ;
wire  BBC ;
wire  BBD ;
wire  BBE ;
wire  BBF ;
wire  BBG ;
wire  BBH ;
wire  BBI ;
wire  BBJ ;
wire  BBK ;
wire  BBL ;
wire  BBM ;
wire  BBN ;
wire  BBO ;
wire  BBP ;
wire  bca ;
wire  bcb ;
wire  bcc ;
wire  bcd ;
wire  bce ;
wire  bcf ;
wire  bcg ;
wire  bch ;
wire  bci ;
wire  bcj ;
wire  bck ;
wire  bcl ;
wire  bcm ;
wire  bcn ;
wire  bco ;
wire  bcp ;
wire  bda ;
wire  bdb ;
wire  bdc ;
wire  bdd ;
wire  bde ;
wire  bdf ;
wire  bdg ;
wire  bdh ;
wire  bdi ;
wire  bdj ;
wire  bdk ;
wire  bdl ;
wire  bdm ;
wire  bdn ;
wire  bdo ;
wire  bdp ;
wire  bea ;
wire  beb ;
wire  bec ;
wire  bed ;
wire  bee ;
wire  bef ;
wire  beg ;
wire  beh ;
wire  bei ;
wire  bej ;
wire  bek ;
wire  bel ;
wire  bem ;
wire  ben ;
wire  beo ;
wire  bep ;
wire  CAA ;
wire  cab ;
wire  cac ;
wire  cad ;
wire  cae ;
wire  caf ;
wire  cag ;
wire  cah ;
wire  cai ;
wire  caj ;
wire  cak ;
wire  cal ;
wire  cam ;
wire  can ;
wire  cao ;
wire  cap ;
wire  cba ;
wire  cbb ;
wire  cbc ;
wire  cbd ;
wire  cbe ;
wire  cbf ;
wire  cbg ;
wire  cbh ;
wire  cbi ;
wire  cbj ;
wire  cbk ;
wire  cbl ;
wire  cbm ;
wire  cbn ;
wire  cbo ;
wire  cbp ;
wire  cca ;
wire  ccb ;
wire  ccc ;
wire  ccd ;
wire  cce ;
wire  ccf ;
wire  ccg ;
wire  cch ;
wire  cci ;
wire  ccj ;
wire  cck ;
wire  ccl ;
wire  ccm ;
wire  ccn ;
wire  cco ;
wire  ccp ;
wire  CDA ;
wire  cdb ;
wire  cdc ;
wire  cdd ;
wire  cde ;
wire  cdf ;
wire  cdg ;
wire  cdh ;
wire  cdi ;
wire  cdj ;
wire  cdk ;
wire  cdl ;
wire  cdm ;
wire  cdn ;
wire  cdo ;
wire  cdp ;
wire  cea ;
wire  ceb ;
wire  cec ;
wire  ced ;
wire  cee ;
wire  cef ;
wire  ceg ;
wire  ceh ;
wire  cei ;
wire  cej ;
wire  cek ;
wire  cel ;
wire  cem ;
wire  cen ;
wire  ceo ;
wire  cep ;
wire  cfa ;
wire  cfb ;
wire  cfc ;
wire  cfd ;
wire  cfe ;
wire  cff ;
wire  cfg ;
wire  cfh ;
wire  cfi ;
wire  cfj ;
wire  cfk ;
wire  cfl ;
wire  cfm ;
wire  daf ;
wire  dag ;
wire  dah ;
wire  dai ;
wire  daj ;
wire  dak ;
wire  dal ;
wire  dam ;
wire  dan ;
wire  dao ;
wire  dap ;
wire  dba ;
wire  DBB ;
wire  DBC ;
wire  DBD ;
wire  DBE ;
wire  DBF ;
wire  DBG ;
wire  DBH ;
wire  DBI ;
wire  dbn ;
wire  dbo ;
wire  dbp ;
wire  dca ;
wire  dcb ;
wire  dcc ;
wire  dcd ;
wire  dce ;
wire  dcf ;
wire  dcg ;
wire  dch ;
wire  dci ;
wire  dcj ;
wire  dck ;
wire  dcl ;
wire  dcm ;
wire  dda ;
wire  ddb ;
wire  ddc ;
wire  ddd ;
wire  dde ;
wire  DDF ;
wire  DDG ;
wire  DDH ;
wire  DDI ;
wire  DDJ ;
wire  DDK ;
wire  DDL ;
wire  DDM ;
wire  deb ;
wire  dec ;
wire  ded ;
wire  dee ;
wire  def ;
wire  deg ;
wire  deh ;
wire  dei ;
wire  dej ;
wire  dek ;
wire  del ;
wire  dem ;
wire  DEN ;
wire  DEO ;
wire  DEP ;
wire  DFA ;
wire  DFB ;
wire  DFC ;
wire  DFD ;
wire  DFE ;
wire  dga ;
wire  dgb ;
wire  dgc ;
wire  dgd ;
wire  dge ;
wire  DGF ;
wire  DGG ;
wire  DGH ;
wire  DGI ;
wire  dgk ;
wire  dgl ;
wire  dgm ;
wire  dgn ;
wire  dgo ;
wire  dgp ;
wire  dha ;
wire  DHB ;
wire  DHC ;
wire  DHD ;
wire  DHE ;
wire  dhg ;
wire  dhh ;
wire  dhi ;
wire  dhj ;
wire  dhk ;
wire  dhl ;
wire  dhm ;
wire  DHN ;
wire  DHO ;
wire  DHP ;
wire  DIA ;
wire  dic ;
wire  did ;
wire  die ;
wire  dif ;
wire  dig ;
wire  dih ;
wire  dii ;
wire  dij ;
wire  dik ;
wire  dil ;
wire  dim ;
wire  din ;
wire  dio ;
wire  dip ;
wire  eaa ;
wire  EAA ;
wire  eab ;
wire  EAB ;
wire  eac ;
wire  EAC ;
wire  ead ;
wire  EAD ;
wire  eae ;
wire  EAE ;
wire  eaf ;
wire  EAF ;
wire  eag ;
wire  EAG ;
wire  eah ;
wire  EAH ;
wire  eai ;
wire  EAI ;
wire  eaj ;
wire  EAJ ;
wire  eak ;
wire  EAK ;
wire  eal ;
wire  EAL ;
wire  eam ;
wire  EAM ;
wire  ean ;
wire  EAN ;
wire  eao ;
wire  EAO ;
wire  eap ;
wire  EAP ;
wire  eaq ;
wire  EAQ ;
wire  ear ;
wire  EAR ;
wire  eas ;
wire  EAS ;
wire  eat ;
wire  EAT ;
wire  eau ;
wire  EAU ;
wire  eav ;
wire  EAV ;
wire  eaw ;
wire  EAW ;
wire  eax ;
wire  EAX ;
wire  eba ;
wire  EBA ;
wire  ebb ;
wire  EBB ;
wire  ebc ;
wire  EBC ;
wire  ebd ;
wire  EBD ;
wire  ebe ;
wire  EBE ;
wire  ebf ;
wire  EBF ;
wire  ebg ;
wire  EBG ;
wire  ebh ;
wire  EBH ;
wire  ebi ;
wire  EBI ;
wire  ebj ;
wire  EBJ ;
wire  ebk ;
wire  EBK ;
wire  ebl ;
wire  EBL ;
wire  ebm ;
wire  EBM ;
wire  ebn ;
wire  EBN ;
wire  ebo ;
wire  EBO ;
wire  ebp ;
wire  EBP ;
wire  ebq ;
wire  EBQ ;
wire  eca ;
wire  ECA ;
wire  ecb ;
wire  ECB ;
wire  ecc ;
wire  ECC ;
wire  ecd ;
wire  ECD ;
wire  ece ;
wire  ECE ;
wire  ecf ;
wire  ECF ;
wire  ecg ;
wire  ECG ;
wire  ech ;
wire  ECH ;
wire  eci ;
wire  ECI ;
wire  ecj ;
wire  ECJ ;
wire  eck ;
wire  ECK ;
wire  ecl ;
wire  ECL ;
wire  ecm ;
wire  ECM ;
wire  ecn ;
wire  ECN ;
wire  eco ;
wire  ECO ;
wire  ecp ;
wire  ECP ;
wire  ecq ;
wire  ECQ ;
wire  ecr ;
wire  ECR ;
wire  ecs ;
wire  ECS ;
wire  ect ;
wire  ECT ;
wire  ecu ;
wire  ECU ;
wire  ecv ;
wire  ECV ;
wire  ecw ;
wire  ECW ;
wire  ecx ;
wire  ECX ;
wire  eda ;
wire  EDA ;
wire  edb ;
wire  EDB ;
wire  edc ;
wire  EDC ;
wire  edd ;
wire  EDD ;
wire  ede ;
wire  EDE ;
wire  edf ;
wire  EDF ;
wire  edg ;
wire  EDG ;
wire  edh ;
wire  EDH ;
wire  edi ;
wire  EDI ;
wire  edj ;
wire  EDJ ;
wire  edk ;
wire  EDK ;
wire  edl ;
wire  EDL ;
wire  edm ;
wire  EDM ;
wire  edn ;
wire  EDN ;
wire  edo ;
wire  EDO ;
wire  edp ;
wire  EDP ;
wire  edq ;
wire  EDQ ;
wire  edr ;
wire  EDR ;
wire  eea ;
wire  EEA ;
wire  eeb ;
wire  EEB ;
wire  eec ;
wire  EEC ;
wire  eed ;
wire  EED ;
wire  eee ;
wire  EEE ;
wire  eef ;
wire  EEF ;
wire  eeg ;
wire  EEG ;
wire  eeh ;
wire  EEH ;
wire  eei ;
wire  EEI ;
wire  eej ;
wire  EEJ ;
wire  eek ;
wire  EEK ;
wire  eel ;
wire  EEL ;
wire  eem ;
wire  EEM ;
wire  een ;
wire  EEN ;
wire  eeo ;
wire  EEO ;
wire  eep ;
wire  EEP ;
wire  eeq ;
wire  EEQ ;
wire  eer ;
wire  EER ;
wire  ees ;
wire  EES ;
wire  eet ;
wire  EET ;
wire  eeu ;
wire  EEU ;
wire  eev ;
wire  EEV ;
wire  eew ;
wire  EEW ;
wire  eex ;
wire  EEX ;
wire  efa ;
wire  EFA ;
wire  efb ;
wire  EFB ;
wire  efc ;
wire  EFC ;
wire  efd ;
wire  EFD ;
wire  efe ;
wire  EFE ;
wire  eff ;
wire  EFF ;
wire  efg ;
wire  EFG ;
wire  efh ;
wire  EFH ;
wire  efi ;
wire  EFI ;
wire  efj ;
wire  EFJ ;
wire  efk ;
wire  EFK ;
wire  efl ;
wire  EFL ;
wire  efm ;
wire  EFM ;
wire  efn ;
wire  EFN ;
wire  efo ;
wire  EFO ;
wire  efp ;
wire  EFP ;
wire  efq ;
wire  EFQ ;
wire  efr ;
wire  EFR ;
wire  efs ;
wire  EFS ;
wire  ega ;
wire  EGA ;
wire  egb ;
wire  EGB ;
wire  egc ;
wire  EGC ;
wire  egd ;
wire  EGD ;
wire  ege ;
wire  EGE ;
wire  egf ;
wire  EGF ;
wire  egg ;
wire  EGG ;
wire  egh ;
wire  EGH ;
wire  egi ;
wire  EGI ;
wire  egj ;
wire  EGJ ;
wire  egk ;
wire  EGK ;
wire  egl ;
wire  EGL ;
wire  egm ;
wire  EGM ;
wire  egn ;
wire  EGN ;
wire  ego ;
wire  EGO ;
wire  egp ;
wire  EGP ;
wire  egq ;
wire  EGQ ;
wire  egr ;
wire  EGR ;
wire  egs ;
wire  EGS ;
wire  egt ;
wire  EGT ;
wire  egu ;
wire  EGU ;
wire  egv ;
wire  EGV ;
wire  egw ;
wire  EGW ;
wire  egx ;
wire  EGX ;
wire  eha ;
wire  EHA ;
wire  ehb ;
wire  EHB ;
wire  ehc ;
wire  EHC ;
wire  ehd ;
wire  EHD ;
wire  ehe ;
wire  EHE ;
wire  ehf ;
wire  EHF ;
wire  ehg ;
wire  EHG ;
wire  ehh ;
wire  EHH ;
wire  ehi ;
wire  EHI ;
wire  ehj ;
wire  EHJ ;
wire  ehk ;
wire  EHK ;
wire  ehl ;
wire  EHL ;
wire  ehm ;
wire  EHM ;
wire  ehn ;
wire  EHN ;
wire  eho ;
wire  EHO ;
wire  ehp ;
wire  EHP ;
wire  ehq ;
wire  EHQ ;
wire  ehr ;
wire  EHR ;
wire  ehs ;
wire  EHS ;
wire  eht ;
wire  EHT ;
wire  eia ;
wire  EIA ;
wire  eib ;
wire  EIB ;
wire  eic ;
wire  EIC ;
wire  eid ;
wire  EID ;
wire  eie ;
wire  EIE ;
wire  eif ;
wire  EIF ;
wire  eig ;
wire  EIG ;
wire  eih ;
wire  EIH ;
wire  eii ;
wire  EII ;
wire  eij ;
wire  EIJ ;
wire  eik ;
wire  EIK ;
wire  eil ;
wire  EIL ;
wire  eim ;
wire  EIM ;
wire  ein ;
wire  EIN ;
wire  eio ;
wire  EIO ;
wire  eip ;
wire  EIP ;
wire  eiq ;
wire  EIQ ;
wire  eir ;
wire  EIR ;
wire  eis ;
wire  EIS ;
wire  eit ;
wire  EIT ;
wire  eiu ;
wire  EIU ;
wire  eiv ;
wire  EIV ;
wire  eiw ;
wire  EIW ;
wire  eix ;
wire  EIX ;
wire  eja ;
wire  EJA ;
wire  ejb ;
wire  EJB ;
wire  ejc ;
wire  EJC ;
wire  ejd ;
wire  EJD ;
wire  eje ;
wire  EJE ;
wire  ejf ;
wire  EJF ;
wire  ejg ;
wire  EJG ;
wire  ejh ;
wire  EJH ;
wire  eji ;
wire  EJI ;
wire  ejj ;
wire  EJJ ;
wire  ejk ;
wire  EJK ;
wire  ejl ;
wire  EJL ;
wire  ejm ;
wire  EJM ;
wire  ejn ;
wire  EJN ;
wire  ejo ;
wire  EJO ;
wire  ejp ;
wire  EJP ;
wire  ejq ;
wire  EJQ ;
wire  ejr ;
wire  EJR ;
wire  ejs ;
wire  EJS ;
wire  ejt ;
wire  EJT ;
wire  eju ;
wire  EJU ;
wire  eka ;
wire  EKA ;
wire  ekb ;
wire  EKB ;
wire  ekc ;
wire  EKC ;
wire  ekd ;
wire  EKD ;
wire  eke ;
wire  EKE ;
wire  ekf ;
wire  EKF ;
wire  ekg ;
wire  EKG ;
wire  ekh ;
wire  EKH ;
wire  eki ;
wire  EKI ;
wire  ekj ;
wire  EKJ ;
wire  ekk ;
wire  EKK ;
wire  ekl ;
wire  EKL ;
wire  ekm ;
wire  EKM ;
wire  ekn ;
wire  EKN ;
wire  eko ;
wire  EKO ;
wire  ekp ;
wire  EKP ;
wire  ekq ;
wire  EKQ ;
wire  ekr ;
wire  EKR ;
wire  eks ;
wire  EKS ;
wire  ekt ;
wire  EKT ;
wire  eku ;
wire  EKU ;
wire  ekv ;
wire  EKV ;
wire  ekw ;
wire  EKW ;
wire  ekx ;
wire  EKX ;
wire  ela ;
wire  ELA ;
wire  elb ;
wire  ELB ;
wire  elc ;
wire  ELC ;
wire  eld ;
wire  ELD ;
wire  ele ;
wire  ELE ;
wire  elf ;
wire  ELF ;
wire  elg ;
wire  ELG ;
wire  elh ;
wire  ELH ;
wire  eli ;
wire  ELI ;
wire  elj ;
wire  ELJ ;
wire  elk ;
wire  ELK ;
wire  ell ;
wire  ELL ;
wire  elm ;
wire  ELM ;
wire  eln ;
wire  ELN ;
wire  elo ;
wire  ELO ;
wire  elp ;
wire  ELP ;
wire  elq ;
wire  ELQ ;
wire  elr ;
wire  ELR ;
wire  els ;
wire  ELS ;
wire  elt ;
wire  ELT ;
wire  elu ;
wire  ELU ;
wire  elv ;
wire  ELV ;
wire  ema ;
wire  EMA ;
wire  emb ;
wire  EMB ;
wire  emc ;
wire  EMC ;
wire  emd ;
wire  EMD ;
wire  eme ;
wire  EME ;
wire  emf ;
wire  EMF ;
wire  emg ;
wire  EMG ;
wire  emh ;
wire  EMH ;
wire  emi ;
wire  EMI ;
wire  emj ;
wire  EMJ ;
wire  emk ;
wire  EMK ;
wire  eml ;
wire  EML ;
wire  emm ;
wire  EMM ;
wire  emn ;
wire  EMN ;
wire  emo ;
wire  EMO ;
wire  emp ;
wire  EMP ;
wire  emq ;
wire  EMQ ;
wire  emr ;
wire  EMR ;
wire  ems ;
wire  EMS ;
wire  emt ;
wire  EMT ;
wire  emu ;
wire  EMU ;
wire  emv ;
wire  EMV ;
wire  emw ;
wire  EMW ;
wire  emx ;
wire  EMX ;
wire  ena ;
wire  ENA ;
wire  enb ;
wire  ENB ;
wire  enc ;
wire  ENC ;
wire  endd ;
wire  ENDD  ;
wire  ene ;
wire  ENE ;
wire  enf ;
wire  ENF ;
wire  eng ;
wire  ENG ;
wire  enh ;
wire  ENH ;
wire  eni ;
wire  ENI ;
wire  enj ;
wire  ENJ ;
wire  enk ;
wire  ENK ;
wire  enl ;
wire  ENL ;
wire  enm ;
wire  ENM ;
wire  enn ;
wire  ENN ;
wire  eno ;
wire  ENO ;
wire  enp ;
wire  ENP ;
wire  enq ;
wire  ENQ ;
wire  enr ;
wire  ENR ;
wire  ens ;
wire  ENS ;
wire  ent ;
wire  ENT ;
wire  enu ;
wire  ENU ;
wire  env ;
wire  ENV ;
wire  enw ;
wire  ENW ;
wire  eoa ;
wire  EOA ;
wire  eob ;
wire  EOB ;
wire  eoc ;
wire  EOC ;
wire  eod ;
wire  EOD ;
wire  eoe ;
wire  EOE ;
wire  eof ;
wire  EOF ;
wire  eog ;
wire  EOG ;
wire  eoh ;
wire  EOH ;
wire  eoi ;
wire  EOI ;
wire  eoj ;
wire  EOJ ;
wire  eok ;
wire  EOK ;
wire  eol ;
wire  EOL ;
wire  eom ;
wire  EOM ;
wire  eon ;
wire  EON ;
wire  eoo ;
wire  EOO ;
wire  eop ;
wire  EOP ;
wire  eoq ;
wire  EOQ ;
wire  eor ;
wire  EOR ;
wire  eos ;
wire  EOS ;
wire  eot ;
wire  EOT ;
wire  eou ;
wire  EOU ;
wire  eov ;
wire  EOV ;
wire  eow ;
wire  EOW ;
wire  eox ;
wire  EOX ;
wire  epa ;
wire  EPA ;
wire  epb ;
wire  EPB ;
wire  epc ;
wire  EPC ;
wire  epd ;
wire  EPD ;
wire  epe ;
wire  EPE ;
wire  epf ;
wire  EPF ;
wire  epg ;
wire  EPG ;
wire  eph ;
wire  EPH ;
wire  epi ;
wire  EPI ;
wire  epj ;
wire  EPJ ;
wire  epk ;
wire  EPK ;
wire  epl ;
wire  EPL ;
wire  epm ;
wire  EPM ;
wire  epn ;
wire  EPN ;
wire  epo ;
wire  EPO ;
wire  epp ;
wire  EPP ;
wire  epq ;
wire  EPQ ;
wire  epr ;
wire  EPR ;
wire  eps ;
wire  EPS ;
wire  ept ;
wire  EPT ;
wire  epu ;
wire  EPU ;
wire  epv ;
wire  EPV ;
wire  epw ;
wire  EPW ;
wire  epx ;
wire  EPX ;
wire  eqb ;
wire  EQB ;
wire  eqc ;
wire  EQC ;
wire  eqd ;
wire  EQD ;
wire  eqe ;
wire  EQE ;
wire  eqf ;
wire  EQF ;
wire  eqg ;
wire  EQG ;
wire  eqh ;
wire  EQH ;
wire  eqi ;
wire  EQI ;
wire  eqj ;
wire  EQJ ;
wire  eqk ;
wire  EQK ;
wire  eql ;
wire  EQL ;
wire  eqm ;
wire  EQM ;
wire  eqn ;
wire  EQN ;
wire  eqo ;
wire  EQO ;
wire  eqp ;
wire  EQP ;
wire  eqq ;
wire  EQQ ;
wire  eqr ;
wire  EQR ;
wire  eqs ;
wire  EQS ;
wire  eqt ;
wire  EQT ;
wire  equ ;
wire  EQU ;
wire  eqv ;
wire  EQV ;
wire  eqw ;
wire  EQW ;
wire  eqx ;
wire  EQX ;
wire  era ;
wire  ERA ;
wire  erb ;
wire  ERB ;
wire  erc ;
wire  ERC ;
wire  erd ;
wire  ERD ;
wire  ere ;
wire  ERE ;
wire  erf ;
wire  ERF ;
wire  erg ;
wire  ERG ;
wire  erh ;
wire  ERH ;
wire  eri ;
wire  ERI ;
wire  erj ;
wire  ERJ ;
wire  erk ;
wire  ERK ;
wire  erl ;
wire  ERL ;
wire  erm ;
wire  ERM ;
wire  ern ;
wire  ERN ;
wire  ero ;
wire  ERO ;
wire  erp ;
wire  ERP ;
wire  erq ;
wire  ERQ ;
wire  err ;
wire  ERR ;
wire  ers ;
wire  ERS ;
wire  ert ;
wire  ERT ;
wire  eru ;
wire  ERU ;
wire  erv ;
wire  ERV ;
wire  erw ;
wire  ERW ;
wire  erx ;
wire  ERX ;
wire  faa ;
wire  fab ;
wire  fac ;
wire  fad ;
wire  fae ;
wire  faf ;
wire  fag ;
wire  fah ;
wire  fai ;
wire  faj ;
wire  fak ;
wire  fal ;
wire  fam ;
wire  fan ;
wire  FBA ;
wire  FBB ;
wire  FBC ;
wire  FBD ;
wire  FBE ;
wire  FBF ;
wire  FBG ;
wire  FBH ;
wire  FBI ;
wire  FBJ ;
wire  FBK ;
wire  FBL ;
wire  FBM ;
wire  FBN ;
wire  fca ;
wire  fcb ;
wire  fcc ;
wire  fcd ;
wire  fce ;
wire  fcf ;
wire  fcg ;
wire  fch ;
wire  fci ;
wire  fcj ;
wire  fck ;
wire  fcl ;
wire  fcm ;
wire  fcn ;
wire  fco ;
wire  FDB ;
wire  FDC ;
wire  FDD ;
wire  FDE ;
wire  FDF ;
wire  FDG ;
wire  FDH ;
wire  FDI ;
wire  FDJ ;
wire  FDK ;
wire  FDL ;
wire  FDM ;
wire  FDN ;
wire  FDO ;
wire  fea ;
wire  feb ;
wire  fec ;
wire  fed ;
wire  fee ;
wire  fef ;
wire  feg ;
wire  feh ;
wire  fei ;
wire  fej ;
wire  fek ;
wire  fel ;
wire  fem ;
wire  fen ;
wire  feo ;
wire  fep ;
wire  FFC ;
wire  FFD ;
wire  FFE ;
wire  FFF ;
wire  FFG ;
wire  FFH ;
wire  FFI ;
wire  FFJ ;
wire  FFK ;
wire  FFL ;
wire  FFM ;
wire  FFN ;
wire  FFO ;
wire  FFP ;
wire  fga ;
wire  fgb ;
wire  fgc ;
wire  fgd ;
wire  fge ;
wire  fgf ;
wire  fgg ;
wire  fgh ;
wire  fgi ;
wire  fgj ;
wire  fgk ;
wire  fgl ;
wire  fgm ;
wire  fgn ;
wire  fgo ;
wire  FHA ;
wire  FHB ;
wire  FHC ;
wire  FHD ;
wire  FHE ;
wire  FHF ;
wire  FHG ;
wire  FHH ;
wire  FHI ;
wire  FHJ ;
wire  FHK ;
wire  FHL ;
wire  FHM ;
wire  FHN ;
wire  FHO ;
wire  fia ;
wire  fib ;
wire  fic ;
wire  fid ;
wire  fie ;
wire  fif ;
wire  fig ;
wire  fih ;
wire  fii ;
wire  fij ;
wire  fik ;
wire  fil ;
wire  fim ;
wire  fin ;
wire  fio ;
wire  fip ;
wire  FJB ;
wire  FJC ;
wire  FJD ;
wire  FJE ;
wire  FJF ;
wire  FJG ;
wire  FJH ;
wire  FJI ;
wire  FJJ ;
wire  FJK ;
wire  FJL ;
wire  FJM ;
wire  FJN ;
wire  FJO ;
wire  FJP ;
wire  fka ;
wire  fkb ;
wire  fkc ;
wire  fkd ;
wire  fke ;
wire  fkf ;
wire  fkg ;
wire  fkh ;
wire  fki ;
wire  fkj ;
wire  fkk ;
wire  fkl ;
wire  fkm ;
wire  fkn ;
wire  fko ;
wire  fkp ;
wire  fkq ;
wire  FLC ;
wire  FLD ;
wire  FLE ;
wire  FLF ;
wire  FLG ;
wire  FLH ;
wire  FLI ;
wire  FLJ ;
wire  FLK ;
wire  FLL ;
wire  FLM ;
wire  FLN ;
wire  FLO ;
wire  FLP ;
wire  FLQ ;
wire  fma ;
wire  fmb ;
wire  fmc ;
wire  fmd ;
wire  fme ;
wire  fmf ;
wire  fmg ;
wire  fmh ;
wire  fmi ;
wire  fmj ;
wire  fmk ;
wire  fml ;
wire  fmm ;
wire  fmn ;
wire  fmo ;
wire  fmp ;
wire  FNA ;
wire  FNB ;
wire  FNC ;
wire  FND ;
wire  FNE ;
wire  FNF ;
wire  FNG ;
wire  FNH ;
wire  FNI ;
wire  FNJ ;
wire  FNK ;
wire  FNL ;
wire  FNM ;
wire  FNN ;
wire  FNO ;
wire  FNP ;
wire  foa ;
wire  fob ;
wire  foc ;
wire  fod ;
wire  foe ;
wire  fof ;
wire  fog ;
wire  foh ;
wire  foi ;
wire  foj ;
wire  fok ;
wire  fol ;
wire  fom ;
wire  fon ;
wire  foo ;
wire  fop ;
wire  foq ;
wire  FPB ;
wire  FPC ;
wire  FPD ;
wire  FPE ;
wire  FPF ;
wire  FPG ;
wire  FPH ;
wire  FPI ;
wire  FPJ ;
wire  FPK ;
wire  FPL ;
wire  FPM ;
wire  FPN ;
wire  FPO ;
wire  FPP ;
wire  FPQ ;
wire  fqa ;
wire  fqb ;
wire  fqc ;
wire  fqd ;
wire  fqe ;
wire  fqf ;
wire  fqg ;
wire  fqh ;
wire  fqi ;
wire  fqj ;
wire  fqk ;
wire  fql ;
wire  fqm ;
wire  fqn ;
wire  fqo ;
wire  fqp ;
wire  gaa ;
wire  GAA ;
wire  gab ;
wire  GAB ;
wire  gac ;
wire  GAC ;
wire  gad ;
wire  GAD ;
wire  gba ;
wire  GBA ;
wire  gbb ;
wire  GBB ;
wire  gbc ;
wire  GBC ;
wire  gbd ;
wire  GBD ;
wire  gca ;
wire  GCA ;
wire  gcb ;
wire  GCB ;
wire  gcc ;
wire  GCC ;
wire  gcd ;
wire  GCD ;
wire  gce ;
wire  GCE ;
wire  gcf ;
wire  GCF ;
wire  gcg ;
wire  GCG ;
wire  gch ;
wire  GCH ;
wire  gci ;
wire  GCI ;
wire  gda ;
wire  GDA ;
wire  gdb ;
wire  GDB ;
wire  gdc ;
wire  GDC ;
wire  gdd ;
wire  GDD ;
wire  gde ;
wire  GDE ;
wire  gdf ;
wire  GDF ;
wire  gdg ;
wire  GDG ;
wire  gdh ;
wire  GDH ;
wire  gdi ;
wire  GDI ;
wire  gea ;
wire  GEA ;
wire  geb ;
wire  GEB ;
wire  gec ;
wire  GEC ;
wire  ged ;
wire  GED ;
wire  gee ;
wire  GEE ;
wire  gef ;
wire  GEF ;
wire  geg ;
wire  GEG ;
wire  geh ;
wire  GEH ;
wire  gei ;
wire  GEI ;
wire  gej ;
wire  GEJ ;
wire  gfa ;
wire  GFA ;
wire  gfb ;
wire  GFB ;
wire  gfc ;
wire  GFC ;
wire  gfd ;
wire  GFD ;
wire  gfe ;
wire  GFE ;
wire  gff ;
wire  GFF ;
wire  gfg ;
wire  GFG ;
wire  gfh ;
wire  GFH ;
wire  gfi ;
wire  GFI ;
wire  gfj ;
wire  GFJ ;
wire  gga ;
wire  GGA ;
wire  ggb ;
wire  GGB ;
wire  ggc ;
wire  GGC ;
wire  ggd ;
wire  GGD ;
wire  gge ;
wire  GGE ;
wire  ggf ;
wire  GGF ;
wire  ggg ;
wire  GGG ;
wire  ggh ;
wire  GGH ;
wire  ggi ;
wire  GGI ;
wire  gha ;
wire  GHA ;
wire  ghb ;
wire  GHB ;
wire  ghc ;
wire  GHC ;
wire  ghd ;
wire  GHD ;
wire  ghe ;
wire  GHE ;
wire  ghf ;
wire  GHF ;
wire  ghg ;
wire  GHG ;
wire  ghh ;
wire  GHH ;
wire  ghi ;
wire  GHI ;
wire  gia ;
wire  GIA ;
wire  gib ;
wire  GIB ;
wire  gic ;
wire  GIC ;
wire  gid ;
wire  GID ;
wire  gie ;
wire  GIE ;
wire  gif ;
wire  GIF ;
wire  gig ;
wire  GIG ;
wire  gih ;
wire  GIH ;
wire  gii ;
wire  GII ;
wire  gij ;
wire  GIJ ;
wire  gja ;
wire  GJA ;
wire  gjb ;
wire  GJB ;
wire  gjc ;
wire  GJC ;
wire  gjd ;
wire  GJD ;
wire  gje ;
wire  GJE ;
wire  gjf ;
wire  GJF ;
wire  gjg ;
wire  GJG ;
wire  gjh ;
wire  GJH ;
wire  gji ;
wire  GJI ;
wire  gjj ;
wire  GJJ ;
wire  gka ;
wire  GKA ;
wire  gkb ;
wire  GKB ;
wire  gkc ;
wire  GKC ;
wire  gkd ;
wire  GKD ;
wire  gke ;
wire  GKE ;
wire  gkf ;
wire  GKF ;
wire  gkg ;
wire  GKG ;
wire  gkh ;
wire  GKH ;
wire  gki ;
wire  GKI ;
wire  gkj ;
wire  GKJ ;
wire  gla ;
wire  GLA ;
wire  glb ;
wire  GLB ;
wire  glc ;
wire  GLC ;
wire  gld ;
wire  GLD ;
wire  gle ;
wire  GLE ;
wire  glf ;
wire  GLF ;
wire  glg ;
wire  GLG ;
wire  glh ;
wire  GLH ;
wire  gli ;
wire  GLI ;
wire  glj ;
wire  GLJ ;
wire  gma ;
wire  GMA ;
wire  gmb ;
wire  GMB ;
wire  gmc ;
wire  GMC ;
wire  gmd ;
wire  GMD ;
wire  gme ;
wire  GME ;
wire  gmf ;
wire  GMF ;
wire  gmg ;
wire  GMG ;
wire  gmh ;
wire  GMH ;
wire  gmi ;
wire  GMI ;
wire  gmj ;
wire  GMJ ;
wire  gna ;
wire  GNA ;
wire  gnb ;
wire  GNB ;
wire  gnc ;
wire  GNC ;
wire  gnd ;
wire  GND ;
wire  gne ;
wire  GNE ;
wire  gnf ;
wire  GNF ;
wire  gng ;
wire  GNG ;
wire  gnh ;
wire  GNH ;
wire  gni ;
wire  GNI ;
wire  gnj ;
wire  GNJ ;
wire  goa ;
wire  GOA ;
wire  gob ;
wire  GOB ;
wire  goc ;
wire  GOC ;
wire  god ;
wire  GOD ;
wire  goe ;
wire  GOE ;
wire  gof ;
wire  GOF ;
wire  gog ;
wire  GOG ;
wire  goh ;
wire  GOH ;
wire  goi ;
wire  GOI ;
wire  goj ;
wire  GOJ ;
wire  gok ;
wire  GOK ;
wire  gpa ;
wire  GPA ;
wire  gpb ;
wire  GPB ;
wire  gpc ;
wire  GPC ;
wire  gpd ;
wire  GPD ;
wire  gpe ;
wire  GPE ;
wire  gpf ;
wire  GPF ;
wire  gpg ;
wire  GPG ;
wire  gph ;
wire  GPH ;
wire  gpi ;
wire  GPI ;
wire  gpj ;
wire  GPJ ;
wire  gpk ;
wire  GPK ;
wire  gqa ;
wire  GQA ;
wire  gqb ;
wire  GQB ;
wire  gqc ;
wire  GQC ;
wire  gqd ;
wire  GQD ;
wire  gqe ;
wire  GQE ;
wire  gqf ;
wire  GQF ;
wire  gqg ;
wire  GQG ;
wire  gqh ;
wire  GQH ;
wire  gqi ;
wire  GQI ;
wire  gqj ;
wire  GQJ ;
wire  gra ;
wire  GRA ;
wire  grb ;
wire  GRB ;
wire  grc ;
wire  GRC ;
wire  grd ;
wire  GRD ;
wire  gre ;
wire  GRE ;
wire  grf ;
wire  GRF ;
wire  grg ;
wire  GRG ;
wire  grh ;
wire  GRH ;
wire  gri ;
wire  GRI ;
wire  grj ;
wire  GRJ ;
wire  haa ;
wire  hab ;
wire  HBA ;
wire  HBB ;
wire  hca ;
wire  hcb ;
wire  hcc ;
wire  hcd ;
wire  hce ;
wire  HDA ;
wire  HDB ;
wire  HDC ;
wire  HDD ;
wire  HDE ;
wire  hea ;
wire  heb ;
wire  hec ;
wire  hed ;
wire  hee ;
wire  hef ;
wire  heg ;
wire  HFA ;
wire  HFB ;
wire  HFC ;
wire  HFD ;
wire  HFE ;
wire  HFF ;
wire  hga ;
wire  hgb ;
wire  hgc ;
wire  hgd ;
wire  hge ;
wire  hgf ;
wire  hgg ;
wire  HHA ;
wire  HHB ;
wire  HHC ;
wire  HHD ;
wire  HHE ;
wire  HHF ;
wire  HHG ;
wire  hia ;
wire  hib ;
wire  hic ;
wire  hid ;
wire  hie ;
wire  hif ;
wire  hig ;
wire  hih ;
wire  HJA ;
wire  HJB ;
wire  HJC ;
wire  HJD ;
wire  HJE ;
wire  HJF ;
wire  hka ;
wire  hkb ;
wire  hkc ;
wire  hkd ;
wire  hke ;
wire  hkf ;
wire  hkg ;
wire  hkh ;
wire  HLA ;
wire  HLB ;
wire  HLC ;
wire  HLD ;
wire  HLE ;
wire  HLF ;
wire  HLG ;
wire  hma ;
wire  hmb ;
wire  hmc ;
wire  hmd ;
wire  hme ;
wire  hmf ;
wire  hmg ;
wire  HNA ;
wire  HNB ;
wire  HNC ;
wire  HND ;
wire  HNE ;
wire  HNF ;
wire  HNG ;
wire  hoa ;
wire  hob ;
wire  hoc ;
wire  hod ;
wire  hoe ;
wire  hof ;
wire  hog ;
wire  HPA ;
wire  HPB ;
wire  HPC ;
wire  HPD ;
wire  HPE ;
wire  HPF ;
wire  HPG ;
wire  hqa ;
wire  hqb ;
wire  hqc ;
wire  hqd ;
wire  hqe ;
wire  hqf ;
wire  hqg ;
wire  hqh ;
wire  hqi ;
wire  iaa ;
wire  iab ;
wire  iac ;
wire  iad ;
wire  iae ;
wire  iaf ;
wire  iag ;
wire  iah ;
wire  iai ;
wire  iaj ;
wire  iak ;
wire  ial ;
wire  iam ;
wire  ian ;
wire  iao ;
wire  iap ;
wire  iba ;
wire  ibb ;
wire  ibc ;
wire  ibd ;
wire  ibe ;
wire  ibf ;
wire  ibg ;
wire  ibh ;
wire  ibi ;
wire  ibj ;
wire  ibk ;
wire  ibl ;
wire  ibm ;
wire  ibn ;
wire  ibo ;
wire  ibp ;
wire  ica ;
wire  icb ;
wire  icc ;
wire  icd ;
wire  ice ;
wire  icf ;
wire  icg ;
wire  ich ;
wire  ici ;
wire  icj ;
wire  ick ;
wire  icl ;
wire  icm ;
wire  icn ;
wire  ico ;
wire  icp ;
wire  ida ;
wire  idb ;
wire  idc ;
wire  idd ;
wire  ide ;
wire  idf ;
wire  idg ;
wire  idh ;
wire  idi ;
wire  idj ;
wire  idk ;
wire  idl ;
wire  idm ;
wire  idn ;
wire  ido ;
wire  idp ;
wire  iea ;
wire  ieb ;
wire  iec ;
wire  ied ;
wire  iee ;
wire  ief ;
wire  ieg ;
wire  ieh ;
wire  iei ;
wire  iej ;
wire  iek ;
wire  iel ;
wire  iem ;
wire  ien ;
wire  ieo ;
wire  iep ;
wire  ieq ;
wire  ier ;
wire  ies ;
wire  iet ;
wire  ieu ;
wire  iev ;
wire  iew ;
wire  iex ;
wire  iey ;
wire  iez ;
wire  ifa ;
wire  ifb ;
wire  ifc ;
wire  ifd ;
wire  ife ;
wire  ifff  ;
wire  ifg ;
wire  ifh ;
wire  ifi ;
wire  ifj ;
wire  ifk ;
wire  ifl ;
wire  ifm ;
wire  ifn ;
wire  ifo ;
wire  ifp ;
wire  iga ;
wire  iha ;
wire  ika ;
wire  imm ;
wire  imr ;
wire  ims ;
wire  ira ;
wire  isa ;
wire  ita ;
wire  jba ;
wire  JBA ;
wire  jca ;
wire  JCA ;
wire  jcb ;
wire  JCB ;
wire  jda ;
wire  JDA ;
wire  jdb ;
wire  JDB ;
wire  jea ;
wire  JEA ;
wire  jeb ;
wire  JEB ;
wire  jec ;
wire  JEC ;
wire  jed ;
wire  JED ;
wire  jfa ;
wire  JFA ;
wire  jfb ;
wire  JFB ;
wire  jfc ;
wire  JFC ;
wire  jfd ;
wire  JFD ;
wire  jga ;
wire  JGA ;
wire  jgb ;
wire  JGB ;
wire  jgc ;
wire  JGC ;
wire  jgd ;
wire  JGD ;
wire  jha ;
wire  JHA ;
wire  jhb ;
wire  JHB ;
wire  jhc ;
wire  JHC ;
wire  jhd ;
wire  JHD ;
wire  jia ;
wire  JIA ;
wire  jib ;
wire  JIB ;
wire  jic ;
wire  JIC ;
wire  jid ;
wire  JID ;
wire  jie ;
wire  JIE ;
wire  jja ;
wire  JJA ;
wire  jjb ;
wire  JJB ;
wire  jjc ;
wire  JJC ;
wire  jjd ;
wire  JJD ;
wire  jje ;
wire  JJE ;
wire  jka ;
wire  JKA ;
wire  jkb ;
wire  JKB ;
wire  jkc ;
wire  JKC ;
wire  jkd ;
wire  JKD ;
wire  jla ;
wire  JLA ;
wire  jlb ;
wire  JLB ;
wire  jlc ;
wire  JLC ;
wire  jld ;
wire  JLD ;
wire  jma ;
wire  JMA ;
wire  jmb ;
wire  JMB ;
wire  jmc ;
wire  JMC ;
wire  jmd ;
wire  JMD ;
wire  jna ;
wire  JNA ;
wire  jnb ;
wire  JNB ;
wire  jnc ;
wire  JNC ;
wire  jnd ;
wire  JND ;
wire  joa ;
wire  JOA ;
wire  job ;
wire  JOB ;
wire  joc ;
wire  JOC ;
wire  jod ;
wire  JOD ;
wire  jpa ;
wire  JPA ;
wire  jpb ;
wire  JPB ;
wire  jpc ;
wire  JPC ;
wire  jpd ;
wire  JPD ;
wire  jqa ;
wire  JQA ;
wire  jqb ;
wire  JQB ;
wire  jqc ;
wire  JQC ;
wire  jqd ;
wire  JQD ;
wire  jqe ;
wire  JQE ;
wire  jra ;
wire  JRA ;
wire  jrb ;
wire  JRB ;
wire  jrc ;
wire  JRC ;
wire  jrd ;
wire  JRD ;
wire  jre ;
wire  JRE ;
wire  kca ;
wire  kcb ;
wire  KDA ;
wire  kea ;
wire  keb ;
wire  KFA ;
wire  KFB ;
wire  kga ;
wire  kgb ;
wire  kgc ;
wire  KHA ;
wire  KHB ;
wire  KHC ;
wire  kia ;
wire  kib ;
wire  kic ;
wire  KJA ;
wire  KJB ;
wire  KJC ;
wire  kka ;
wire  kkb ;
wire  kkc ;
wire  kkd ;
wire  kke ;
wire  KLA ;
wire  KLB ;
wire  KLC ;
wire  kma ;
wire  kmb ;
wire  kmc ;
wire  kmd ;
wire  KNA ;
wire  KNB ;
wire  KNC ;
wire  koa ;
wire  kob ;
wire  koc ;
wire  kod ;
wire  KPA ;
wire  KPB ;
wire  KPC ;
wire  kqa ;
wire  kqb ;
wire  kqc ;
wire  kqd ;
wire  lda ;
wire  LDA ;
wire  lea ;
wire  LEA ;
wire  lfa ;
wire  LFA ;
wire  lga ;
wire  LGA ;
wire  lha ;
wire  LHA ;
wire  lia ;
wire  LIA ;
wire  lib ;
wire  LIB ;
wire  lja ;
wire  LJA ;
wire  ljb ;
wire  LJB ;
wire  lka ;
wire  LKA ;
wire  lkb ;
wire  LKB ;
wire  lla ;
wire  LLA ;
wire  llb ;
wire  LLB ;
wire  lma ;
wire  LMA ;
wire  lmb ;
wire  LMB ;
wire  lna ;
wire  LNA ;
wire  lnb ;
wire  LNB ;
wire  loa ;
wire  LOA ;
wire  lob ;
wire  LOB ;
wire  lpa ;
wire  LPA ;
wire  lpb ;
wire  LPB ;
wire  lqa ;
wire  LQA ;
wire  lqb ;
wire  LQB ;
wire  lra ;
wire  LRA ;
wire  lrb ;
wire  LRB ;
wire  MFA ;
wire  mga ;
wire  mgb ;
wire  MHA ;
wire  mia ;
wire  MJA ;
wire  mka ;
wire  mkb ;
wire  MLA ;
wire  MLB ;
wire  mma ;
wire  mmb ;
wire  mmc ;
wire  MNA ;
wire  moa ;
wire  mob ;
wire  moc ;
wire  MPA ;
wire  mqa ;
wire  mqb ;
wire  mqc ;
wire  nha ;
wire  NHA ;
wire  nma ;
wire  NMA ;
wire  nna ;
wire  NNA ;
wire  noa ;
wire  NOA ;
wire  npa ;
wire  NPA ;
wire  nqa ;
wire  NQA ;
wire  nra ;
wire  NRA ;
wire  oaa ;
wire  oab ;
wire  oac ;
wire  oad ;
wire  oae ;
wire  oaf ;
wire  oag ;
wire  oah ;
wire  oai ;
wire  oaj ;
wire  oak ;
wire  oal ;
wire  oam ;
wire  oan ;
wire  oao ;
wire  oap ;
wire  oba ;
wire  obb ;
wire  obc ;
wire  obd ;
wire  obe ;
wire  obf ;
wire  obg ;
wire  obh ;
wire  obi ;
wire  obj ;
wire  obk ;
wire  obl ;
wire  obm ;
wire  obn ;
wire  obo ;
wire  obp ;
wire  ocg ;
wire  och ;
wire  oci ;
wire  ocj ;
wire  ock ;
wire  ocl ;
wire  ocm ;
wire  ocn ;
wire  oco ;
wire  ocp ;
wire  oda ;
wire  odb ;
wire  odc ;
wire  odd ;
wire  ode ;
wire  odf ;
wire  odg ;
wire  odh ;
wire  odi ;
wire  odj ;
wire  odk ;
wire  odl ;
wire  odm ;
wire  odn ;
wire  odo ;
wire  odp ;
wire  oea ;
wire  oeb ;
wire  oec ;
wire  oed ;
wire  oee ;
wire  oef ;
wire  oeg ;
wire  oeh ;
wire  oei ;
wire  oej ;
wire  oek ;
wire  oel ;
wire  oem ;
wire  oen ;
wire  oeo ;
wire  oep ;
wire  ofg ;
wire  ofh ;
wire  ofi ;
wire  ofj ;
wire  ofk ;
wire  ofl ;
wire  ofm ;
wire  ofn ;
wire  ofo ;
wire  ofp ;
wire  OGA ;
wire  OGB ;
wire  OGC ;
wire  OGD ;
wire  OGE ;
wire  OGF ;
wire  OGG ;
wire  OGH ;
wire  OGI ;
wire  OGJ ;
wire  OGK ;
wire  OGL ;
wire  OGM ;
wire  OGN ;
wire  OGO ;
wire  OGP ;
wire  OHA ;
wire  OHB ;
wire  OHC ;
wire  OHD ;
wire  OHE ;
wire  OHF ;
wire  OHG ;
wire  ohh ;
wire  ohi ;
wire  ohj ;
wire  ohk ;
wire  OIH ;
wire  OII ;
wire  OIJ ;
wire  OKA ;
wire  OKB ;
wire  OKC ;
wire  okd ;
wire  oke ;
wire  okf ;
wire  OLD ;
wire  OMA ;
wire  omb ;
wire  ONB ;
wire  opk ;
wire  opm ;
wire  opo ;
wire  opq ;
wire  opr ;
wire  OQJ ;
wire  OQK ;
wire  OQM ;
wire  OQO ;
wire  OQQ ;
wire  qaa ;
wire  qab ;
wire  qac ;
wire  qad ;
wire  qae ;
wire  qaf ;
wire  qag ;
wire  qah ;
wire  qai ;
wire  qga ;
wire  qha ;
wire  qka ;
wire  qmm ;
wire  qmr ;
wire  qms ;
wire  qra ;
wire  qsa ;
wire  qta ;
wire  tam ;
wire  tar ;
wire  tas ;
wire  tga ;
wire  TGB ;
wire  tgc ;
wire  TGD ;
wire  tge ;
wire  TGF ;
wire  tha ;
wire  THB ;
wire  thc ;
wire  THD ;
wire  the ;
wire  THF ;
wire  tka ;
wire  TKB ;
wire  tkc ;
wire  TKD ;
wire  tke ;
wire  TKF ;
wire  tra ;
wire  trb ;
wire  TRC ;
wire  tsa ;
wire  TSB ;
wire  tsc ;
wire  TSD ;
wire  tse ;
wire  TSF ;
wire  tta ;
wire  TTB ;
wire  ttc ;
wire  TTD ;
wire  tte ;
wire  TTF ;
wire  ZZI ;
wire  ZZO ;
assign ZZI = 1'b1;
assign ZZO = 1'b0;
assign EBO =  DCG & CDC  ; 
assign ebo = ~EBO;  //complement 
assign EBP =  DCH & CDB  ; 
assign ebp = ~EBP;  //complement 
assign EBQ =  DCI & CDA  ; 
assign ebq = ~EBQ;  //complement 
assign EDP =  DCH & CDC  ; 
assign edp = ~EDP;  //complement 
assign EDQ =  DCI & CDB  ; 
assign edq = ~EDQ;  //complement 
assign EDR =  DCJ & CDA  ; 
assign edr = ~EDR;  //complement 
assign EFQ =  DCI & CDC  ; 
assign efq = ~EFQ;  //complement 
assign EFR =  DCJ & CDB  ; 
assign efr = ~EFR;  //complement 
assign EFS =  DCK & CDA  ; 
assign efs = ~EFS;  //complement 
assign EHR =  DCJ & CDC  ; 
assign ehr = ~EHR;  //complement 
assign EHS =  DCK & CDB  ; 
assign ehs = ~EHS;  //complement 
assign EHT =  DCL & CDA  ; 
assign eht = ~EHT;  //complement 
assign fan = ~FAN;  //complement 
assign FBN = ~fbn;  //complement 
assign fco = ~FCO;  //complement 
assign FDO = ~fdo;  //complement 
assign fep = ~FEP;  //complement 
assign FFP = ~ffp;  //complement 
assign fgo = ~FGO;  //complement 
assign FHO = ~fho;  //complement 
assign EBL =  DCD & CDF  ; 
assign ebl = ~EBL;  //complement 
assign EBM =  DCE & CDE  ; 
assign ebm = ~EBM;  //complement 
assign EBN =  DCF & CDD  ; 
assign ebn = ~EBN;  //complement 
assign fem = ~FEM;  //complement 
assign FFM = ~ffm;  //complement 
assign EFN =  DCF & CDF  ; 
assign efn = ~EFN;  //complement 
assign EFO =  DCG & CDE  ; 
assign efo = ~EFO;  //complement 
assign EFP =  DCH & CDD  ; 
assign efp = ~EFP;  //complement 
assign EHO =  DCG & CDF  ; 
assign eho = ~EHO;  //complement 
assign EHP =  DCH & CDE  ; 
assign ehp = ~EHP;  //complement 
assign EHQ =  DCI & CDD  ; 
assign ehq = ~EHQ;  //complement 
assign fam = ~FAM;  //complement 
assign FBM = ~fbm;  //complement 
assign fcn = ~FCN;  //complement 
assign FDN = ~fdn;  //complement 
assign feo = ~FEO;  //complement 
assign FFO = ~ffo;  //complement 
assign fgn = ~FGN;  //complement 
assign FHN = ~fhn;  //complement 
assign EBI =  DCA & CDI  ; 
assign ebi = ~EBI;  //complement 
assign EBJ =  DCB & CDH  ; 
assign ebj = ~EBJ;  //complement 
assign EBK =  DCC & CDG  ; 
assign ebk = ~EBK;  //complement 
assign EDJ =  DCB & CDI  ; 
assign edj = ~EDJ;  //complement 
assign EDK =  DCC & CDH  ; 
assign edk = ~EDK;  //complement 
assign EDL =  DCD & CDG  ; 
assign edl = ~EDL;  //complement 
assign EFK =  DCC & CDI  ; 
assign efk = ~EFK;  //complement 
assign EFL =  DCD & CDH  ; 
assign efl = ~EFL;  //complement 
assign EFM =  DCE & CDG  ; 
assign efm = ~EFM;  //complement 
assign EHL =  DCD & CDI  ; 
assign ehl = ~EHL;  //complement 
assign EHM =  DCE & CDH  ; 
assign ehm = ~EHM;  //complement 
assign EHN =  DCF & CDG  ; 
assign ehn = ~EHN;  //complement 
assign fal = ~FAL;  //complement 
assign FBL = ~fbl;  //complement 
assign fcm = ~FCM;  //complement 
assign FDM = ~fdm;  //complement 
assign fgm = ~FGM;  //complement 
assign FHM = ~fhm;  //complement 
assign EBF =  DBN & CDL  ; 
assign ebf = ~EBF;  //complement 
assign EBG =  DBO & CDK  ; 
assign ebg = ~EBG;  //complement 
assign EBH =  DBP & CDJ  ; 
assign ebh = ~EBH;  //complement 
assign EDG =  DBO & CDL  ; 
assign edg = ~EDG;  //complement 
assign EDH =  DBP & CDK  ; 
assign edh = ~EDH;  //complement 
assign EDI =  DCA & CDJ  ; 
assign edi = ~EDI;  //complement 
assign EDM =  DCE & CDF  ; 
assign edm = ~EDM;  //complement 
assign EDN =  DCF & CDE  ; 
assign edn = ~EDN;  //complement 
assign EDO =  DCG & CDD  ; 
assign edo = ~EDO;  //complement 
assign EHI =  DCA & CDL  ; 
assign ehi = ~EHI;  //complement 
assign EHJ =  DCB & CDK  ; 
assign ehj = ~EHJ;  //complement 
assign EHK =  DCC & CDJ  ; 
assign ehk = ~EHK;  //complement 
assign fak = ~FAK;  //complement 
assign FBK = ~fbk;  //complement 
assign fcl = ~FCL;  //complement 
assign FDL = ~fdl;  //complement 
assign EFH =  DBP & CDL  ; 
assign efh = ~EFH;  //complement 
assign EFI =  DCA & CDK  ; 
assign efi = ~EFI;  //complement 
assign EFJ =  DCB & CDJ  ; 
assign efj = ~EFJ;  //complement 
assign fgl = ~FGL;  //complement 
assign FHL = ~fhl;  //complement 
assign EJS =  DCK & CDC  ; 
assign ejs = ~EJS;  //complement 
assign EJT =  DCL & CDB  ; 
assign ejt = ~EJT;  //complement 
assign EJU =  DCM & CDA  ; 
assign eju = ~EJU;  //complement 
assign CDA = ~cda;  //complement 
assign cdb = ~CDB;  //complement 
assign cdc = ~CDC;  //complement 
assign ELT =  DIL & CAC  ; 
assign elt = ~ELT;  //complement 
assign ELU =  DIM & CAB  ; 
assign elu = ~ELU;  //complement 
assign ELV =  DIN & CAA  ; 
assign elv = ~ELV;  //complement 
assign fip = ~FIP;  //complement 
assign FJP = ~fjp;  //complement 
assign dcj = ~DCJ;  //complement 
assign dck = ~DCK;  //complement 
assign dcl = ~DCL;  //complement 
assign dcm = ~DCM;  //complement 
assign fkq = ~FKQ;  //complement 
assign FLQ = ~flq;  //complement 
assign EJP =  DCH & CDF  ; 
assign ejp = ~EJP;  //complement 
assign EJQ =  DCI & CDE  ; 
assign ejq = ~EJQ;  //complement 
assign EJR =  DCJ & CDD  ; 
assign ejr = ~EJR;  //complement 
assign cdd = ~CDD;  //complement 
assign cde = ~CDE;  //complement 
assign cdf = ~CDF;  //complement 
assign ELQ =  DII & CAF  ; 
assign elq = ~ELQ;  //complement 
assign ELR =  DIJ & CAE  ; 
assign elr = ~ELR;  //complement 
assign ELS =  DIK & CAD  ; 
assign els = ~ELS;  //complement 
assign fen = ~FEN;  //complement 
assign FFN = ~ffn;  //complement 
assign fio = ~FIO;  //complement 
assign FJO = ~fjo;  //complement 
assign dcf = ~DCF;  //complement 
assign dcg = ~DCG;  //complement 
assign dch = ~DCH;  //complement 
assign dci = ~DCI;  //complement 
assign fkp = ~FKP;  //complement 
assign FLP = ~flp;  //complement 
assign EJN =  DCF & CDH  ; 
assign ejn = ~EJN;  //complement 
assign EJM =  DCE & CDI  ; 
assign ejm = ~EJM;  //complement 
assign EJO =  DCG & CDG  ; 
assign ejo = ~EJO;  //complement 
assign cdg = ~CDG;  //complement 
assign cdh = ~CDH;  //complement 
assign cdi = ~CDI;  //complement 
assign ELN =  DIF & CAI  ; 
assign eln = ~ELN;  //complement 
assign ELO =  DIG & CAH  ; 
assign elo = ~ELO;  //complement 
assign ELP =  DIH & CAG  ; 
assign elp = ~ELP;  //complement 
assign fin = ~FIN;  //complement 
assign FJN = ~fjn;  //complement 
assign dcb = ~DCB;  //complement 
assign dcd = ~DCD;  //complement 
assign dcc = ~DCC;  //complement 
assign dce = ~DCE;  //complement 
assign fko = ~FKO;  //complement 
assign FLO = ~flo;  //complement 
assign EJJ =  DCB & CDL  ; 
assign ejj = ~EJJ;  //complement 
assign EJK =  DCC & CDK  ; 
assign ejk = ~EJK;  //complement 
assign EJL =  DCD & CDJ  ; 
assign ejl = ~EJL;  //complement 
assign cdj = ~CDJ;  //complement 
assign cdk = ~CDK;  //complement 
assign cdl = ~CDL;  //complement 
assign ELK =  DIC & CAL  ; 
assign elk = ~ELK;  //complement 
assign ELM =  DIE & CAJ  ; 
assign elm = ~ELM;  //complement 
assign ELL =  DID & CAK  ; 
assign ell = ~ELL;  //complement 
assign fim = ~FIM;  //complement 
assign FJM = ~fjm;  //complement 
assign dbn = ~DBN;  //complement 
assign dbo = ~DBO;  //complement 
assign dbp = ~DBP;  //complement 
assign dca = ~DCA;  //complement 
assign fkn = ~FKN;  //complement 
assign FLN = ~fln;  //complement 
assign ENU =  DIM & CAC  ; 
assign enu = ~ENU;  //complement 
assign ENV =  DIN & CAB  ; 
assign env = ~ENV;  //complement 
assign ENW =  DIO & CAA  ; 
assign enw = ~ENW;  //complement 
assign EPV =  DIN & CAC  ; 
assign epv = ~EPV;  //complement 
assign EPW =  DIO & CAB  ; 
assign epw = ~EPW;  //complement 
assign EPX =  DIP & CAA  ; 
assign epx = ~EPX;  //complement 
assign ERW =  DIO & CAC  ; 
assign erw = ~ERW;  //complement 
assign ERX =  DIP & CAB  ; 
assign erx = ~ERX;  //complement 
assign ERP =  DIH & CAJ  ; 
assign erp = ~ERP;  //complement 
assign CAA = ~caa;  //complement 
assign cab = ~CAB;  //complement 
assign cac = ~CAC;  //complement 
assign fmp = ~FMP;  //complement 
assign FNP = ~fnp;  //complement 
assign foq = ~FOQ;  //complement 
assign FPQ = ~fpq;  //complement 
assign fqp = ~FQP;  //complement 
assign OGP = ~ogp;  //complement 
assign din = ~DIN;  //complement 
assign dio = ~DIO;  //complement 
assign dip = ~DIP;  //complement 
assign ENR =  DIJ & CAF  ; 
assign enr = ~ENR;  //complement 
assign ENS =  DIK & CAE  ; 
assign ens = ~ENS;  //complement 
assign ENT =  DIL & CAD  ; 
assign ent = ~ENT;  //complement 
assign EPS =  DIK & CAF  ; 
assign eps = ~EPS;  //complement 
assign EPT =  DIL & CAE  ; 
assign ept = ~EPT;  //complement 
assign ERV =  DIN & CAD  ; 
assign erv = ~ERV;  //complement 
assign ERT =  DIL & CAF  ; 
assign ert = ~ERT;  //complement 
assign ERU =  DIM & CAE  ; 
assign eru = ~ERU;  //complement 
assign cad = ~CAD;  //complement 
assign cae = ~CAE;  //complement 
assign caf = ~CAF;  //complement 
assign fmo = ~FMO;  //complement 
assign FNO = ~fno;  //complement 
assign fop = ~FOP;  //complement 
assign FPP = ~fpp;  //complement 
assign fqo = ~FQO;  //complement 
assign OGO = ~ogo;  //complement 
assign dij = ~DIJ;  //complement 
assign dik = ~DIK;  //complement 
assign dil = ~DIL;  //complement 
assign dim = ~DIM;  //complement 
assign ENO =  DEG & CAI  ; 
assign eno = ~ENO;  //complement 
assign ENP =  DIH & CAH  ; 
assign enp = ~ENP;  //complement 
assign ENQ =  DII & CAG  ; 
assign enq = ~ENQ;  //complement 
assign EPP =  DIH & CAI  ; 
assign epp = ~EPP;  //complement 
assign EPQ =  DII & CAH  ; 
assign epq = ~EPQ;  //complement 
assign EPR =  DIJ & CAG  ; 
assign epr = ~EPR;  //complement 
assign ERQ =  DII & CAI  ; 
assign erq = ~ERQ;  //complement 
assign ERR =  DIJ & CAH  ; 
assign err = ~ERR;  //complement 
assign ERS =  DIK & CAG  ; 
assign ers = ~ERS;  //complement 
assign cag = ~CAG;  //complement 
assign cah = ~CAH;  //complement 
assign cai = ~CAI;  //complement 
assign fmn = ~FMN;  //complement 
assign FNN = ~fnn;  //complement 
assign foo = ~FOO;  //complement 
assign FPO = ~fpo;  //complement 
assign fqn = ~FQN;  //complement 
assign OGN = ~ogn;  //complement 
assign dif = ~DIF;  //complement 
assign dig = ~DIG;  //complement 
assign dih = ~DIH;  //complement 
assign dii = ~DII;  //complement 
assign ENL =  DID & CAL  ; 
assign enl = ~ENL;  //complement 
assign ENM =  DIE & CAK  ; 
assign enm = ~ENM;  //complement 
assign ENN =  DIF & CAJ  ; 
assign enn = ~ENN;  //complement 
assign EPM =  DIE & CAL  ; 
assign epm = ~EPM;  //complement 
assign EPN =  DIF & CAK  ; 
assign epn = ~EPN;  //complement 
assign EPO =  DIG & CAJ  ; 
assign epo = ~EPO;  //complement 
assign EPU =  DIM & CAD  ; 
assign epu = ~EPU;  //complement 
assign ERN =  DIF & CAL  ; 
assign ern = ~ERN;  //complement 
assign ERO =  DIG & CAK  ; 
assign ero = ~ERO;  //complement 
assign caj = ~CAJ;  //complement 
assign cak = ~CAK;  //complement 
assign cal = ~CAL;  //complement 
assign fmm = ~FMM;  //complement 
assign FNM = ~fnm;  //complement 
assign fon = ~FON;  //complement 
assign FPN = ~fpn;  //complement 
assign fqm = ~FQM;  //complement 
assign OGM = ~ogm;  //complement 
assign dic = ~DIC;  //complement 
assign did = ~DID;  //complement 
assign die = ~DIE;  //complement 
assign faj = ~FAJ;  //complement 
assign FBJ = ~fbj;  //complement 
assign fck = ~FCK;  //complement 
assign FDK = ~fdk;  //complement 
assign fel = ~FEL;  //complement 
assign FFL = ~ffl;  //complement 
assign fgk = ~FGK;  //complement 
assign FHK = ~fhk;  //complement 
assign EBC =  DEK & CDO  ; 
assign ebc = ~EBC;  //complement 
assign EBD =  DEL & CDN  ; 
assign ebd = ~EBD;  //complement 
assign EBE =  DEM & CDM  ; 
assign ebe = ~EBE;  //complement 
assign EDD =  DEL & CDO  ; 
assign edd = ~EDD;  //complement 
assign EDE =  DEM & CDN  ; 
assign ede = ~EDE;  //complement 
assign EDF =  DEN & CDM  ; 
assign edf = ~EDF;  //complement 
assign EFE =  DEM & CDO  ; 
assign efe = ~EFE;  //complement 
assign EFF =  DEN & CDN  ; 
assign eff = ~EFF;  //complement 
assign EFG =  DEO & CDM  ; 
assign efg = ~EFG;  //complement 
assign EHF =  DEN & CDO  ; 
assign ehf = ~EHF;  //complement 
assign EHG =  DEO & CDN  ; 
assign ehg = ~EHG;  //complement 
assign EHH =  DEP & CDM  ; 
assign ehh = ~EHH;  //complement 
assign fai = ~FAI;  //complement 
assign FBI = ~fbi;  //complement 
assign EEW =  DEG & CEE  ; 
assign eew = ~EEW;  //complement 
assign EEX =  DEH & CED  ; 
assign eex = ~EEX;  //complement 
assign fek = ~FEK;  //complement 
assign FFK = ~ffk;  //complement 
assign fgj = ~FGJ;  //complement 
assign FHJ = ~fhj;  //complement 
assign EAX =  DEH & CEB  ; 
assign eax = ~EAX;  //complement 
assign EBA =  DEI & CEA  ; 
assign eba = ~EBA;  //complement 
assign EBB =  DEJ & CDP  ; 
assign ebb = ~EBB;  //complement 
assign EDA =  DEI & CEB  ; 
assign eda = ~EDA;  //complement 
assign EDB =  DEJ & CEA  ; 
assign edb = ~EDB;  //complement 
assign EDC =  DEK & CDP  ; 
assign edc = ~EDC;  //complement 
assign EFB =  DEJ & CEB  ; 
assign efb = ~EFB;  //complement 
assign EFC =  DEK & CEA  ; 
assign efc = ~EFC;  //complement 
assign EFD =  DEL & CDP  ; 
assign efd = ~EFD;  //complement 
assign EHC =  DEK & CEB  ; 
assign ehc = ~EHC;  //complement 
assign EHD =  DEL & CEA  ; 
assign ehd = ~EHD;  //complement 
assign EHE =  DEM & CDP  ; 
assign ehe = ~EHE;  //complement 
assign fah = ~FAH;  //complement 
assign FBH = ~fbh;  //complement 
assign fci = ~FCI;  //complement 
assign FDI = ~fdi;  //complement 
assign fej = ~FEJ;  //complement 
assign FFJ = ~ffj;  //complement 
assign fgi = ~FGI;  //complement 
assign FHI = ~fhi;  //complement 
assign EAU =  DEE & CEE  ; 
assign eau = ~EAU;  //complement 
assign EAV =  DEF & CED  ; 
assign eav = ~EAV;  //complement 
assign EAW =  DEG & CEC  ; 
assign eaw = ~EAW;  //complement 
assign ECV =  DEF & CEE  ; 
assign ecv = ~ECV;  //complement 
assign ECW =  DEG & CED  ; 
assign ecw = ~ECW;  //complement 
assign ECX =  DEH & CEC  ; 
assign ecx = ~ECX;  //complement 
assign EFA =  DEI & CEC  ; 
assign efa = ~EFA;  //complement 
assign EGX =  DEH & CEE  ; 
assign egx = ~EGX;  //complement 
assign EHA =  DEI & CED  ; 
assign eha = ~EHA;  //complement 
assign EHB =  DEJ & CEC  ; 
assign ehb = ~EHB;  //complement 
assign fag = ~FAG;  //complement 
assign FBG = ~fbg;  //complement 
assign fch = ~FCH;  //complement 
assign FDH = ~fdh;  //complement 
assign fcj = ~FCJ;  //complement 
assign FDJ = ~fdj;  //complement 
assign fgh = ~FGH;  //complement 
assign FHH = ~fhh;  //complement 
assign EAR =  DEB & CEH  ; 
assign ear = ~EAR;  //complement 
assign EAS =  DEC & CEG  ; 
assign eas = ~EAS;  //complement 
assign EAT =  DED & CEF  ; 
assign eat = ~EAT;  //complement 
assign ECS =  DEC & CEH  ; 
assign ecs = ~ECS;  //complement 
assign ECT =  DED & CEG  ; 
assign ect = ~ECT;  //complement 
assign ECU =  DEE & CEF  ; 
assign ecu = ~ECU;  //complement 
assign EEU =  DEE & CEG  ; 
assign eeu = ~EEU;  //complement 
assign EET =  DED & CEH  ; 
assign eet = ~EET;  //complement 
assign EEV =  DEF & CEF  ; 
assign eev = ~EEV;  //complement 
assign EGU =  DEE & CEH  ; 
assign egu = ~EGU;  //complement 
assign EGV =  DEF & CEG  ; 
assign egv = ~EGV;  //complement 
assign EGW =  DEG & CEF  ; 
assign egw = ~EGW;  //complement 
assign fil = ~FIL;  //complement 
assign FJL = ~fjl;  //complement 
assign DEN = ~den;  //complement 
assign DEO = ~deo;  //complement 
assign DEP = ~dep;  //complement 
assign DFA = ~dfa;  //complement 
assign fkm = ~FKM;  //complement 
assign FLM = ~flm;  //complement 
assign EJG =  DEO & CDO  ; 
assign ejg = ~EJG;  //complement 
assign EJH =  DEP & CDN  ; 
assign ejh = ~EJH;  //complement 
assign EJI =  DFA & CDM  ; 
assign eji = ~EJI;  //complement 
assign dhk = ~DHK;  //complement 
assign dhl = ~DHL;  //complement 
assign cdm = ~CDM;  //complement 
assign cdn = ~CDN;  //complement 
assign cdo = ~CDO;  //complement 
assign ELH =  DHP & CAO  ; 
assign elh = ~ELH;  //complement 
assign ELI =  DIA & CAN  ; 
assign eli = ~ELI;  //complement 
assign ELJ =  DFB & CAM  ; 
assign elj = ~ELJ;  //complement 
assign fii = ~FII;  //complement 
assign FJI = ~fji;  //complement 
assign fik = ~FIK;  //complement 
assign FJK = ~fjk;  //complement 
assign dej = ~DEJ;  //complement 
assign dek = ~DEK;  //complement 
assign del = ~DEL;  //complement 
assign dem = ~DEM;  //complement 
assign fkl = ~FKL;  //complement 
assign FLL = ~fll;  //complement 
assign EJD =  DEL & CEB  ; 
assign ejd = ~EJD;  //complement 
assign EJE =  DEM & CEA  ; 
assign eje = ~EJE;  //complement 
assign EJF =  DEN & CDP  ; 
assign ejf = ~EJF;  //complement 
assign obb = ~OBB;  //complement 
assign cdp = ~CDP;  //complement 
assign cea = ~CEA;  //complement 
assign ceb = ~CEB;  //complement 
assign ELE =  DHM & CBB  ; 
assign ele = ~ELE;  //complement 
assign ELF =  DHN & CBA  ; 
assign elf = ~ELF;  //complement 
assign ELG =  DHO & CAP  ; 
assign elg = ~ELG;  //complement 
assign fij = ~FIJ;  //complement 
assign FJJ = ~fjj;  //complement 
assign def = ~DEF;  //complement 
assign deg = ~DEG;  //complement 
assign deh = ~DEH;  //complement 
assign dei = ~DEI;  //complement 
assign fkk = ~FKK;  //complement 
assign FLK = ~flk;  //complement 
assign EJA =  DEI & CEE  ; 
assign eja = ~EJA;  //complement 
assign EJB =  DEJ & CED  ; 
assign ejb = ~EJB;  //complement 
assign EJC =  DEK & CEC  ; 
assign ejc = ~EJC;  //complement 
assign cec = ~CEC;  //complement 
assign ced = ~CED;  //complement 
assign cee = ~CEE;  //complement 
assign ELC =  DHK & CBD  ; 
assign elc = ~ELC;  //complement 
assign ELB =  DHJ & CBE  ; 
assign elb = ~ELB;  //complement 
assign ELD =  DHL & CBC  ; 
assign eld = ~ELD;  //complement 
assign cef = ~CEF;  //complement 
assign ceg = ~CEG;  //complement 
assign ceh = ~CEH;  //complement 
assign fei = ~FEI;  //complement 
assign FFI = ~ffi;  //complement 
assign deb = ~DEB;  //complement 
assign dec = ~DEC;  //complement 
assign ded = ~DED;  //complement 
assign dee = ~DEE;  //complement 
assign fkj = ~FKJ;  //complement 
assign FLJ = ~flj;  //complement 
assign EIV =  DEF & CEH  ; 
assign eiv = ~EIV;  //complement 
assign EIW =  DEG & CEG  ; 
assign eiw = ~EIW;  //complement 
assign EIX =  DEH & CEF  ; 
assign eix = ~EIX;  //complement 
assign aad = ~AAD;  //complement 
assign EKW =  DHG & CBH  ; 
assign ekw = ~EKW;  //complement 
assign EKX =  DHH & CBG  ; 
assign ekx = ~EKX;  //complement 
assign ELA =  DHI & CBF  ; 
assign ela = ~ELA;  //complement 
assign fml = ~FML;  //complement 
assign FNL = ~fnl;  //complement 
assign fom = ~FOM;  //complement 
assign FPM = ~fpm;  //complement 
assign fql = ~FQL;  //complement 
assign OGL = ~ogl;  //complement 
assign DFB = ~dfb;  //complement 
assign DFC = ~dfc;  //complement 
assign DFD = ~dfd;  //complement 
assign DFE = ~dfe;  //complement 
assign ENI =  DIA & CAO  ; 
assign eni = ~ENI;  //complement 
assign ENK =  DFC & CAM  ; 
assign enk = ~ENK;  //complement 
assign ENJ =  DFB & CAN  ; 
assign enj = ~ENJ;  //complement 
assign EPJ =  DFB & CAO  ; 
assign epj = ~EPJ;  //complement 
assign EPK =  DFC & CAN  ; 
assign epk = ~EPK;  //complement 
assign EPL =  DFD & CAM  ; 
assign epl = ~EPL;  //complement 
assign ERK =  DFC & CAO  ; 
assign erk = ~ERK;  //complement 
assign ERL =  DFD & CAN  ; 
assign erl = ~ERL;  //complement 
assign ERM =  DFE & CAM  ; 
assign erm = ~ERM;  //complement 
assign cam = ~CAM;  //complement 
assign can = ~CAN;  //complement 
assign cao = ~CAO;  //complement 
assign fmk = ~FMK;  //complement 
assign FNK = ~fnk;  //complement 
assign fol = ~FOL;  //complement 
assign FPL = ~fpl;  //complement 
assign fqk = ~FQK;  //complement 
assign OGK = ~ogk;  //complement 
assign DHN = ~dhn;  //complement 
assign DHO = ~dho;  //complement 
assign DHP = ~dhp;  //complement 
assign DIA = ~dia;  //complement 
assign ENF =  DHN & CBB  ; 
assign enf = ~ENF;  //complement 
assign ENG =  DHO & CBA  ; 
assign eng = ~ENG;  //complement 
assign ENH =  DHP & CAP  ; 
assign enh = ~ENH;  //complement 
assign EPG =  DHO & CBB  ; 
assign epg = ~EPG;  //complement 
assign EPH =  DHP & CBA  ; 
assign eph = ~EPH;  //complement 
assign EPI =  DIA & CAP  ; 
assign epi = ~EPI;  //complement 
assign ERH =  DHP & CBB  ; 
assign erh = ~ERH;  //complement 
assign ERI =  DIA & CBA  ; 
assign eri = ~ERI;  //complement 
assign ERJ =  DFB & CAP  ; 
assign erj = ~ERJ;  //complement 
assign cap = ~CAP;  //complement 
assign cba = ~CBA;  //complement 
assign cbb = ~CBB;  //complement 
assign fmj = ~FMJ;  //complement 
assign FNJ = ~fnj;  //complement 
assign fok = ~FOK;  //complement 
assign FPK = ~fpk;  //complement 
assign fqj = ~FQJ;  //complement 
assign OGJ = ~ogj;  //complement 
assign dhj = ~DHJ;  //complement 
assign dhm = ~DHM;  //complement 
assign ENC =  DHK & CBE  ; 
assign enc = ~ENC;  //complement 
assign ENDD  =  DHL & CBD  ; 
assign endd = ~ENDD ;  //complement 
assign ENE =  DHM & CBC  ; 
assign ene = ~ENE;  //complement 
assign EPD =  DHL & CBE  ; 
assign epd = ~EPD;  //complement 
assign EPE =  DHM & CBD  ; 
assign epe = ~EPE;  //complement 
assign EPF =  DHN & CBC  ; 
assign epf = ~EPF;  //complement 
assign ERE =  DHM & CBE  ; 
assign ere = ~ERE;  //complement 
assign ERF =  DHN & CBD  ; 
assign erf = ~ERF;  //complement 
assign ERG =  DHO & CBC  ; 
assign erg = ~ERG;  //complement 
assign cbc = ~CBC;  //complement 
assign cbd = ~CBD;  //complement 
assign cbe = ~CBE;  //complement 
assign fmi = ~FMI;  //complement 
assign FNI = ~fni;  //complement 
assign foj = ~FOJ;  //complement 
assign FPJ = ~fpj;  //complement 
assign fqi = ~FQI;  //complement 
assign OGI = ~ogi;  //complement 
assign tra = ~TRA;  //complement 
assign dhg = ~DHG;  //complement 
assign dhh = ~DHH;  //complement 
assign dhi = ~DHI;  //complement 
assign EMX =  DHH & CBH  ; 
assign emx = ~EMX;  //complement 
assign ENA =  DHI & CBG  ; 
assign ena = ~ENA;  //complement 
assign ENB =  DHJ & CBF  ; 
assign enb = ~ENB;  //complement 
assign EPA =  DHI & CBH  ; 
assign epa = ~EPA;  //complement 
assign EPB =  DHJ & CBG  ; 
assign epb = ~EPB;  //complement 
assign EPC =  DHK & CBF  ; 
assign epc = ~EPC;  //complement 
assign ERB =  DHJ & CBH  ; 
assign erb = ~ERB;  //complement 
assign ERC =  DHK & CBG  ; 
assign erc = ~ERC;  //complement 
assign ERD =  DHL & CBF  ; 
assign erd = ~ERD;  //complement 
assign cbf = ~CBF;  //complement 
assign cbg = ~CBG;  //complement 
assign cbh = ~CBH;  //complement 
assign GCG =  FBJ & fbn & fbf  |  fbj & FBN & fbf  |  fbj & fbn & FBF  |  FBJ & FBN & FBF  ; 
assign gcg = ~GCG; //complement 
assign gdg =  FBJ & fbn & fbf  |  fbj & FBN & fbf  |  fbj & fbn & FBF  |  fbj & fbn & fbf  ; 
assign GDG = ~gdg;  //complement 
assign GEH =  FDK & fdo & fdg  |  fdk & FDO & fdg  |  fdk & fdo & FDG  |  FDK & FDO & FDG  ; 
assign geh = ~GEH; //complement 
assign gfh =  FDK & fdo & fdg  |  fdk & FDO & fdg  |  fdk & fdo & FDG  |  fdk & fdo & fdg  ; 
assign GFH = ~gfh;  //complement 
assign GGG =  FFL & ffp & ffh  |  ffl & FFP & ffh  |  ffl & ffp & FFH  |  FFL & FFP & FFH  ; 
assign ggg = ~GGG; //complement 
assign ghg =  FFL & ffp & ffh  |  ffl & FFP & ffh  |  ffl & ffp & FFH  |  ffl & ffp & ffh  ; 
assign GHG = ~ghg;  //complement 
assign GIH =  FHO & fhk & fhg  |  fho & FHK & fhg  |  fho & fhk & FHG  |  FHO & FHK & FHG  ; 
assign gih = ~GIH; //complement 
assign gjh =  FHO & fhk & fhg  |  fho & FHK & fhg  |  fho & fhk & FHG  |  fho & fhk & fhg  ; 
assign GJH = ~gjh;  //complement 
assign GAD =  FAN & faj & fai  |  fan & FAJ & fai  |  fan & faj & FAI  |  FAN & FAJ & FAI  ; 
assign gad = ~GAD; //complement 
assign gbd =  FAN & faj & fai  |  fan & FAJ & fai  |  fan & faj & FAI  |  fan & faj & fai  ; 
assign GBD = ~gbd;  //complement 
assign GCD =  FCO & fcj & fck  |  fco & FCJ & fck  |  fco & fcj & FCK  |  FCO & FCJ & FCK  ; 
assign gcd = ~GCD; //complement 
assign gdd =  FCO & fcj & fck  |  fco & FCJ & fck  |  fco & fcj & FCK  |  fco & fcj & fck  ; 
assign GDD = ~gdd;  //complement 
assign GEE =  FEP & fel & fek  |  fep & FEL & fek  |  fep & fel & FEK  |  FEP & FEL & FEK  ; 
assign gee = ~GEE; //complement 
assign gfe =  FEP & fel & fek  |  fep & FEL & fek  |  fep & fel & FEK  |  fep & fel & fek  ; 
assign GFE = ~gfe;  //complement 
assign GGD =  FGO & fgk & fgj  |  fgo & FGK & fgj  |  fgo & fgk & FGJ  |  FGO & FGK & FGJ  ; 
assign ggd = ~GGD; //complement 
assign ghd =  FGO & fgk & fgj  |  fgo & FGK & fgj  |  fgo & fgk & FGJ  |  fgo & fgk & fgj  ; 
assign GHD = ~ghd;  //complement 
assign hcc = ~HCC;  //complement 
assign HDC = ~hdc;  //complement 
assign hcb = ~HCB;  //complement 
assign HDB = ~hdb;  //complement 
assign heb = ~HEB;  //complement 
assign HFB = ~hfb;  //complement 
assign hgb = ~HGB;  //complement 
assign HHB = ~hhb;  //complement 
assign hih = ~HIH;  //complement 
assign GCH =  FBH & fbi & fbm  |  fbh & FBI & fbm  |  fbh & fbi & FBM  |  FBH & FBI & FBM  ; 
assign gch = ~GCH; //complement 
assign gdh =  FBH & fbi & fbm  |  fbh & FBI & fbm  |  fbh & fbi & FBM  |  fbh & fbi & fbm  ; 
assign GDH = ~gdh;  //complement 
assign GEI =  FDI & fdj & fdn  |  fdi & FDJ & fdn  |  fdi & fdj & FDN  |  FDI & FDJ & FDN  ; 
assign gei = ~GEI; //complement 
assign gfi =  FDI & fdj & fdn  |  fdi & FDJ & fdn  |  fdi & fdj & FDN  |  fdi & fdj & fdn  ; 
assign GFI = ~gfi;  //complement 
assign GGH =  FFO & ffj & ffk  |  ffo & FFJ & ffk  |  ffo & ffj & FFK  |  FFO & FFJ & FFK  ; 
assign ggh = ~GGH; //complement 
assign ghh =  FFO & ffj & ffk  |  ffo & FFJ & ffk  |  ffo & ffj & FFK  |  ffo & ffj & ffk  ; 
assign GHH = ~ghh;  //complement 
assign GII =  FHN & fhi & fhj  |  fhn & FHI & fhj  |  fhn & fhi & FHJ  |  FHN & FHI & FHJ  ; 
assign gii = ~GII; //complement 
assign gji =  FHN & fhi & fhj  |  fhn & FHI & fhj  |  fhn & fhi & FHJ  |  fhn & fhi & fhj  ; 
assign GJI = ~gji;  //complement 
assign GAC =  FAL & fam & fah  |  fal & FAM & fah  |  fal & fam & FAH  |  FAL & FAM & FAH  ; 
assign gac = ~GAC; //complement 
assign gbc =  FAL & fam & fah  |  fal & FAM & fah  |  fal & fam & FAH  |  fal & fam & fah  ; 
assign GBC = ~gbc;  //complement 
assign GCC =  FCM & fcn & fci  |  fcm & FCN & fci  |  fcm & fcn & FCI  |  FCM & FCN & FCI  ; 
assign gcc = ~GCC; //complement 
assign gdc =  FCM & fcn & fci  |  fcm & FCN & fci  |  fcm & fcn & FCI  |  fcm & fcn & fci  ; 
assign GDC = ~gdc;  //complement 
assign GED =  FEN & feo & fej  |  fen & FEO & fej  |  fen & feo & FEJ  |  FEN & FEO & FEJ  ; 
assign ged = ~GED; //complement 
assign gfd =  FEN & feo & fej  |  fen & FEO & fej  |  fen & feo & FEJ  |  fen & feo & fej  ; 
assign GFD = ~gfd;  //complement 
assign GGC =  FGN & fgm & fgi  |  fgn & FGM & fgi  |  fgn & fgm & FGI  |  FGN & FGM & FGI  ; 
assign ggc = ~GGC; //complement 
assign ghc =  FGN & fgm & fgi  |  fgn & FGM & fgi  |  fgn & fgm & FGI  |  fgn & fgm & fgi  ; 
assign GHC = ~ghc;  //complement 
assign hab = ~HAB;  //complement 
assign HBB = ~hbb;  //complement 
assign hed = ~HED;  //complement 
assign HFD = ~hfd;  //complement 
assign hgd = ~HGD;  //complement 
assign HHD = ~hhd;  //complement 
assign hid = ~HID;  //complement 
assign HJD = ~hjd;  //complement 
assign GCI =  FBK & fbl & fbg  |  fbk & FBL & fbg  |  fbk & fbl & FBG  |  FBK & FBL & FBG  ; 
assign gci = ~GCI; //complement 
assign gdi =  FBK & fbl & fbg  |  fbk & FBL & fbg  |  fbk & fbl & FBG  |  fbk & fbl & fbg  ; 
assign GDI = ~gdi;  //complement 
assign GEJ =  FDL & fdm & fdh  |  fdl & FDM & fdh  |  fdl & fdm & FDH  |  FDL & FDM & FDH  ; 
assign gej = ~GEJ; //complement 
assign gfj =  FDL & fdm & fdh  |  fdl & FDM & fdh  |  fdl & fdm & FDH  |  fdl & fdm & fdh  ; 
assign GFJ = ~gfj;  //complement 
assign GGI =  FFM & ffn & ffi  |  ffm & FFN & ffi  |  ffm & ffn & FFI  |  FFM & FFN & FFI  ; 
assign ggi = ~GGI; //complement 
assign ghi =  FFM & ffn & ffi  |  ffm & FFN & ffi  |  ffm & ffn & FFI  |  ffm & ffn & ffi  ; 
assign GHI = ~ghi;  //complement 
assign GIJ =  FHL & fhm & fhh  |  fhl & FHM & fhh  |  fhl & fhm & FHH  |  FHL & FHM & FHH  ; 
assign gij = ~GIJ; //complement 
assign gjj =  FHL & fhm & fhh  |  fhl & FHM & fhh  |  fhl & fhm & FHH  |  fhl & fhm & fhh  ; 
assign GJJ = ~gjj;  //complement 
assign GAB =  FAG & fak & fac  |  fag & FAK & fac  |  fag & fak & FAC  |  FAG & FAK & FAC  ; 
assign gab = ~GAB; //complement 
assign gbb =  FAG & fak & fac  |  fag & FAK & fac  |  fag & fak & FAC  |  fag & fak & fac  ; 
assign GBB = ~gbb;  //complement 
assign GCB =  FCH & fcl & fcd  |  fch & FCL & fcd  |  fch & fcl & FCD  |  FCH & FCL & FCD  ; 
assign gcb = ~GCB; //complement 
assign gdb =  FCH & fcl & fcd  |  fch & FCL & fcd  |  fch & fcl & FCD  |  fch & fcl & fcd  ; 
assign GDB = ~gdb;  //complement 
assign GEC =  FEM & fei & fee  |  fem & FEI & fee  |  fem & fei & FEE  |  FEM & FEI & FEE  ; 
assign gec = ~GEC; //complement 
assign gfc =  FEM & fei & fee  |  fem & FEI & fee  |  fem & fei & FEE  |  fem & fei & fee  ; 
assign GFC = ~gfc;  //complement 
assign GGB =  FGL & fgh & fgd  |  fgl & FGH & fgd  |  fgl & fgh & FGD  |  FGL & FGH & FGD  ; 
assign ggb = ~GGB; //complement 
assign ghb =  FGL & fgh & fgd  |  fgl & FGH & fgd  |  fgl & fgh & FGD  |  fgl & fgh & fgd  ; 
assign GHB = ~ghb;  //complement 
assign GKH =  FJP & fjl & fjh  |  fjp & FJL & fjh  |  fjp & fjl & FJH  |  FJP & FJL & FJH  ; 
assign gkh = ~GKH; //complement 
assign glh =  FJP & fjl & fjh  |  fjp & FJL & fjh  |  fjp & fjl & FJH  |  fjp & fjl & fjh  ; 
assign GLH = ~glh;  //complement 
assign GMH =  FLQ & flm & fli  |  flq & FLM & fli  |  flq & flm & FLI  |  FLQ & FLM & FLI  ; 
assign gmh = ~GMH; //complement 
assign gnh =  FLQ & flm & fli  |  flq & FLM & fli  |  flq & flm & FLI  |  flq & flm & fli  ; 
assign GNH = ~gnh;  //complement 
assign GOI =  FNL & fnp & fnh  |  fnl & FNP & fnh  |  fnl & fnp & FNH  |  FNL & FNP & FNH  ; 
assign goi = ~GOI; //complement 
assign gpi =  FNL & fnp & fnh  |  fnl & FNP & fnh  |  fnl & fnp & FNH  |  fnl & fnp & fnh  ; 
assign GPI = ~gpi;  //complement 
assign GIE =  FIK & fil & fip  |  fik & FIL & fip  |  fik & fil & FIP  |  FIK & FIL & FIP  ; 
assign gie = ~GIE; //complement 
assign gje =  FIK & fil & fip  |  fik & FIL & fip  |  fik & fil & FIP  |  fik & fil & fip  ; 
assign GJE = ~gje;  //complement 
assign GKE =  FKQ & fkm & fkl  |  fkq & FKM & fkl  |  fkq & fkm & FKL  |  FKQ & FKM & FKL  ; 
assign gke = ~GKE; //complement 
assign gle =  FKQ & fkm & fkl  |  fkq & FKM & fkl  |  fkq & fkm & FKL  |  fkq & fkm & fkl  ; 
assign GLE = ~gle;  //complement 
assign GME =  FMK & fml & fmp  |  fmk & FML & fmp  |  fmk & fml & FMP  |  FMK & FML & FMP  ; 
assign gme = ~GME; //complement 
assign gne =  FMK & fml & fmp  |  fmk & FML & fmp  |  fmk & fml & FMP  |  fmk & fml & fmp  ; 
assign GNE = ~gne;  //complement 
assign hib = ~HIB;  //complement 
assign HJB = ~hjb;  //complement 
assign hmb = ~HMB;  //complement 
assign HNB = ~hnb;  //complement 
assign hob = ~HOB;  //complement 
assign HPB = ~hpb;  //complement 
assign GKI =  FJO & fjj & fjk  |  fjo & FJJ & fjk  |  fjo & fjj & FJK  |  FJO & FJJ & FJK  ; 
assign gki = ~GKI; //complement 
assign gli =  FJO & fjj & fjk  |  fjo & FJJ & fjk  |  fjo & fjj & FJK  |  fjo & fjj & fjk  ; 
assign GLI = ~gli;  //complement 
assign hkb = ~HKB;  //complement 
assign HLB = ~hlb;  //complement 
assign GMI =  FLP & flk & fll  |  flp & FLK & fll  |  flp & flk & FLL  |  FLP & FLK & FLL  ; 
assign gmi = ~GMI; //complement 
assign gni =  FLP & flk & fll  |  flp & FLK & fll  |  flp & flk & FLL  |  flp & flk & fll  ; 
assign GNI = ~gni;  //complement 
assign GOJ =  FNJ & fnk & fno  |  fnj & FNK & fno  |  fnj & fnk & FNO  |  FNJ & FNK & FNO  ; 
assign goj = ~GOJ; //complement 
assign gpj =  FNJ & fnk & fno  |  fnj & FNK & fno  |  fnj & fnk & FNO  |  fnj & fnk & fno  ; 
assign GPJ = ~gpj;  //complement 
assign GID =  FIN & fio & fij  |  fin & FIO & fij  |  fin & fio & FIJ  |  FIN & FIO & FIJ  ; 
assign gid = ~GID; //complement 
assign gjd =  FIN & fio & fij  |  fin & FIO & fij  |  fin & fio & FIJ  |  fin & fio & fij  ; 
assign GJD = ~gjd;  //complement 
assign hkg = ~HKG;  //complement 
assign HLG = ~hlg;  //complement 
assign GKD =  FKO & fkp & fkk  |  fko & FKP & fkk  |  fko & fkp & FKK  |  FKO & FKP & FKK  ; 
assign gkd = ~GKD; //complement 
assign gld =  FKO & fkp & fkk  |  fko & FKP & fkk  |  fko & fkp & FKK  |  fko & fkp & fkk  ; 
assign GLD = ~gld;  //complement 
assign GMD =  FMN & fmo & fmj  |  fmn & FMO & fmj  |  fmn & fmo & FMJ  |  FMN & FMO & FMJ  ; 
assign gmd = ~GMD; //complement 
assign gnd =  FMN & fmo & fmj  |  fmn & FMO & fmj  |  fmn & fmo & FMJ  |  fmn & fmo & fmj  ; 
assign GND = ~gnd;  //complement 
assign hkd = ~HKD;  //complement 
assign HLD = ~hld;  //complement 
assign hmd = ~HMD;  //complement 
assign HND = ~hnd;  //complement 
assign hod = ~HOD;  //complement 
assign HPD = ~hpd;  //complement 
assign GKJ =  FJM & fjn & fji  |  fjm & FJN & fji  |  fjm & fjn & FJI  |  FJM & FJN & FJI  ; 
assign gkj = ~GKJ; //complement 
assign glj =  FJM & fjn & fji  |  fjm & FJN & fji  |  fjm & fjn & FJI  |  fjm & fjn & fji  ; 
assign GLJ = ~glj;  //complement 
assign GMJ =  FLN & flo & flj  |  fln & FLO & flj  |  fln & flo & FLJ  |  FLN & FLO & FLJ  ; 
assign gmj = ~GMJ; //complement 
assign gnj =  FLN & flo & flj  |  fln & FLO & flj  |  fln & flo & FLJ  |  fln & flo & flj  ; 
assign GNJ = ~gnj;  //complement 
assign GOK =  FNI & fnm & fnn  |  fni & FNM & fnn  |  fni & fnm & FNN  |  FNI & FNM & FNN  ; 
assign gok = ~GOK; //complement 
assign gpk =  FNI & fnm & fnn  |  fni & FNM & fnn  |  fni & fnm & FNN  |  fni & fnm & fnn  ; 
assign GPK = ~gpk;  //complement 
assign GIC =  FIM & fii & fie  |  fim & FII & fie  |  fim & fii & FIE  |  FIM & FII & FIE  ; 
assign gic = ~GIC; //complement 
assign gjc =  FIM & fii & fie  |  fim & FII & fie  |  fim & fii & FIE  |  fim & fii & fie  ; 
assign GJC = ~gjc;  //complement 
assign GKC =  FKN & fkj & fkf  |  fkn & FKJ & fkf  |  fkn & fkj & FKF  |  FKN & FKJ & FKF  ; 
assign gkc = ~GKC; //complement 
assign glc =  FKN & fkj & fkf  |  fkn & FKJ & fkf  |  fkn & fkj & FKF  |  fkn & fkj & fkf  ; 
assign GLC = ~glc;  //complement 
assign GMC =  FMM & fmi & fme  |  fmm & FMI & fme  |  fmm & fmi & FME  |  FMM & FMI & FME  ; 
assign gmc = ~GMC; //complement 
assign gnc =  FMM & fmi & fme  |  fmm & FMI & fme  |  fmm & fmi & FME  |  fmm & fmi & fme  ; 
assign GNC = ~gnc;  //complement 
assign GQH =  FPM & fpq & fpi  |  fpm & FPQ & fpi  |  fpm & fpq & FPI  |  FPM & FPQ & FPI  ; 
assign gqh = ~GQH; //complement 
assign grh =  FPM & fpq & fpi  |  fpm & FPQ & fpi  |  fpm & fpq & FPI  |  fpm & fpq & fpi  ; 
assign GRH = ~grh;  //complement 
assign ohh = ~OHH;  //complement 
assign OIH = ~oih;  //complement 
assign aab = ~AAB;  //complement 
assign oba = ~OBA;  //complement 
assign GOF =  FOQ & fol & fom  |  foq & FOL & fom  |  foq & fol & FOM  |  FOQ & FOL & FOM  ; 
assign gof = ~GOF; //complement 
assign gpf =  FOQ & fol & fom  |  foq & FOL & fom  |  foq & fol & FOM  |  foq & fol & fom  ; 
assign GPF = ~gpf;  //complement 
assign GQE =  FQK & fql & fqp  |  fqk & FQL & fqp  |  fqk & fql & FQP  |  FQK & FQL & FQP  ; 
assign gqe = ~GQE; //complement 
assign gre =  FQK & fql & fqp  |  fqk & FQL & fqp  |  fqk & fql & FQP  |  fqk & fql & fqp  ; 
assign GRE = ~gre;  //complement 
assign bda = ~BDA;  //complement 
assign bdb = ~BDB;  //complement 
assign bea = ~BEA;  //complement 
assign beb = ~BEB;  //complement 
assign oab = ~OAB;  //complement 
assign hqb = ~HQB;  //complement 
assign OHB = ~ohb;  //complement 
assign qga = ~QGA;  //complement 
assign qha = ~QHA;  //complement 
assign qka = ~QKA;  //complement 
assign BBA = ~bba;  //complement 
assign BBB = ~bbb;  //complement 
assign bca = ~BCA;  //complement 
assign bcb = ~BCB;  //complement 
assign oda = ~ODA;  //complement 
assign oea = ~OEA;  //complement 
assign GQI =  FPK & fpl & fpp  |  fpk & FPL & fpp  |  fpk & fpl & FPP  |  FPK & FPL & FPP  ; 
assign gqi = ~GQI; //complement 
assign gri =  FPK & fpl & fpp  |  fpk & FPL & fpp  |  fpk & fpl & FPP  |  fpk & fpl & fpp  ; 
assign GRI = ~gri;  //complement 
assign ohi = ~OHI;  //complement 
assign OII = ~oii;  //complement 
assign ohk = ~OHK;  //complement 
assign baa = ~BAA;  //complement 
assign bab = ~BAB;  //complement 
assign odb = ~ODB;  //complement 
assign oeb = ~OEB;  //complement 
assign obd = ~OBD;  //complement 
assign GQD =  FQN & fqo & fqj  |  fqn & FQO & fqj  |  fqn & fqo & FQJ  |  FQN & FQO & FQJ  ; 
assign gqd = ~GQD; //complement 
assign grd =  FQN & fqo & fqj  |  fqn & FQO & fqj  |  fqn & fqo & FQJ  |  fqn & fqo & fqj  ; 
assign GRD = ~grd;  //complement 
assign bac = ~BAC;  //complement 
assign bad = ~BAD;  //complement 
assign odd = ~ODD;  //complement 
assign oed = ~OED;  //complement 
assign hqd = ~HQD;  //complement 
assign OHD = ~ohd;  //complement 
assign qra = ~QRA;  //complement 
assign qsa = ~QSA;  //complement 
assign qta = ~QTA;  //complement 
assign BBC = ~bbc;  //complement 
assign BBD = ~bbd;  //complement 
assign bcc = ~BCC;  //complement 
assign bcd = ~BCD;  //complement 
assign odc = ~ODC;  //complement 
assign oec = ~OEC;  //complement 
assign GQJ =  FPN & fpo & fpj  |  fpn & FPO & fpj  |  fpn & fpo & FPJ  |  FPN & FPO & FPJ  ; 
assign gqj = ~GQJ; //complement 
assign grj =  FPN & fpo & fpj  |  fpn & FPO & fpj  |  fpn & fpo & FPJ  |  fpn & fpo & fpj  ; 
assign GRJ = ~grj;  //complement 
assign ohj = ~OHJ;  //complement 
assign OIJ = ~oij;  //complement 
assign bdc = ~BDC;  //complement 
assign bdd = ~BDD;  //complement 
assign bec = ~BEC;  //complement 
assign bed = ~BED;  //complement 
assign oad = ~OAD;  //complement 
assign GOD =  FON & foj & fof  |  fon & FOJ & fof  |  fon & foj & FOF  |  FON & FOJ & FOF  ; 
assign god = ~GOD; //complement 
assign gpd =  FON & foj & fof  |  fon & FOJ & fof  |  fon & foj & FOF  |  fon & foj & fof  ; 
assign GPD = ~gpd;  //complement 
assign GQC =  FQM & fqi & fqe  |  fqm & FQI & fqe  |  fqm & fqi & FQE  |  FQM & FQI & FQE  ; 
assign gqc = ~GQC; //complement 
assign grc =  FQM & fqi & fqe  |  fqm & FQI & fqe  |  fqm & fqi & FQE  |  fqm & fqi & fqe  ; 
assign GRC = ~grc;  //complement 
assign aac = ~AAC;  //complement 
assign oac = ~OAC;  //complement 
assign obc = ~OBC;  //complement 
assign GOE =  FOO & fop & fok  |  foo & FOP & fok  |  foo & fop & FOK  |  FOO & FOP & FOK  ; 
assign goe = ~GOE; //complement 
assign gpe =  FOO & fop & fok  |  foo & FOP & fok  |  foo & fop & FOK  |  foo & fop & fok  ; 
assign GPE = ~gpe;  //complement 
assign kga = ~KGA;  //complement 
assign KHA = ~kha;  //complement 
assign kia = ~KIA;  //complement 
assign KJA = ~kja;  //complement 
assign JEB =  HDB & heb & hec  |  hdb & HEB & hec  |  hdb & heb & HEC  |  HDB & HEB & HEC  ; 
assign jeb = ~JEB; //complement 
assign jfb =  HDB & heb & hec  |  hdb & HEB & hec  |  hdb & heb & HEC  |  hdb & heb & hec  ; 
assign JFB = ~jfb;  //complement 
assign LIA =  KIA & kha & kic  |  kia & KHA & kic  |  kia & kha & KIC  |  KIA & KHA & KIC  ; 
assign lia = ~LIA; //complement 
assign lja =  KIA & kha & kic  |  kia & KHA & kic  |  kia & kha & KIC  |  kia & kha & kic  ; 
assign LJA = ~lja;  //complement 
assign JCA =  HCC & hcb & hba  |  hcc & HCB & hba  |  hcc & hcb & HBA  |  HCC & HCB & HBA  ; 
assign jca = ~JCA; //complement 
assign jda =  HCC & hcb & hba  |  hcc & HCB & hba  |  hcc & hcb & HBA  |  hcc & hcb & hba  ; 
assign JDA = ~jda;  //complement 
assign JGB =  HFB & hgb & hgc  |  hfb & HGB & hgc  |  hfb & hgb & HGC  |  HFB & HGB & HGC  ; 
assign jgb = ~JGB; //complement 
assign jhb =  HFB & hgb & hgc  |  hfb & HGB & hgc  |  hfb & hgb & HGC  |  hfb & hgb & hgc  ; 
assign JHB = ~jhb;  //complement 
assign JIB =  HHB & hih & hib  |  hhb & HIH & hib  |  hhb & hih & HIB  |  HHB & HIH & HIB  ; 
assign jib = ~JIB; //complement 
assign jjb =  HHB & hih & hib  |  hhb & HIH & hib  |  hhb & hih & HIB  |  hhb & hih & hib  ; 
assign JJB = ~jjb;  //complement 
assign OQJ = ~oqj;  //complement 
assign kic = ~KIC;  //complement 
assign KJC = ~kjc;  //complement 
assign kca = ~KCA;  //complement 
assign KDA = ~kda;  //complement 
assign kcb = ~KCB;  //complement 
assign nha =  MGB & mga & mfa  |  mgb & MGA & mfa  |  mgb & mga & MFA  |  mgb & mga & mfa  ; 
assign NHA = ~nha;  //complement 
assign kgc = ~KGC;  //complement 
assign KHC = ~khc;  //complement 
assign mgb = ~MGB;  //complement 
assign mia = ~MIA;  //complement 
assign MJA = ~mja;  //complement 
assign jba =  HAA & hab  |  haa & HAB  |  haa & hab  |  haa & hab  ; 
assign JBA = ~jba;  //complement 
assign JEC =  HED & hdd & heg  |  hed & HDD & heg  |  hed & hdd & HEG  |  HED & HDD & HEG  ; 
assign jec = ~JEC; //complement 
assign jfc =  HED & hdd & heg  |  hed & HDD & heg  |  hed & hdd & HEG  |  hed & hdd & heg  ; 
assign JFC = ~jfc;  //complement 
assign JGC =  HFD & hgd & hfe  |  hfd & HGD & hfe  |  hfd & hgd & HFE  |  HFD & HGD & HFE  ; 
assign jgc = ~JGC; //complement 
assign jhc =  HFD & hgd & hfe  |  hfd & HGD & hfe  |  hfd & hgd & HFE  |  hfd & hgd & hfe  ; 
assign JHC = ~jhc;  //complement 
assign JIC =  HID & hhd & hhe  |  hid & HHD & hhe  |  hid & hhd & HHE  |  HID & HHD & HHE  ; 
assign jic = ~JIC; //complement 
assign jjc =  HID & hhd & hhe  |  hid & HHD & hhe  |  hid & hhd & HHE  |  hid & hhd & hhe  ; 
assign JJC = ~jjc;  //complement 
assign kka = ~KKA;  //complement 
assign KLA = ~kla;  //complement 
assign kma = ~KMA;  //complement 
assign KNA = ~kna;  //complement 
assign mqc = ~MQC;  //complement 
assign koa = ~KOA;  //complement 
assign KPA = ~kpa;  //complement 
assign mka = ~MKA;  //complement 
assign MLA = ~mla;  //complement 
assign LMA =  KMA & kla & kmc  |  kma & KLA & kmc  |  kma & kla & KMC  |  KMA & KLA & KMC  ; 
assign lma = ~LMA; //complement 
assign lna =  KMA & kla & kmc  |  kma & KLA & kmc  |  kma & kla & KMC  |  kma & kla & kmc  ; 
assign LNA = ~lna;  //complement 
assign hmg = ~HMG;  //complement 
assign HNG = ~hng;  //complement 
assign JKB =  HJB & hkc & hkb  |  hjb & HKC & hkb  |  hjb & hkc & HKB  |  HJB & HKC & HKB  ; 
assign jkb = ~JKB; //complement 
assign jlb =  HJB & hkc & hkb  |  hjb & HKC & hkb  |  hjb & hkc & HKB  |  hjb & hkc & hkb  ; 
assign JLB = ~jlb;  //complement 
assign JMB =  HMB & hlb & hmc  |  hmb & HLB & hmc  |  hmb & hlb & HMC  |  HMB & HLB & HMC  ; 
assign jmb = ~JMB; //complement 
assign jnb =  HMB & hlb & hmc  |  hmb & HLB & hmc  |  hmb & hlb & HMC  |  hmb & hlb & hmc  ; 
assign JNB = ~jnb;  //complement 
assign JOB =  HOB & hnb & hog  |  hob & HNB & hog  |  hob & hnb & HOG  |  HOB & HNB & HOG  ; 
assign job = ~JOB; //complement 
assign jpb =  HOB & hnb & hog  |  hob & HNB & hog  |  hob & hnb & HOG  |  hob & hnb & hog  ; 
assign JPB = ~jpb;  //complement 
assign kkc = ~KKC;  //complement 
assign KLC = ~klc;  //complement 
assign kke = ~KKE;  //complement 
assign NMA =  MMA & mmc & mmb  |  mma & MMC & mmb  |  mma & mmc & MMB  |  MMA & MMC & MMB  ; 
assign nma = ~NMA; //complement 
assign nna =  MMA & mmc & mmb  |  mma & MMC & mmb  |  mma & mmc & MMB  |  mma & mmc & mmb  ; 
assign NNA = ~nna;  //complement 
assign kmc = ~KMC;  //complement 
assign KNC = ~knc;  //complement 
assign mmc = ~MMC;  //complement 
assign koc = ~KOC;  //complement 
assign KPC = ~kpc;  //complement 
assign moc = ~MOC;  //complement 
assign opk = ~OPK;  //complement 
assign OQK = ~oqk;  //complement 
assign opm = ~OPM;  //complement 
assign OQM = ~oqm;  //complement 
assign moa = ~MOA;  //complement 
assign MPA = ~mpa;  //complement 
assign mob = ~MOB;  //complement 
assign NOA =  MOA & mob & moc  |  moa & MOB & moc  |  moa & mob & MOC  |  MOA & MOB & MOC  ; 
assign noa = ~NOA; //complement 
assign npa =  MOA & mob & moc  |  moa & MOB & moc  |  moa & mob & MOC  |  moa & mob & moc  ; 
assign NPA = ~npa;  //complement 
assign JKC =  HKD & hjd & hje  |  hkd & HJD & hje  |  hkd & hjd & HJE  |  HKD & HJD & HJE  ; 
assign jkc = ~JKC; //complement 
assign jlc =  HKD & hjd & hje  |  hkd & HJD & hje  |  hkd & hjd & HJE  |  hkd & hjd & hje  ; 
assign JLC = ~jlc;  //complement 
assign JMC =  HMD & hld & hlg  |  hmd & HLD & hlg  |  hmd & hld & HLG  |  HMD & HLD & HLG  ; 
assign jmc = ~JMC; //complement 
assign jnc =  HMD & hld & hlg  |  hmd & HLD & hlg  |  hmd & hld & HLG  |  hmd & hld & hlg  ; 
assign JNC = ~jnc;  //complement 
assign JOC =  HOD & hnd & hne  |  hod & HND & hne  |  hod & hnd & HNE  |  HOD & HND & HNE  ; 
assign joc = ~JOC; //complement 
assign jpc =  HOD & hnd & hne  |  hod & HND & hne  |  hod & hnd & HNE  |  hod & hnd & hne  ; 
assign JPC = ~jpc;  //complement 
assign tha = ~THA;  //complement 
assign thc = ~THC;  //complement 
assign the = ~THE;  //complement 
assign aae = ~AAE;  //complement 
assign aaf = ~AAF;  //complement 
assign oae = ~OAE;  //complement 
assign obe = ~OBE;  //complement 
assign hog = ~HOG;  //complement 
assign HPG = ~hpg;  //complement 
assign hqg = ~HQG;  //complement 
assign OHG = ~ohg;  //complement 
assign bde = ~BDE;  //complement 
assign bdf = ~BDF;  //complement 
assign bee = ~BEE;  //complement 
assign bef = ~BEF;  //complement 
assign oaf = ~OAF;  //complement 
assign obf = ~OBF;  //complement 
assign JQB =  HQG & hqb & hpb  |  hqg & HQB & hpb  |  hqg & hqb & HPB  |  HQG & HQB & HPB  ; 
assign jqb = ~JQB; //complement 
assign jrb =  HQG & hqb & hpb  |  hqg & HQB & hpb  |  hqg & hqb & HPB  |  hqg & hqb & hpb  ; 
assign JRB = ~jrb;  //complement 
assign BBE = ~bbe;  //complement 
assign BBF = ~bbf;  //complement 
assign bce = ~BCE;  //complement 
assign bcf = ~BCF;  //complement 
assign ode = ~ODE;  //complement 
assign oee = ~OEE;  //complement 
assign kqc = ~KQC;  //complement 
assign OKC = ~okc;  //complement 
assign okf = ~OKF;  //complement 
assign tta = ~TTA;  //complement 
assign ttc = ~TTC;  //complement 
assign tte = ~TTE;  //complement 
assign bae = ~BAE;  //complement 
assign baf = ~BAF;  //complement 
assign odf = ~ODF;  //complement 
assign oef = ~OEF;  //complement 
assign och = ~OCH;  //complement 
assign TTB = ~ttb;  //complement 
assign TTD = ~ttd;  //complement 
assign TTF = ~ttf;  //complement 
assign bag = ~BAG;  //complement 
assign bah = ~BAH;  //complement 
assign odh = ~ODH;  //complement 
assign oeh = ~OEH;  //complement 
assign ofh = ~OFH;  //complement 
assign JQC =  HQD & hpd & hpe  |  hqd & HPD & hpe  |  hqd & hpd & HPE  |  HQD & HPD & HPE  ; 
assign jqc = ~JQC; //complement 
assign jrc =  HQD & hpd & hpe  |  hqd & HPD & hpe  |  hqd & hpd & HPE  |  hqd & hpd & hpe  ; 
assign JRC = ~jrc;  //complement 
assign omb = ~OMB;  //complement 
assign BBG = ~bbg;  //complement 
assign BBH = ~bbh;  //complement 
assign bcg = ~BCG;  //complement 
assign bch = ~BCH;  //complement 
assign odg = ~ODG;  //complement 
assign oeg = ~OEG;  //complement 
assign ofg = ~OFG;  //complement 
assign okd = ~OKD;  //complement 
assign OLD = ~old;  //complement 
assign bdg = ~BDG;  //complement 
assign bdh = ~BDH;  //complement 
assign beg = ~BEG;  //complement 
assign beh = ~BEH;  //complement 
assign oah = ~OAH;  //complement 
assign obh = ~OBH;  //complement 
assign THB = ~thb;  //complement 
assign THD = ~thd;  //complement 
assign THF = ~thf;  //complement 
assign aag = ~AAG;  //complement 
assign aah = ~AAH;  //complement 
assign oag = ~OAG;  //complement 
assign obg = ~OBG;  //complement 
assign ocg = ~OCG;  //complement 
assign JEA =  HEA & hda & hdc  |  hea & HDA & hdc  |  hea & hda & HDC  |  HEA & HDA & HDC  ; 
assign jea = ~JEA; //complement 
assign jfa =  HEA & hda & hdc  |  hea & HDA & hdc  |  hea & hda & HDC  |  hea & hda & hdc  ; 
assign JFA = ~jfa;  //complement 
assign JGA =  HFA & hga & hfc  |  hfa & HGA & hfc  |  hfa & hga & HFC  |  HFA & HGA & HFC  ; 
assign jga = ~JGA; //complement 
assign jha =  HFA & hga & hfc  |  hfa & HGA & hfc  |  hfa & hga & HFC  |  hfa & hga & hfc  ; 
assign JHA = ~jha;  //complement 
assign JIA =  HIA & hha & hhc  |  hia & HHA & hhc  |  hia & hha & HHC  |  HIA & HHA & HHC  ; 
assign jia = ~JIA; //complement 
assign jja =  HIA & hha & hhc  |  hia & HHA & hhc  |  hia & hha & HHC  |  hia & hha & hhc  ; 
assign JJA = ~jja;  //complement 
assign opq = ~OPQ;  //complement 
assign OQQ = ~oqq;  //complement 
assign opr = ~OPR;  //complement 
assign kea = ~KEA;  //complement 
assign KFA = ~kfa;  //complement 
assign MFA = ~mfa;  //complement 
assign LEA =  KDA & kea & keb  |  kda & KEA & keb  |  kda & kea & KEB  |  KDA & KEA & KEB  ; 
assign lea = ~LEA; //complement 
assign lfa =  KDA & kea & keb  |  kda & KEA & keb  |  kda & kea & KEB  |  kda & kea & keb  ; 
assign LFA = ~lfa;  //complement 
assign JIE =  HIC & hig & hhg  |  hic & HIG & hhg  |  hic & hig & HHG  |  HIC & HIG & HHG  ; 
assign jie = ~JIE; //complement 
assign jje =  HIC & hig & hhg  |  hic & HIG & hhg  |  hic & hig & HHG  |  hic & hig & hhg  ; 
assign JJE = ~jje;  //complement 
assign lda =  KCA & kcb  |  kca & KCB  |  kca & kcb  ; 
assign LDA = ~lda; //complement 
assign mga = ~MGA;  //complement 
assign MHA = ~mha;  //complement 
assign LGA =  KGB & kfb & kgc  |  kgb & KFB & kgc  |  kgb & kfb & KGC  |  KGB & KFB & KGC  ; 
assign lga = ~LGA; //complement 
assign lha =  KGB & kfb & kgc  |  kgb & KFB & kgc  |  kgb & kfb & KGC  |  kgb & kfb & kgc  ; 
assign LHA = ~lha;  //complement 
assign LIB =  KIB & khb & khc  |  kib & KHB & khc  |  kib & khb & KHC  |  KIB & KHB & KHC  ; 
assign lib = ~LIB; //complement 
assign ljb =  KIB & khb & khc  |  kib & KHB & khc  |  kib & khb & KHC  |  kib & khb & khc  ; 
assign LJB = ~ljb;  //complement 
assign JCB =  HBB & hcd & hce  |  hbb & HCD & hce  |  hbb & hcd & HCE  |  HBB & HCD & HCE  ; 
assign jcb = ~JCB; //complement 
assign jdb =  HBB & hcd & hce  |  hbb & HCD & hce  |  hbb & hcd & HCE  |  hbb & hcd & hce  ; 
assign JDB = ~jdb;  //complement 
assign keb = ~KEB;  //complement 
assign KFB = ~kfb;  //complement 
assign kgb = ~KGB;  //complement 
assign KHB = ~khb;  //complement 
assign kib = ~KIB;  //complement 
assign KJB = ~kjb;  //complement 
assign ONB = ~onb;  //complement 
assign JED =  HEE & hde & hef  |  hee & HDE & hef  |  hee & hde & HEF  |  HEE & HDE & HEF  ; 
assign jed = ~JED; //complement 
assign jfd =  HEE & hde & hef  |  hee & HDE & hef  |  hee & hde & HEF  |  hee & hde & hef  ; 
assign JFD = ~jfd;  //complement 
assign JGD =  HGE & hgf & hff  |  hge & HGF & hff  |  hge & hgf & HFF  |  HGE & HGF & HFF  ; 
assign jgd = ~JGD; //complement 
assign jhd =  HGE & hgf & hff  |  hge & HGF & hff  |  hge & hgf & HFF  |  hge & hgf & hff  ; 
assign JHD = ~jhd;  //complement 
assign JID =  HIE & hif & hhf  |  hie & HIF & hhf  |  hie & hif & HHF  |  HIE & HIF & HHF  ; 
assign jid = ~JID; //complement 
assign jjd =  HIE & hif & hhf  |  hie & HIF & hhf  |  hie & hif & HHF  |  hie & hif & hhf  ; 
assign JJD = ~jjd;  //complement 
assign JKA =  HJA & hka & hjc  |  hja & HKA & hjc  |  hja & hka & HJC  |  HJA & HKA & HJC  ; 
assign jka = ~JKA; //complement 
assign jla =  HJA & hka & hjc  |  hja & HKA & hjc  |  hja & hka & HJC  |  hja & hka & hjc  ; 
assign JLA = ~jla;  //complement 
assign JMA =  HMA & hla & hmg  |  hma & HLA & hmg  |  hma & hla & HMG  |  HMA & HLA & HMG  ; 
assign jma = ~JMA; //complement 
assign jna =  HMA & hla & hmg  |  hma & HLA & hmg  |  hma & hla & HMG  |  hma & hla & hmg  ; 
assign JNA = ~jna;  //complement 
assign JOA =  HOA & hna & hng  |  hoa & HNA & hng  |  hoa & hna & HNG  |  HOA & HNA & HNG  ; 
assign joa = ~JOA; //complement 
assign jpa =  HOA & hna & hng  |  hoa & HNA & hng  |  hoa & hna & HNG  |  hoa & hna & hng  ; 
assign JPA = ~jpa;  //complement 
assign LOA =  KNA & koa & koc  |  kna & KOA & koc  |  kna & koa & KOC  |  KNA & KOA & KOC  ; 
assign loa = ~LOA; //complement 
assign lpa =  KNA & koa & koc  |  kna & KOA & koc  |  kna & koa & KOC  |  kna & koa & koc  ; 
assign LPA = ~lpa;  //complement 
assign NQA =  MQA & mqb & mqc  |  mqa & MQB & mqc  |  mqa & mqb & MQC  |  MQA & MQB & MQC  ; 
assign nqa = ~NQA; //complement 
assign nra =  MQA & mqb & mqc  |  mqa & MQB & mqc  |  mqa & mqb & MQC  |  mqa & mqb & mqc  ; 
assign NRA = ~nra;  //complement 
assign mqa = ~MQA;  //complement 
assign OMA = ~oma;  //complement 
assign mqb = ~MQB;  //complement 
assign LKA =  KKC & kke & kjc  |  kkc & KKE & kjc  |  kkc & kke & KJC  |  KKC & KKE & KJC  ; 
assign lka = ~LKA; //complement 
assign lla =  KKC & kke & kjc  |  kkc & KKE & kjc  |  kkc & kke & KJC  |  kkc & kke & kjc  ; 
assign LLA = ~lla;  //complement 
assign mma = ~MMA;  //complement 
assign MNA = ~mna;  //complement 
assign mmb = ~MMB;  //complement 
assign opo = ~OPO;  //complement 
assign OQO = ~oqo;  //complement 
assign LQA =  KPC & kqc & kqa  |  kpc & KQC & kqa  |  kpc & kqc & KQA  |  KPC & KQC & KQA  ; 
assign lqa = ~LQA; //complement 
assign lra =  KPC & kqc & kqa  |  kpc & KQC & kqa  |  kpc & kqc & KQA  |  kpc & kqc & kqa  ; 
assign LRA = ~lra;  //complement 
assign LKB =  KKB & kkd & kjb  |  kkb & KKD & kjb  |  kkb & kkd & KJB  |  KKB & KKD & KJB  ; 
assign lkb = ~LKB; //complement 
assign llb =  KKB & kkd & kjb  |  kkb & KKD & kjb  |  kkb & kkd & KJB  |  kkb & kkd & kjb  ; 
assign LLB = ~llb;  //complement 
assign mkb = ~MKB;  //complement 
assign MLB = ~mlb;  //complement 
assign LMB =  KMB & kmd & klb  |  kmb & KMD & klb  |  kmb & kmd & KLB  |  KMB & KMD & KLB  ; 
assign lmb = ~LMB; //complement 
assign lnb =  KMB & kmd & klb  |  kmb & KMD & klb  |  kmb & kmd & KLB  |  kmb & kmd & klb  ; 
assign LNB = ~lnb;  //complement 
assign LOB =  KOB & kod & knb  |  kob & KOD & knb  |  kob & kod & KNB  |  KOB & KOD & KNB  ; 
assign lob = ~LOB; //complement 
assign lpb =  KOB & kod & knb  |  kob & KOD & knb  |  kob & kod & KNB  |  kob & kod & knb  ; 
assign LPB = ~lpb;  //complement 
assign kkb = ~KKB;  //complement 
assign KLB = ~klb;  //complement 
assign kkd = ~KKD;  //complement 
assign kmb = ~KMB;  //complement 
assign KNB = ~knb;  //complement 
assign kmd = ~KMD;  //complement 
assign kob = ~KOB;  //complement 
assign KPB = ~kpb;  //complement 
assign kod = ~KOD;  //complement 
assign JKD =  HKE & hkh & hkf  |  hke & HKH & hkf  |  hke & hkh & HKF  |  HKE & HKH & HKF  ; 
assign jkd = ~JKD; //complement 
assign jld =  HKE & hkh & hkf  |  hke & HKH & hkf  |  hke & hkh & HKF  |  hke & hkh & hkf  ; 
assign JLD = ~jld;  //complement 
assign JMD =  HME & hmf & hle  |  hme & HMF & hle  |  hme & hmf & HLE  |  HME & HMF & HLE  ; 
assign jmd = ~JMD; //complement 
assign jnd =  HME & hmf & hle  |  hme & HMF & hle  |  hme & hmf & HLE  |  hme & hmf & hle  ; 
assign JND = ~jnd;  //complement 
assign JOD =  HOE & hof & hnf  |  hoe & HOF & hnf  |  hoe & hof & HNF  |  HOE & HOF & HNF  ; 
assign jod = ~JOD; //complement 
assign jpd =  HOE & hof & hnf  |  hoe & HOF & hnf  |  hoe & hof & HNF  |  hoe & hof & hnf  ; 
assign JPD = ~jpd;  //complement 
assign JQA =  HQA & hpa & hpg  |  hqa & HPA & hpg  |  hqa & hpa & HPG  |  HQA & HPA & HPG  ; 
assign jqa = ~JQA; //complement 
assign jra =  HQA & hpa & hpg  |  hqa & HPA & hpg  |  hqa & hpa & HPG  |  hqa & hpa & hpg  ; 
assign JRA = ~jra;  //complement 
assign tsa = ~TSA;  //complement 
assign tsc = ~TSC;  //complement 
assign tse = ~TSE;  //complement 
assign aai = ~AAI;  //complement 
assign aaj = ~AAJ;  //complement 
assign oai = ~OAI;  //complement 
assign obi = ~OBI;  //complement 
assign oci = ~OCI;  //complement 
assign bdi = ~BDI;  //complement 
assign bdj = ~BDJ;  //complement 
assign bei = ~BEI;  //complement 
assign bej = ~BEJ;  //complement 
assign oaj = ~OAJ;  //complement 
assign obj = ~OBJ;  //complement 
assign ocj = ~OCJ;  //complement 
assign kqa = ~KQA;  //complement 
assign OKA = ~oka;  //complement 
assign oke = ~OKE;  //complement 
assign BBI = ~bbi;  //complement 
assign BBJ = ~bbj;  //complement 
assign bci = ~BCI;  //complement 
assign bcj = ~BCJ;  //complement 
assign odi = ~ODI;  //complement 
assign oei = ~OEI;  //complement 
assign ofi = ~OFI;  //complement 
assign bck = ~BCK;  //complement 
assign tga = ~TGA;  //complement 
assign tgc = ~TGC;  //complement 
assign tge = ~TGE;  //complement 
assign bai = ~BAI;  //complement 
assign baj = ~BAJ;  //complement 
assign odj = ~ODJ;  //complement 
assign oej = ~OEJ;  //complement 
assign ofj = ~OFJ;  //complement 
assign obl = ~OBL;  //complement 
assign TGB = ~tgb;  //complement 
assign TGD = ~tgd;  //complement 
assign TGF = ~tgf;  //complement 
assign bak = ~BAK;  //complement 
assign bal = ~BAL;  //complement 
assign odl = ~ODL;  //complement 
assign oel = ~OEL;  //complement 
assign ofl = ~OFL;  //complement 
assign kqb = ~KQB;  //complement 
assign OKB = ~okb;  //complement 
assign kqd = ~KQD;  //complement 
assign LQB =  KQB & kqd & kpb  |  kqb & KQD & kpb  |  kqb & kqd & KPB  |  KQB & KQD & KPB  ; 
assign lqb = ~LQB; //complement 
assign lrb =  KQB & kqd & kpb  |  kqb & KQD & kpb  |  kqb & kqd & KPB  |  kqb & kqd & kpb  ; 
assign LRB = ~lrb;  //complement 
assign BBK = ~bbk;  //complement 
assign BBL = ~bbl;  //complement 
assign bcl = ~BCL;  //complement 
assign odk = ~ODK;  //complement 
assign oek = ~OEK;  //complement 
assign ofk = ~OFK;  //complement 
assign JQD =  HQE & hqi & hqf  |  hqe & HQI & hqf  |  hqe & hqi & HQF  |  HQE & HQI & HQF  ; 
assign jqd = ~JQD; //complement 
assign jrd =  HQE & hqi & hqf  |  hqe & HQI & hqf  |  hqe & hqi & HQF  |  hqe & hqi & hqf  ; 
assign JRD = ~jrd;  //complement 
assign JQE =  HQC & hqh & hpc  |  hqc & HQH & hpc  |  hqc & hqh & HPC  |  HQC & HQH & HPC  ; 
assign jqe = ~JQE; //complement 
assign jre =  HQC & hqh & hpc  |  hqc & HQH & hpc  |  hqc & hqh & HPC  |  hqc & hqh & hpc  ; 
assign JRE = ~jre;  //complement 
assign bdk = ~BDK;  //complement 
assign bdl = ~BDL;  //complement 
assign bek = ~BEK;  //complement 
assign bel = ~BEL;  //complement 
assign oal = ~OAL;  //complement 
assign ocl = ~OCL;  //complement 
assign TSB = ~tsb;  //complement 
assign TSD = ~tsd;  //complement 
assign TSF = ~tsf;  //complement 
assign aak = ~AAK;  //complement 
assign aal = ~AAL;  //complement 
assign oak = ~OAK;  //complement 
assign obk = ~OBK;  //complement 
assign ock = ~OCK;  //complement 
assign hca = ~HCA;  //complement 
assign HDA = ~hda;  //complement 
assign hea = ~HEA;  //complement 
assign HFA = ~hfa;  //complement 
assign hga = ~HGA;  //complement 
assign HHA = ~hha;  //complement 
assign hia = ~HIA;  //complement 
assign HJA = ~hja;  //complement 
assign GAA =  FAA & fab & faf  |  faa & FAB & faf  |  faa & fab & FAF  |  FAA & FAB & FAF  ; 
assign gaa = ~GAA; //complement 
assign gba =  FAA & fab & faf  |  faa & FAB & faf  |  faa & fab & FAF  |  faa & fab & faf  ; 
assign GBA = ~gba;  //complement 
assign GCA =  FCB & fcc & fcg  |  fcb & FCC & fcg  |  fcb & fcc & FCG  |  FCB & FCC & FCG  ; 
assign gca = ~GCA; //complement 
assign gda =  FCB & fcc & fcg  |  fcb & FCC & fcg  |  fcb & fcc & FCG  |  fcb & fcc & fcg  ; 
assign GDA = ~gda;  //complement 
assign GEB =  FEH & fec & fed  |  feh & FEC & fed  |  feh & fec & FED  |  FEH & FEC & FED  ; 
assign geb = ~GEB; //complement 
assign gfb =  FEH & fec & fed  |  feh & FEC & fed  |  feh & fec & FED  |  feh & fec & fed  ; 
assign GFB = ~gfb;  //complement 
assign GGA =  FGG & fgc & fgb  |  fgg & FGC & fgb  |  fgg & fgc & FGB  |  FGG & FGC & FGB  ; 
assign gga = ~GGA; //complement 
assign gha =  FGG & fgc & fgb  |  fgg & FGC & fgb  |  fgg & fgc & FGB  |  fgg & fgc & fgb  ; 
assign GHA = ~gha;  //complement 
assign GCF =  FBE & fba & fbb  |  fbe & FBA & fbb  |  fbe & fba & FBB  |  FBE & FBA & FBB  ; 
assign gcf = ~GCF; //complement 
assign gdf =  FBE & fba & fbb  |  fbe & FBA & fbb  |  fbe & fba & FBB  |  fbe & fba & fbb  ; 
assign GDF = ~gdf;  //complement 
assign GGF =  FFC & ffg & ffd  |  ffc & FFG & ffd  |  ffc & ffg & FFD  |  FFC & FFG & FFD  ; 
assign ggf = ~GGF; //complement 
assign ghf =  FFC & ffg & ffd  |  ffc & FFG & ffd  |  ffc & ffg & FFD  |  ffc & ffg & ffd  ; 
assign GHF = ~ghf;  //complement 
assign GIG =  FHB & fhc & fhf  |  fhb & FHC & fhf  |  fhb & fhc & FHF  |  FHB & FHC & FHF  ; 
assign gig = ~GIG; //complement 
assign gjg =  FHB & fhc & fhf  |  fhb & FHC & fhf  |  fhb & fhc & FHF  |  fhb & fhc & fhf  ; 
assign GJG = ~gjg;  //complement 
assign GGE =  FFF & ffe & fge  |  fff & FFE & fge  |  fff & ffe & FGE  |  FFF & FFE & FGE  ; 
assign gge = ~GGE; //complement 
assign ghe =  FFF & ffe & fge  |  fff & FFE & fge  |  fff & ffe & FGE  |  fff & ffe & fge  ; 
assign GHE = ~ghe;  //complement 
assign hec = ~HEC;  //complement 
assign HFC = ~hfc;  //complement 
assign hgc = ~HGC;  //complement 
assign HHC = ~hhc;  //complement 
assign hic = ~HIC;  //complement 
assign HJC = ~hjc;  //complement 
assign hig = ~HIG;  //complement 
assign hcd = ~HCD;  //complement 
assign HDD = ~hdd;  //complement 
assign heg = ~HEG;  //complement 
assign GEA =  FEA & feb & feg  |  fea & FEB & feg  |  fea & feb & FEG  |  FEA & FEB & FEG  ; 
assign gea = ~GEA; //complement 
assign gfa =  FEA & feb & feg  |  fea & FEB & feg  |  fea & feb & FEG  |  fea & feb & feg  ; 
assign GFA = ~gfa;  //complement 
assign hgg = ~HGG;  //complement 
assign HHG = ~hhg;  //complement 
assign GCE =  FCE & fbd & fbc  |  fce & FBD & fbc  |  fce & fbd & FBC  |  FCE & FBD & FBC  ; 
assign gce = ~GCE; //complement 
assign gde =  FCE & fbd & fbc  |  fce & FBD & fbc  |  fce & fbd & FBC  |  fce & fbd & fbc  ; 
assign GDE = ~gde;  //complement 
assign GEF =  FEF & fde & fdd  |  fef & FDE & fdd  |  fef & fde & FDD  |  FEF & FDE & FDD  ; 
assign gef = ~GEF; //complement 
assign gff =  FEF & fde & fdd  |  fef & FDE & fdd  |  fef & fde & FDD  |  fef & fde & fdd  ; 
assign GFF = ~gff;  //complement 
assign haa = ~HAA;  //complement 
assign HBA = ~hba;  //complement 
assign GIF =  FHA & fhe & fhd  |  fha & FHE & fhd  |  fha & fhe & FHD  |  FHA & FHE & FHD  ; 
assign gif = ~GIF; //complement 
assign gjf =  FHA & fhe & fhd  |  fha & FHE & fhd  |  fha & fhe & FHD  |  fha & fhe & fhd  ; 
assign GJF = ~gjf;  //complement 
assign hce = ~HCE;  //complement 
assign HDE = ~hde;  //complement 
assign hee = ~HEE;  //complement 
assign HFE = ~hfe;  //complement 
assign GEG =  FDF & fdb & fdc  |  fdf & FDB & fdc  |  fdf & fdb & FDC  |  FDF & FDB & FDC  ; 
assign geg = ~GEG; //complement 
assign gfg =  FDF & fdb & fdc  |  fdf & FDB & fdc  |  fdf & fdb & FDC  |  fdf & fdb & fdc  ; 
assign GFG = ~gfg;  //complement 
assign hie = ~HIE;  //complement 
assign HJE = ~hje;  //complement 
assign hge = ~HGE;  //complement 
assign HHE = ~hhe;  //complement 
assign hef = ~HEF;  //complement 
assign HFF = ~hff;  //complement 
assign hgf = ~HGF;  //complement 
assign HHF = ~hhf;  //complement 
assign hif = ~HIF;  //complement 
assign HJF = ~hjf;  //complement 
assign hka = ~HKA;  //complement 
assign HLA = ~hla;  //complement 
assign hma = ~HMA;  //complement 
assign HNA = ~hna;  //complement 
assign hoa = ~HOA;  //complement 
assign HPA = ~hpa;  //complement 
assign GIB =  FIH & fic & fid  |  fih & FIC & fid  |  fih & fic & FID  |  FIH & FIC & FID  ; 
assign gib = ~GIB; //complement 
assign gjb =  FIH & fic & fid  |  fih & FIC & fid  |  fih & fic & FID  |  fih & fic & fid  ; 
assign GJB = ~gjb;  //complement 
assign GKB =  FKI & fkd & fke  |  fki & FKD & fke  |  fki & fkd & FKE  |  FKI & FKD & FKE  ; 
assign gkb = ~GKB; //complement 
assign glb =  FKI & fkd & fke  |  fki & FKD & fke  |  fki & fkd & FKE  |  fki & fkd & fke  ; 
assign GLB = ~glb;  //complement 
assign GMB =  FMH & fmc & fmd  |  fmh & FMC & fmd  |  fmh & fmc & FMD  |  FMH & FMC & FMD  ; 
assign gmb = ~GMB; //complement 
assign gnb =  FMH & fmc & fmd  |  fmh & FMC & fmd  |  fmh & fmc & FMD  |  fmh & fmc & fmd  ; 
assign GNB = ~gnb;  //complement 
assign GKG =  FJC & fjd & fjg  |  fjc & FJD & fjg  |  fjc & fjd & FJG  |  FJC & FJD & FJG  ; 
assign gkg = ~GKG; //complement 
assign glg =  FJC & fjd & fjg  |  fjc & FJD & fjg  |  fjc & fjd & FJG  |  fjc & fjd & fjg  ; 
assign GLG = ~glg;  //complement 
assign GMG =  FLH & fld & fle  |  flh & FLD & fle  |  flh & fld & FLE  |  FLH & FLD & FLE  ; 
assign gmg = ~GMG; //complement 
assign gng =  FLH & fld & fle  |  flh & FLD & fle  |  flh & fld & FLE  |  flh & fld & fle  ; 
assign GNG = ~gng;  //complement 
assign GOH =  FNC & fnd & fng  |  fnc & FND & fng  |  fnc & fnd & FNG  |  FNC & FND & FNG  ; 
assign goh = ~GOH; //complement 
assign gph =  FNC & fnd & fng  |  fnc & FND & fng  |  fnc & fnd & FNG  |  fnc & fnd & fng  ; 
assign GPH = ~gph;  //complement 
assign hkc = ~HKC;  //complement 
assign HLC = ~hlc;  //complement 
assign hmc = ~HMC;  //complement 
assign HNC = ~hnc;  //complement 
assign hoc = ~HOC;  //complement 
assign HPC = ~hpc;  //complement 
assign GIA =  FIF & fig & fib  |  fif & FIG & fib  |  fif & fig & FIB  |  FIF & FIG & FIB  ; 
assign gia = ~GIA; //complement 
assign gja =  FIF & fig & fib  |  fif & FIG & fib  |  fif & fig & FIB  |  fif & fig & fib  ; 
assign GJA = ~gja;  //complement 
assign hoe = ~HOE;  //complement 
assign HPE = ~hpe;  //complement 
assign GKA =  FKG & fkh & fkc  |  fkg & FKH & fkc  |  fkg & fkh & FKC  |  FKG & FKH & FKC  ; 
assign gka = ~GKA; //complement 
assign gla =  FKG & fkh & fkc  |  fkg & FKH & fkc  |  fkg & fkh & FKC  |  fkg & fkh & fkc  ; 
assign GLA = ~gla;  //complement 
assign GMA =  FMF & fmg & fmb  |  fmf & FMG & fmb  |  fmf & fmg & FMB  |  FMF & FMG & FMB  ; 
assign gma = ~GMA; //complement 
assign gna =  FMF & fmg & fmb  |  fmf & FMG & fmb  |  fmf & fmg & FMB  |  fmf & fmg & fmb  ; 
assign GNA = ~gna;  //complement 
assign GKF =  FJB & fje & fjf  |  fjb & FJE & fjf  |  fjb & fje & FJF  |  FJB & FJE & FJF  ; 
assign gkf = ~GKF; //complement 
assign glf =  FJB & fje & fjf  |  fjb & FJE & fjf  |  fjb & fje & FJF  |  fjb & fje & fjf  ; 
assign GLF = ~glf;  //complement 
assign GMF =  FLF & flg & flc  |  flf & FLG & flc  |  flf & flg & FLC  |  FLF & FLG & FLC  ; 
assign gmf = ~GMF; //complement 
assign gnf =  FLF & flg & flc  |  flf & FLG & flc  |  flf & flg & FLC  |  flf & flg & flc  ; 
assign GNF = ~gnf;  //complement 
assign GOG =  FNE & fnf & fnb  |  fne & FNF & fnb  |  fne & fnf & FNB  |  FNE & FNF & FNB  ; 
assign gog = ~GOG; //complement 
assign gpg =  FNE & fnf & fnb  |  fne & FNF & fnb  |  fne & fnf & FNB  |  fne & fnf & fnb  ; 
assign GPG = ~gpg;  //complement 
assign hke = ~HKE;  //complement 
assign HLE = ~hle;  //complement 
assign hkh = ~HKH;  //complement 
assign hme = ~HME;  //complement 
assign HNE = ~hne;  //complement 
assign hkf = ~HKF;  //complement 
assign HLF = ~hlf;  //complement 
assign hmf = ~HMF;  //complement 
assign HNF = ~hnf;  //complement 
assign hof = ~HOF;  //complement 
assign HPF = ~hpf;  //complement 
assign hqa = ~HQA;  //complement 
assign OHA = ~oha;  //complement 
assign tka = ~TKA;  //complement 
assign tke = ~TKE;  //complement 
assign aam = ~AAM;  //complement 
assign aan = ~AAN;  //complement 
assign oam = ~OAM;  //complement 
assign obm = ~OBM;  //complement 
assign ocm = ~OCM;  //complement 
assign GOC =  FOD & foe & foi  |  fod & FOE & foi  |  fod & foe & FOI  |  FOD & FOE & FOI  ; 
assign goc = ~GOC; //complement 
assign gpc =  FOD & foe & foi  |  fod & FOE & foi  |  fod & foe & FOI  |  fod & foe & foi  ; 
assign GPC = ~gpc;  //complement 
assign GQB =  FQC & fqd & fqh  |  fqc & FQD & fqh  |  fqc & fqd & FQH  |  FQC & FQD & FQH  ; 
assign gqb = ~GQB; //complement 
assign grb =  FQC & fqd & fqh  |  fqc & FQD & fqh  |  fqc & fqd & FQH  |  fqc & fqd & fqh  ; 
assign GRB = ~grb;  //complement 
assign bdm = ~BDM;  //complement 
assign bdn = ~BDN;  //complement 
assign bem = ~BEM;  //complement 
assign ben = ~BEN;  //complement 
assign oan = ~OAN;  //complement 
assign obn = ~OBN;  //complement 
assign ocn = ~OCN;  //complement 
assign GQG =  FPD & fpe & fph  |  fpd & FPE & fph  |  fpd & fpe & FPH  |  FPD & FPE & FPH  ; 
assign gqg = ~GQG; //complement 
assign grg =  FPD & fpe & fph  |  fpd & FPE & fph  |  fpd & fpe & FPH  |  fpd & fpe & fph  ; 
assign GRG = ~grg;  //complement 
assign ocp = ~OCP;  //complement 
assign BBM = ~bbm;  //complement 
assign BBN = ~bbn;  //complement 
assign bcm = ~BCM;  //complement 
assign bcn = ~BCN;  //complement 
assign odm = ~ODM;  //complement 
assign oem = ~OEM;  //complement 
assign ofm = ~OFM;  //complement 
assign bco = ~BCO;  //complement 
assign BBP = ~bbp;  //complement 
assign hqc = ~HQC;  //complement 
assign OHC = ~ohc;  //complement 
assign hqh = ~HQH;  //complement 
assign bam = ~BAM;  //complement 
assign ban = ~BAN;  //complement 
assign odn = ~ODN;  //complement 
assign oen = ~OEN;  //complement 
assign ofn = ~OFN;  //complement 
assign GOB =  FOG & foh & foc  |  fog & FOH & foc  |  fog & foh & FOC  |  FOG & FOH & FOC  ; 
assign gob = ~GOB; //complement 
assign gpb =  FOG & foh & foc  |  fog & FOH & foc  |  fog & foh & FOC  |  fog & foh & foc  ; 
assign GPB = ~gpb;  //complement 
assign GQA =  FQB & fqg & fqf  |  fqb & FQG & fqf  |  fqb & fqg & FQF  |  FQB & FQG & FQF  ; 
assign gqa = ~GQA; //complement 
assign gra =  FQB & fqg & fqf  |  fqb & FQG & fqf  |  fqb & fqg & FQF  |  fqb & fqg & fqf  ; 
assign GRA = ~gra;  //complement 
assign bao = ~BAO;  //complement 
assign bap = ~BAP;  //complement 
assign odp = ~ODP;  //complement 
assign oep = ~OEP;  //complement 
assign ofp = ~OFP;  //complement 
assign GQF =  FPF & fpg & fpc  |  fpf & FPG & fpc  |  fpf & fpg & FPC  |  FPF & FPG & FPC  ; 
assign gqf = ~GQF; //complement 
assign grf =  FPF & fpg & fpc  |  fpf & FPG & fpc  |  fpf & fpg & FPC  |  fpf & fpg & fpc  ; 
assign GRF = ~grf;  //complement 
assign BBO = ~bbo;  //complement 
assign bcp = ~BCP;  //complement 
assign odo = ~ODO;  //complement 
assign oeo = ~OEO;  //complement 
assign ofo = ~OFO;  //complement 
assign hqe = ~HQE;  //complement 
assign OHE = ~ohe;  //complement 
assign hqi = ~HQI;  //complement 
assign GOA =  FNA & foa & fob  |  fna & FOA & fob  |  fna & foa & FOB  |  FNA & FOA & FOB  ; 
assign goa = ~GOA; //complement 
assign gpa =  FNA & foa & fob  |  fna & FOA & fob  |  fna & foa & FOB  |  fna & foa & fob  ; 
assign GPA = ~gpa;  //complement 
assign bdo = ~BDO;  //complement 
assign bdp = ~BDP;  //complement 
assign beo = ~BEO;  //complement 
assign bep = ~BEP;  //complement 
assign oap = ~OAP;  //complement 
assign obp = ~OBP;  //complement 
assign hqf = ~HQF;  //complement 
assign OHF = ~ohf;  //complement 
assign TKB = ~tkb;  //complement 
assign tkc = ~TKC;  //complement 
assign TKD = ~tkd;  //complement 
assign TKF = ~tkf;  //complement 
assign aao = ~AAO;  //complement 
assign aap = ~AAP;  //complement 
assign oao = ~OAO;  //complement 
assign obo = ~OBO;  //complement 
assign oco = ~OCO;  //complement 
assign EAO =  DAO & CEK  ; 
assign eao = ~EAO;  //complement 
assign EAQ =  DBA & CEI  ; 
assign eaq = ~EAQ;  //complement 
assign EAP =  DAP & CEJ  ; 
assign eap = ~EAP;  //complement 
assign ECP =  DAP & CEK  ; 
assign ecp = ~ECP;  //complement 
assign ECQ =  DBA & CEJ  ; 
assign ecq = ~ECQ;  //complement 
assign ECR =  DBB & CEI  ; 
assign ecr = ~ECR;  //complement 
assign EEQ =  DBA & CEK  ; 
assign eeq = ~EEQ;  //complement 
assign EER =  DBB & CEJ  ; 
assign eer = ~EER;  //complement 
assign EES =  DBC & CEI  ; 
assign ees = ~EES;  //complement 
assign EGR =  DBB & CEK  ; 
assign egr = ~EGR;  //complement 
assign EGS =  DBC & CEJ  ; 
assign egs = ~EGS;  //complement 
assign EGT =  DBD & CEI  ; 
assign egt = ~EGT;  //complement 
assign faf = ~FAF;  //complement 
assign FBF = ~fbf;  //complement 
assign fcg = ~FCG;  //complement 
assign FDG = ~fdg;  //complement 
assign fca = ~FCA;  //complement 
assign feh = ~FEH;  //complement 
assign FFH = ~ffh;  //complement 
assign fgg = ~FGG;  //complement 
assign FHG = ~fhg;  //complement 
assign EAL =  DAL & CEN  ; 
assign eal = ~EAL;  //complement 
assign EAN =  DAN & CEL  ; 
assign ean = ~EAN;  //complement 
assign ECN =  DAN & CEM  ; 
assign ecn = ~ECN;  //complement 
assign EGN =  DAN & CEO  ; 
assign egn = ~EGN;  //complement 
assign EEN =  DAN & CEN  ; 
assign een = ~EEN;  //complement 
assign EEO =  DAO & CEM  ; 
assign eeo = ~EEO;  //complement 
assign EEP =  DAP & CEL  ; 
assign eep = ~EEP;  //complement 
assign EGO =  DAO & CEN  ; 
assign ego = ~EGO;  //complement 
assign EGP =  DAP & CEM  ; 
assign egp = ~EGP;  //complement 
assign EGQ =  DBA & CEL  ; 
assign egq = ~EGQ;  //complement 
assign fae = ~FAE;  //complement 
assign FBE = ~fbe;  //complement 
assign fcf = ~FCF;  //complement 
assign FDF = ~fdf;  //complement 
assign feb = ~FEB;  //complement 
assign feg = ~FEG;  //complement 
assign FFG = ~ffg;  //complement 
assign fgf = ~FGF;  //complement 
assign FHF = ~fhf;  //complement 
assign EAI =  DAI & CFA  ; 
assign eai = ~EAI;  //complement 
assign EAJ =  DAJ & CEP  ; 
assign eaj = ~EAJ;  //complement 
assign EAK =  DAK & CEO  ; 
assign eak = ~EAK;  //complement 
assign ECJ =  DAJ & CFA  ; 
assign ecj = ~ECJ;  //complement 
assign ECK =  DAK & CEP  ; 
assign eck = ~ECK;  //complement 
assign ECL =  DAL & CEO  ; 
assign ecl = ~ECL;  //complement 
assign EEK =  DAK & CFA  ; 
assign eek = ~EEK;  //complement 
assign EEL =  DAL & CEP  ; 
assign eel = ~EEL;  //complement 
assign EEM =  DAM & CEO  ; 
assign eem = ~EEM;  //complement 
assign EAM =  DAM & CEM  ; 
assign eam = ~EAM;  //complement 
assign EGL =  DAL & CFA  ; 
assign egl = ~EGL;  //complement 
assign EGM =  DAM & CEP  ; 
assign egm = ~EGM;  //complement 
assign fad = ~FAD;  //complement 
assign FBD = ~fbd;  //complement 
assign fce = ~FCE;  //complement 
assign FDE = ~fde;  //complement 
assign fef = ~FEF;  //complement 
assign FFF = ~fff;  //complement 
assign fge = ~FGE;  //complement 
assign FHE = ~fhe;  //complement 
assign EAF =  DAF & CFD  ; 
assign eaf = ~EAF;  //complement 
assign EAG =  DAG & CFC  ; 
assign eag = ~EAG;  //complement 
assign EAH =  DAH & CFB  ; 
assign eah = ~EAH;  //complement 
assign ECG =  DAG & CFD  ; 
assign ecg = ~ECG;  //complement 
assign ECH =  DAH & CFC  ; 
assign ech = ~ECH;  //complement 
assign ECI =  DAI & CFB  ; 
assign eci = ~ECI;  //complement 
assign EEH =  DAH & CFD  ; 
assign eeh = ~EEH;  //complement 
assign EEJ =  DAJ & CFB  ; 
assign eej = ~EEJ;  //complement 
assign EGI =  DAI & CFD  ; 
assign egi = ~EGI;  //complement 
assign EGJ =  DAJ & CFC  ; 
assign egj = ~EGJ;  //complement 
assign EGK =  DAK & CFB  ; 
assign egk = ~EGK;  //complement 
assign fac = ~FAC;  //complement 
assign FBC = ~fbc;  //complement 
assign fcd = ~FCD;  //complement 
assign FDD = ~fdd;  //complement 
assign fee = ~FEE;  //complement 
assign FFE = ~ffe;  //complement 
assign fgd = ~FGD;  //complement 
assign FHD = ~fhd;  //complement 
assign EIS =  DBC & CEK  ; 
assign eis = ~EIS;  //complement 
assign EIT =  DBD & CEJ  ; 
assign eit = ~EIT;  //complement 
assign EIU =  DBE & CEI  ; 
assign eiu = ~EIU;  //complement 
assign oaa = ~OAA;  //complement 
assign cei = ~CEI;  //complement 
assign cej = ~CEJ;  //complement 
assign cek = ~CEK;  //complement 
assign EKS =  DHC & CBL  ; 
assign eks = ~EKS;  //complement 
assign EKT =  DHD & CBK  ; 
assign ekt = ~EKT;  //complement 
assign EKU =  DHE & CBJ  ; 
assign eku = ~EKU;  //complement 
assign fih = ~FIH;  //complement 
assign FJH = ~fjh;  //complement 
assign aaa = ~AAA;  //complement 
assign DBB = ~dbb;  //complement 
assign DBC = ~dbc;  //complement 
assign DBD = ~dbd;  //complement 
assign DBE = ~dbe;  //complement 
assign fki = ~FKI;  //complement 
assign FLI = ~fli;  //complement 
assign EIP =  DAP & CEN  ; 
assign eip = ~EIP;  //complement 
assign EIQ =  DBA & CEM  ; 
assign eiq = ~EIQ;  //complement 
assign EIR =  DBB & CEL  ; 
assign eir = ~EIR;  //complement 
assign daf = ~DAF;  //complement 
assign dag = ~DAG;  //complement 
assign cel = ~CEL;  //complement 
assign cem = ~CEM;  //complement 
assign cen = ~CEN;  //complement 
assign EKQ =  DHA & CBN  ; 
assign ekq = ~EKQ;  //complement 
assign EKR =  DHB & CBM  ; 
assign ekr = ~EKR;  //complement 
assign EKV =  DBF & CBI  ; 
assign ekv = ~EKV;  //complement 
assign fig = ~FIG;  //complement 
assign FJG = ~fjg;  //complement 
assign dan = ~DAN;  //complement 
assign dao = ~DAO;  //complement 
assign dap = ~DAP;  //complement 
assign dba = ~DBA;  //complement 
assign fkh = ~FKH;  //complement 
assign FLH = ~flh;  //complement 
assign EIM =  DAM & CFA  ; 
assign eim = ~EIM;  //complement 
assign EIN =  DAN & CEP  ; 
assign ein = ~EIN;  //complement 
assign EIO =  DAO & CEO  ; 
assign eio = ~EIO;  //complement 
assign ceo = ~CEO;  //complement 
assign cep = ~CEP;  //complement 
assign cfa = ~CFA;  //complement 
assign EKN =  DGN & CCA  ; 
assign ekn = ~EKN;  //complement 
assign EKO =  DGO & CBP  ; 
assign eko = ~EKO;  //complement 
assign EKP =  DGP & CBO  ; 
assign ekp = ~EKP;  //complement 
assign fif = ~FIF;  //complement 
assign FJF = ~fjf;  //complement 
assign dam = ~DAM;  //complement 
assign daj = ~DAJ;  //complement 
assign dal = ~DAL;  //complement 
assign dak = ~DAK;  //complement 
assign fkg = ~FKG;  //complement 
assign FLG = ~flg;  //complement 
assign TRC = ~trc;  //complement 
assign EIJ =  DAJ & CFD  ; 
assign eij = ~EIJ;  //complement 
assign EIK =  DAK & CFC  ; 
assign eik = ~EIK;  //complement 
assign EIL =  DAL & CFB  ; 
assign eil = ~EIL;  //complement 
assign ECM =  DAM & CEN  ; 
assign ecm = ~ECM;  //complement 
assign ECO =  DAO & CEL  ; 
assign eco = ~ECO;  //complement 
assign EEI =  DAI & CFC  ; 
assign eei = ~EEI;  //complement 
assign cfb = ~CFB;  //complement 
assign cfc = ~CFC;  //complement 
assign cfd = ~CFD;  //complement 
assign EKK =  DGK & CCD  ; 
assign ekk = ~EKK;  //complement 
assign EKL =  DGL & CCC  ; 
assign ekl = ~EKL;  //complement 
assign EKM =  DGM & CCB  ; 
assign ekm = ~EKM;  //complement 
assign fie = ~FIE;  //complement 
assign FJE = ~fje;  //complement 
assign fqf = ~FQF;  //complement 
assign OGF = ~ogf;  //complement 
assign dah = ~DAH;  //complement 
assign dai = ~DAI;  //complement 
assign fkf = ~FKF;  //complement 
assign FLF = ~flf;  //complement 
assign EMU =  DHE & CBK  ; 
assign emu = ~EMU;  //complement 
assign EMV =  DBF & CBJ  ; 
assign emv = ~EMV;  //complement 
assign EMW =  DBG & CBI  ; 
assign emw = ~EMW;  //complement 
assign EOV =  DBF & CBK  ; 
assign eov = ~EOV;  //complement 
assign EOW =  DBG & CBJ  ; 
assign eow = ~EOW;  //complement 
assign EOX =  DBH & CBI  ; 
assign eox = ~EOX;  //complement 
assign EQW =  DBG & CBK  ; 
assign eqw = ~EQW;  //complement 
assign EQX =  DBH & CBJ  ; 
assign eqx = ~EQX;  //complement 
assign ERA =  DBI & CBI  ; 
assign era = ~ERA;  //complement 
assign cbi = ~CBI;  //complement 
assign cbj = ~CBJ;  //complement 
assign cbk = ~CBK;  //complement 
assign fmh = ~FMH;  //complement 
assign FNH = ~fnh;  //complement 
assign foi = ~FOI;  //complement 
assign FPI = ~fpi;  //complement 
assign fqh = ~FQH;  //complement 
assign OGH = ~ogh;  //complement 
assign DBF = ~dbf;  //complement 
assign DBG = ~dbg;  //complement 
assign DBH = ~dbh;  //complement 
assign DBI = ~dbi;  //complement 
assign EMR =  DHB & CBN  ; 
assign emr = ~EMR;  //complement 
assign EMS =  DHC & CBM  ; 
assign ems = ~EMS;  //complement 
assign EMT =  DHD & CBL  ; 
assign emt = ~EMT;  //complement 
assign EOS =  DHC & CBN  ; 
assign eos = ~EOS;  //complement 
assign EOT =  DHD & CBM  ; 
assign eot = ~EOT;  //complement 
assign EOU =  DHE & CBL  ; 
assign eou = ~EOU;  //complement 
assign EQT =  DHD & CBN  ; 
assign eqt = ~EQT;  //complement 
assign EQU =  DHE & CBM  ; 
assign equ = ~EQU;  //complement 
assign EQV =  DBF & CBL  ; 
assign eqv = ~EQV;  //complement 
assign cbl = ~CBL;  //complement 
assign cbm = ~CBM;  //complement 
assign cbn = ~CBN;  //complement 
assign fmg = ~FMG;  //complement 
assign FNG = ~fng;  //complement 
assign foh = ~FOH;  //complement 
assign FPH = ~fph;  //complement 
assign fqg = ~FQG;  //complement 
assign OGG = ~ogg;  //complement 
assign DHB = ~dhb;  //complement 
assign DHC = ~dhc;  //complement 
assign DHD = ~dhd;  //complement 
assign DHE = ~dhe;  //complement 
assign EMO =  DGO & CCA  ; 
assign emo = ~EMO;  //complement 
assign EMP =  DGP & CBP  ; 
assign emp = ~EMP;  //complement 
assign EMQ =  DHA & CBO  ; 
assign emq = ~EMQ;  //complement 
assign EOP =  DGP & CCA  ; 
assign eop = ~EOP;  //complement 
assign EOQ =  DHA & CBP  ; 
assign eoq = ~EOQ;  //complement 
assign EOR =  DHB & CBO  ; 
assign eor = ~EOR;  //complement 
assign EQQ =  DHA & CCA  ; 
assign eqq = ~EQQ;  //complement 
assign EQR =  DHB & CBP  ; 
assign eqr = ~EQR;  //complement 
assign EQS =  DHC & CBO  ; 
assign eqs = ~EQS;  //complement 
assign cbo = ~CBO;  //complement 
assign cbp = ~CBP;  //complement 
assign cca = ~CCA;  //complement 
assign fmf = ~FMF;  //complement 
assign FNF = ~fnf;  //complement 
assign fog = ~FOG;  //complement 
assign FPG = ~fpg;  //complement 
assign trb = ~TRB;  //complement 
assign dgn = ~DGN;  //complement 
assign dgo = ~DGO;  //complement 
assign dgp = ~DGP;  //complement 
assign dha = ~DHA;  //complement 
assign EML =  DGL & CCD  ; 
assign eml = ~EML;  //complement 
assign EMN =  DGN & CCB  ; 
assign emn = ~EMN;  //complement 
assign EMM =  DGM & CCC  ; 
assign emm = ~EMM;  //complement 
assign EOM =  DGM & CCD  ; 
assign eom = ~EOM;  //complement 
assign EON =  DGN & CCC  ; 
assign eon = ~EON;  //complement 
assign EOO =  DGO & CCB  ; 
assign eoo = ~EOO;  //complement 
assign EQN =  DGN & CCD  ; 
assign eqn = ~EQN;  //complement 
assign EQO =  DGO & CCC  ; 
assign eqo = ~EQO;  //complement 
assign EQP =  DGP & CCB  ; 
assign eqp = ~EQP;  //complement 
assign ccb = ~CCB;  //complement 
assign ccc = ~CCC;  //complement 
assign ccd = ~CCD;  //complement 
assign fme = ~FME;  //complement 
assign FNE = ~fne;  //complement 
assign fof = ~FOF;  //complement 
assign FPF = ~fpf;  //complement 
assign fqe = ~FQE;  //complement 
assign OGE = ~oge;  //complement 
assign dgk = ~DGK;  //complement 
assign dgl = ~DGL;  //complement 
assign dgm = ~DGM;  //complement 
assign fab = ~FAB;  //complement 
assign FBB = ~fbb;  //complement 
assign fcc = ~FCC;  //complement 
assign FDC = ~fdc;  //complement 
assign fed = ~FED;  //complement 
assign FFD = ~ffd;  //complement 
assign fgc = ~FGC;  //complement 
assign FHC = ~fhc;  //complement 
assign EAC =  DDC & CFG  ; 
assign eac = ~EAC;  //complement 
assign EAD =  DDD & CFF  ; 
assign ead = ~EAD;  //complement 
assign EAE =  DDE & CFE  ; 
assign eae = ~EAE;  //complement 
assign ECD =  DDD & CFG  ; 
assign ecd = ~ECD;  //complement 
assign ECE =  DDE & CFF  ; 
assign ece = ~ECE;  //complement 
assign ECF =  DDF & CFE  ; 
assign ecf = ~ECF;  //complement 
assign EEE =  DDE & CFG  ; 
assign eee = ~EEE;  //complement 
assign EEF =  DDF & CFF  ; 
assign eef = ~EEF;  //complement 
assign EEG =  DDG & CFE  ; 
assign eeg = ~EEG;  //complement 
assign EGF =  DDF & CFG  ; 
assign egf = ~EGF;  //complement 
assign EGG =  DDG & CFF  ; 
assign egg = ~EGG;  //complement 
assign EGH =  DDH & CFE  ; 
assign egh = ~EGH;  //complement 
assign faa = ~FAA;  //complement 
assign FBA = ~fba;  //complement 
assign tam = ~TAM;  //complement 
assign tar = ~TAR;  //complement 
assign tas = ~TAS;  //complement 
assign fec = ~FEC;  //complement 
assign FFC = ~ffc;  //complement 
assign fgb = ~FGB;  //complement 
assign FHB = ~fhb;  //complement 
assign EAA =  DDA & CFI  ; 
assign eaa = ~EAA;  //complement 
assign EAB =  DDB & CFH  ; 
assign eab = ~EAB;  //complement 
assign ECA =  DDA & CFJ  ; 
assign eca = ~ECA;  //complement 
assign ECB =  DDB & CFI  ; 
assign ecb = ~ECB;  //complement 
assign ECC =  DDC & CFH  ; 
assign ecc = ~ECC;  //complement 
assign EEB =  DDB & CFJ  ; 
assign eeb = ~EEB;  //complement 
assign EEC =  DDC & CFI  ; 
assign eec = ~EEC;  //complement 
assign EED =  DDD & CFH  ; 
assign eed = ~EED;  //complement 
assign EGE =  DDE & CFH  ; 
assign ege = ~EGE;  //complement 
assign EGC =  DDC & CFJ  ; 
assign egc = ~EGC;  //complement 
assign EGD =  DDD & CFE  ; 
assign egd = ~EGD;  //complement 
assign fga = ~FGA;  //complement 
assign FHA = ~fha;  //complement 
assign EEA =  DDA & CFK  ; 
assign eea = ~EEA;  //complement 
assign EGA =  DDA & CFL  ; 
assign ega = ~EGA;  //complement 
assign EGB =  DDB & CFK  ; 
assign egb = ~EGB;  //complement 
assign EIG =  DDG & CFG  ; 
assign eig = ~EIG;  //complement 
assign fea = ~FEA;  //complement 
assign qaa = ~QAA;  //complement 
assign qab = ~QAB;  //complement 
assign fcb = ~FCB;  //complement 
assign FDB = ~fdb;  //complement 
assign fid = ~FID;  //complement 
assign FJD = ~fjd;  //complement 
assign DDF = ~ddf;  //complement 
assign DDG = ~ddg;  //complement 
assign DDH = ~ddh;  //complement 
assign DDI = ~ddi;  //complement 
assign fke = ~FKE;  //complement 
assign FLE = ~fle;  //complement 
assign EIH =  DDH & CFF  ; 
assign eih = ~EIH;  //complement 
assign EII =  DDI & CFE  ; 
assign eii = ~EII;  //complement 
assign cfe = ~CFE;  //complement 
assign cff = ~CFF;  //complement 
assign cfg = ~CFG;  //complement 
assign EKH =  DGH & CCG  ; 
assign ekh = ~EKH;  //complement 
assign EKI =  DGI & CCF  ; 
assign eki = ~EKI;  //complement 
assign EKJ =  DDJ & CCE  ; 
assign ekj = ~EKJ;  //complement 
assign fic = ~FIC;  //complement 
assign FJC = ~fjc;  //complement 
assign ddb = ~DDB;  //complement 
assign ddc = ~DDC;  //complement 
assign ddd = ~DDD;  //complement 
assign dde = ~DDE;  //complement 
assign fkd = ~FKD;  //complement 
assign FLD = ~fld;  //complement 
assign EID =  DDD & CFJ  ; 
assign eid = ~EID;  //complement 
assign EIE =  DDE & CFI  ; 
assign eie = ~EIE;  //complement 
assign EIF =  DDF & CFH  ; 
assign eif = ~EIF;  //complement 
assign fkb = ~FKB;  //complement 
assign cfh = ~CFH;  //complement 
assign cfi = ~CFI;  //complement 
assign cfj = ~CFJ;  //complement 
assign EKE =  DGE & CCJ  ; 
assign eke = ~EKE;  //complement 
assign EKF =  DGF & CCI  ; 
assign ekf = ~EKF;  //complement 
assign EKG =  DGG & CCH  ; 
assign ekg = ~EKG;  //complement 
assign fib = ~FIB;  //complement 
assign FJB = ~fjb;  //complement 
assign fia = ~FIA;  //complement 
assign dda = ~DDA;  //complement 
assign fkc = ~FKC;  //complement 
assign FLC = ~flc;  //complement 
assign EIA =  DDA & CFM  ; 
assign eia = ~EIA;  //complement 
assign EIB =  DDB & CFL  ; 
assign eib = ~EIB;  //complement 
assign EIC =  DDC & CFK  ; 
assign eic = ~EIC;  //complement 
assign cfk = ~CFK;  //complement 
assign cfl = ~CFL;  //complement 
assign cfm = ~CFM;  //complement 
assign EKB =  DGB & CCM  ; 
assign ekb = ~EKB;  //complement 
assign EKC =  DGC & CCL  ; 
assign ekc = ~EKC;  //complement 
assign EKD =  DGD & CCK  ; 
assign ekd = ~EKD;  //complement 
assign qae = ~QAE;  //complement 
assign qaf = ~QAF;  //complement 
assign qai = ~QAI;  //complement 
assign fka = ~FKA;  //complement 
assign qac = ~QAC;  //complement 
assign qad = ~QAD;  //complement 
assign qag = ~QAG;  //complement 
assign qah = ~QAH;  //complement 
assign EKA =  DGA & CCN  ; 
assign eka = ~EKA;  //complement 
assign fmd = ~FMD;  //complement 
assign FND = ~fnd;  //complement 
assign foe = ~FOE;  //complement 
assign FPE = ~fpe;  //complement 
assign fqd = ~FQD;  //complement 
assign OGD = ~ogd;  //complement 
assign DDJ = ~ddj;  //complement 
assign DDK = ~ddk;  //complement 
assign DDL = ~ddl;  //complement 
assign DDM = ~ddm;  //complement 
assign EMI =  DGI & CCG  ; 
assign emi = ~EMI;  //complement 
assign EMJ =  DDJ & CCF  ; 
assign emj = ~EMJ;  //complement 
assign EMK =  DDK & CCE  ; 
assign emk = ~EMK;  //complement 
assign EOJ =  DDJ & CCG  ; 
assign eoj = ~EOJ;  //complement 
assign EOK =  DDK & CCF  ; 
assign eok = ~EOK;  //complement 
assign EOL =  DDL & CCE  ; 
assign eol = ~EOL;  //complement 
assign EQK =  DDK & CCG  ; 
assign eqk = ~EQK;  //complement 
assign EQL =  DDL & CCF  ; 
assign eql = ~EQL;  //complement 
assign EQM =  DDM & CCE  ; 
assign eqm = ~EQM;  //complement 
assign cce = ~CCE;  //complement 
assign ccf = ~CCF;  //complement 
assign ccg = ~CCG;  //complement 
assign fmc = ~FMC;  //complement 
assign FNC = ~fnc;  //complement 
assign fod = ~FOD;  //complement 
assign FPD = ~fpd;  //complement 
assign fqc = ~FQC;  //complement 
assign OGC = ~ogc;  //complement 
assign DGF = ~dgf;  //complement 
assign DGG = ~dgg;  //complement 
assign DGH = ~dgh;  //complement 
assign DGI = ~dgi;  //complement 
assign EMH =  DGH & CCH  ; 
assign emh = ~EMH;  //complement 
assign EMF =  DGF & CCJ  ; 
assign emf = ~EMF;  //complement 
assign EMG =  DGG & CCI  ; 
assign emg = ~EMG;  //complement 
assign EOG =  DGG & CCJ  ; 
assign eog = ~EOG;  //complement 
assign EOH =  DGH & CCI  ; 
assign eoh = ~EOH;  //complement 
assign EOI =  DGI & CCH  ; 
assign eoi = ~EOI;  //complement 
assign EQH =  DGH & CCJ  ; 
assign eqh = ~EQH;  //complement 
assign EQI =  DGI & CCI  ; 
assign eqi = ~EQI;  //complement 
assign EQJ =  DDJ & CCH  ; 
assign eqj = ~EQJ;  //complement 
assign cch = ~CCH;  //complement 
assign cci = ~CCI;  //complement 
assign ccj = ~CCJ;  //complement 
assign fmb = ~FMB;  //complement 
assign FNB = ~fnb;  //complement 
assign foc = ~FOC;  //complement 
assign FPC = ~fpc;  //complement 
assign fqb = ~FQB;  //complement 
assign OGB = ~ogb;  //complement 
assign dgb = ~DGB;  //complement 
assign dgc = ~DGC;  //complement 
assign dgd = ~DGD;  //complement 
assign dge = ~DGE;  //complement 
assign EME =  DGE & CCK  ; 
assign eme = ~EME;  //complement 
assign EMC =  DGC & CCM  ; 
assign emc = ~EMC;  //complement 
assign EMD =  DGD & CCL  ; 
assign emd = ~EMD;  //complement 
assign EOD =  DGD & CCM  ; 
assign eod = ~EOD;  //complement 
assign EOE =  DGE & CCL  ; 
assign eoe = ~EOE;  //complement 
assign EOF =  DGF & CCK  ; 
assign eof = ~EOF;  //complement 
assign EQE =  DGE & CCM  ; 
assign eqe = ~EQE;  //complement 
assign EQF =  DGF & CCL  ; 
assign eqf = ~EQF;  //complement 
assign EQG =  DGG & CCK  ; 
assign eqg = ~EQG;  //complement 
assign cck = ~CCK;  //complement 
assign ccl = ~CCL;  //complement 
assign ccm = ~CCM;  //complement 
assign fma = ~FMA;  //complement 
assign FNA = ~fna;  //complement 
assign fob = ~FOB;  //complement 
assign FPB = ~fpb;  //complement 
assign foa = ~FOA;  //complement 
assign fqa = ~FQA;  //complement 
assign OGA = ~oga;  //complement 
assign dga = ~DGA;  //complement 
assign qmm = ~QMM;  //complement 
assign qmr = ~QMR;  //complement 
assign qms = ~QMS;  //complement 
assign EMB =  DGB & CCN  ; 
assign emb = ~EMB;  //complement 
assign EMA =  DGA & CCO  ; 
assign ema = ~EMA;  //complement 
assign EOA =  DGA & CCP  ; 
assign eoa = ~EOA;  //complement 
assign EOB =  DGB & CCO  ; 
assign eob = ~EOB;  //complement 
assign EOC =  DGC & CCN  ; 
assign eoc = ~EOC;  //complement 
assign EQB =  DGB & CCP  ; 
assign eqb = ~EQB;  //complement 
assign EQC =  DGC & CCO  ; 
assign eqc = ~EQC;  //complement 
assign EQD =  DGD & CCN  ; 
assign eqd = ~EQD;  //complement 
assign ccn = ~CCN;  //complement 
assign cco = ~CCO;  //complement 
assign ccp = ~CCP;  //complement 
assign iaa = ~IAA; //complement 
assign iab = ~IAB; //complement 
assign iac = ~IAC; //complement 
assign iad = ~IAD; //complement 
assign iae = ~IAE; //complement 
assign iaf = ~IAF; //complement 
assign iag = ~IAG; //complement 
assign iah = ~IAH; //complement 
assign iai = ~IAI; //complement 
assign iaj = ~IAJ; //complement 
assign iak = ~IAK; //complement 
assign ial = ~IAL; //complement 
assign iam = ~IAM; //complement 
assign ian = ~IAN; //complement 
assign iao = ~IAO; //complement 
assign iap = ~IAP; //complement 
assign iba = ~IBA; //complement 
assign ibb = ~IBB; //complement 
assign ibc = ~IBC; //complement 
assign ibd = ~IBD; //complement 
assign ibe = ~IBE; //complement 
assign ibf = ~IBF; //complement 
assign ibg = ~IBG; //complement 
assign ibh = ~IBH; //complement 
assign ibi = ~IBI; //complement 
assign ibj = ~IBJ; //complement 
assign ibk = ~IBK; //complement 
assign ibl = ~IBL; //complement 
assign ibm = ~IBM; //complement 
assign ibn = ~IBN; //complement 
assign ibo = ~IBO; //complement 
assign ibp = ~IBP; //complement 
assign ica = ~ICA; //complement 
assign icb = ~ICB; //complement 
assign icc = ~ICC; //complement 
assign icd = ~ICD; //complement 
assign ice = ~ICE; //complement 
assign icf = ~ICF; //complement 
assign icg = ~ICG; //complement 
assign ich = ~ICH; //complement 
assign ici = ~ICI; //complement 
assign icj = ~ICJ; //complement 
assign ick = ~ICK; //complement 
assign icl = ~ICL; //complement 
assign icm = ~ICM; //complement 
assign icn = ~ICN; //complement 
assign ico = ~ICO; //complement 
assign icp = ~ICP; //complement 
assign ida = ~IDA; //complement 
assign idb = ~IDB; //complement 
assign idc = ~IDC; //complement 
assign idd = ~IDD; //complement 
assign ide = ~IDE; //complement 
assign idf = ~IDF; //complement 
assign idg = ~IDG; //complement 
assign idh = ~IDH; //complement 
assign idi = ~IDI; //complement 
assign idj = ~IDJ; //complement 
assign idk = ~IDK; //complement 
assign idl = ~IDL; //complement 
assign idm = ~IDM; //complement 
assign idn = ~IDN; //complement 
assign ido = ~IDO; //complement 
assign idp = ~IDP; //complement 
assign iea = ~IEA; //complement 
assign ieb = ~IEB; //complement 
assign iec = ~IEC; //complement 
assign ied = ~IED; //complement 
assign iee = ~IEE; //complement 
assign ief = ~IEF; //complement 
assign ieg = ~IEG; //complement 
assign ieh = ~IEH; //complement 
assign iei = ~IEI; //complement 
assign iej = ~IEJ; //complement 
assign iek = ~IEK; //complement 
assign iel = ~IEL; //complement 
assign iem = ~IEM; //complement 
assign ien = ~IEN; //complement 
assign ieo = ~IEO; //complement 
assign iep = ~IEP; //complement 
assign ieq = ~IEQ; //complement 
assign ier = ~IER; //complement 
assign ies = ~IES; //complement 
assign iet = ~IET; //complement 
assign ieu = ~IEU; //complement 
assign iev = ~IEV; //complement 
assign iew = ~IEW; //complement 
assign iex = ~IEX; //complement 
assign iey = ~IEY; //complement 
assign iez = ~IEZ; //complement 
assign ifa = ~IFA; //complement 
assign ifb = ~IFB; //complement 
assign ifc = ~IFC; //complement 
assign ifd = ~IFD; //complement 
assign ife = ~IFE; //complement 
assign ifff  = ~IFFF ; //complement 
assign ifg = ~IFG; //complement 
assign ifh = ~IFH; //complement 
assign ifi = ~IFI; //complement 
assign ifj = ~IFJ; //complement 
assign ifk = ~IFK; //complement 
assign ifl = ~IFL; //complement 
assign ifm = ~IFM; //complement 
assign ifn = ~IFN; //complement 
assign ifo = ~IFO; //complement 
assign ifp = ~IFP; //complement 
assign iga = ~IGA; //complement 
assign iha = ~IHA; //complement 
assign ika = ~IKA; //complement 
assign imm = ~IMM; //complement 
assign imr = ~IMR; //complement 
assign ims = ~IMS; //complement 
assign ira = ~IRA; //complement 
assign isa = ~ISA; //complement 
assign ita = ~ITA; //complement 
always@(posedge IZZ )
   begin 
 FAN <=  EBO & ebp & ebq  |  ebo & EBP & ebq  |  ebo & ebp & EBQ  |  EBO & EBP & EBQ  ;
 fbn <=  EBO & ebp & ebq  |  ebo & EBP & ebq  |  ebo & ebp & EBQ  |  ebo & ebp & ebq  ;
 FCO <=  EDP & edq & edr  |  edp & EDQ & edr  |  edp & edq & EDR  |  EDP & EDQ & EDR  ;
 fdo <=  EDP & edq & edr  |  edp & EDQ & edr  |  edp & edq & EDR  |  edp & edq & edr  ;
 FEP <=  EFQ & efr & efs  |  efq & EFR & efs  |  efq & efr & EFS  |  EFQ & EFR & EFS  ;
 ffp <=  EFQ & efr & efs  |  efq & EFR & efs  |  efq & efr & EFS  |  efq & efr & efs  ;
 FGO <=  EHR & ehs & eht  |  ehr & EHS & eht  |  ehr & ehs & EHT  |  EHR & EHS & EHT  ;
 fho <=  EHR & ehs & eht  |  ehr & EHS & eht  |  ehr & ehs & EHT  |  ehr & ehs & eht  ;
 FEM <=  EFH & efi & efj  |  efh & EFI & efj  |  efh & efi & EFJ  |  EFH & EFI & EFJ  ;
 ffm <=  EFH & efi & efj  |  efh & EFI & efj  |  efh & efi & EFJ  |  efh & efi & efj  ;
 FAM <=  EBL & ebm & ebn  |  ebl & EBM & ebn  |  ebl & ebm & EBN  |  EBL & EBM & EBN  ;
 fbm <=  EBL & ebm & ebn  |  ebl & EBM & ebn  |  ebl & ebm & EBN  |  ebl & ebm & ebn  ;
 FCN <=  EDM & edn & edo  |  edm & EDN & edo  |  edm & edn & EDO  |  EDM & EDN & EDO  ;
 fdn <=  EDM & edn & edo  |  edm & EDN & edo  |  edm & edn & EDO  |  edm & edn & edo  ;
 FEO <=  EFN & efo & efp  |  efn & EFO & efp  |  efn & efo & EFP  |  EFN & EFO & EFP  ;
 ffo <=  EFN & efo & efp  |  efn & EFO & efp  |  efn & efo & EFP  |  efn & efo & efp  ;
 FGN <=  EHO & ehp & ehq  |  eho & EHP & ehq  |  eho & ehp & EHQ  |  EHO & EHP & EHQ  ;
 fhn <=  EHO & ehp & ehq  |  eho & EHP & ehq  |  eho & ehp & EHQ  |  eho & ehp & ehq  ;
 FAL <=  EBI & ebj & ebk  |  ebi & EBJ & ebk  |  ebi & ebj & EBK  |  EBI & EBJ & EBK  ;
 fbl <=  EBI & ebj & ebk  |  ebi & EBJ & ebk  |  ebi & ebj & EBK  |  ebi & ebj & ebk  ;
 FCM <=  EDJ & edk & edl  |  edj & EDK & edl  |  edj & edk & EDL  |  EDJ & EDK & EDL  ;
 fdm <=  EDJ & edk & edl  |  edj & EDK & edl  |  edj & edk & EDL  |  edj & edk & edl  ;
 FGM <=  EHL & ehm & ehn  |  ehl & EHM & ehn  |  ehl & ehm & EHN  |  EHL & EHM & EHN  ;
 fhm <=  EHL & ehm & ehn  |  ehl & EHM & ehn  |  ehl & ehm & EHN  |  ehl & ehm & ehn  ;
 FAK <=  EBF & ebg & ebh  |  ebf & EBG & ebh  |  ebf & ebg & EBH  |  EBF & EBG & EBH  ;
 fbk <=  EBF & ebg & ebh  |  ebf & EBG & ebh  |  ebf & ebg & EBH  |  ebf & ebg & ebh  ;
 FCL <=  EDG & edh & edi  |  edg & EDH & edi  |  edg & edh & EDI  |  EDG & EDH & EDI  ;
 fdl <=  EDG & edh & edi  |  edg & EDH & edi  |  edg & edh & EDI  |  edg & edh & edi  ;
 FGL <=  EHI & ehj & ehk  |  ehi & EHJ & ehk  |  ehi & ehj & EHK  |  EHI & EHJ & EHK  ;
 fhl <=  EHI & ehj & ehk  |  ehi & EHJ & ehk  |  ehi & ehj & EHK  |  ehi & ehj & ehk  ;
 cda <= tra & iaa ; 
 CDB <= tra & IAB ; 
 CDC <= tra & IAC ; 
 FIP <=  EJS & ejt & eju  |  ejs & EJT & eju  |  ejs & ejt & EJU  |  EJS & EJT & EJU  ;
 fjp <=  EJS & ejt & eju  |  ejs & EJT & eju  |  ejs & ejt & EJU  |  ejs & ejt & eju  ;
 DCJ <= IFJ ; 
 DCK <= IFK ; 
 DCL <= IFL ; 
 DCM <= IFM ; 
 FKQ <=  ELT & elu & elv  |  elt & ELU & elv  |  elt & elu & ELV  |  ELT & ELU & ELV  ;
 flq <=  ELT & elu & elv  |  elt & ELU & elv  |  elt & elu & ELV  |  elt & elu & elv  ;
 CDD <= IAD ; 
 CDE <= IAE ; 
 CDF <= IAF ; 
 FEN <=  EFK & efl & efm  |  efk & EFL & efm  |  efk & efl & EFM  |  EFK & EFL & EFM  ;
 ffn <=  EFK & efl & efm  |  efk & EFL & efm  |  efk & efl & EFM  |  efk & efl & efm  ;
 FIO <=  EJP & ejq & ejr  |  ejp & EJQ & ejr  |  ejp & ejq & EJR  |  EJP & EJQ & EJR  ;
 fjo <=  EJP & ejq & ejr  |  ejp & EJQ & ejr  |  ejp & ejq & EJR  |  ejp & ejq & ejr  ;
 DCF <= IFFF  ; 
 DCG <= IFG ; 
 DCH <= IFH ; 
 DCI <= IFI ; 
 FKP <=  ELQ & elr & els  |  elq & ELR & els  |  elq & elr & ELS  |  ELQ & ELR & ELS  ;
 flp <=  ELQ & elr & els  |  elq & ELR & els  |  elq & elr & ELS  |  elq & elr & els  ;
 CDG <= IAG ; 
 CDH <= IAH ; 
 CDI <= IAI ; 
 FIN <=  EJM & ejn & ejo  |  ejm & EJN & ejo  |  ejm & ejn & EJO  |  EJM & EJN & EJO  ;
 fjn <=  EJM & ejn & ejo  |  ejm & EJN & ejo  |  ejm & ejn & EJO  |  ejm & ejn & ejo  ;
 DCB <= IFB ; 
 DCD <= IFD ; 
 DCC <= IFC ; 
 DCE <= IFE ; 
 FKO <=  ELN & elo & elp  |  eln & ELO & elp  |  eln & elo & ELP  |  ELN & ELO & ELP  ;
 flo <=  ELN & elo & elp  |  eln & ELO & elp  |  eln & elo & ELP  |  eln & elo & elp  ;
 CDJ <= IAJ ; 
 CDK <= IAK ; 
 CDL <= IAL ; 
 FIM <=  EJJ & ejk & ejl  |  ejj & EJK & ejl  |  ejj & ejk & EJL  |  EJJ & EJK & EJL  ;
 fjm <=  EJJ & ejk & ejl  |  ejj & EJK & ejl  |  ejj & ejk & EJL  |  ejj & ejk & ejl  ;
 DBN <= BAN ; 
 DBO <= BAO ; 
 DBP <= BAP ; 
 DCA <= IFA ; 
 FKN <=  ELK & ell & elm  |  elk & ELL & elm  |  elk & ell & ELM  |  ELK & ELL & ELM  ;
 fln <=  ELK & ell & elm  |  elk & ELL & elm  |  elk & ell & ELM  |  elk & ell & elm  ;
 caa <= tra & iaa ; 
 CAB <= tra & IAB ; 
 CAC <= tra & IAC ; 
 FMP <=  ENU & env & enw  |  enu & ENV & enw  |  enu & env & ENW  |  ENU & ENV & ENW  ;
 fnp <=  ENU & env & enw  |  enu & ENV & enw  |  enu & env & ENW  |  enu & env & enw  ;
 FOQ <=  EPV & epw & epx  |  epv & EPW & epx  |  epv & epw & EPX  |  EPV & EPW & EPX  ;
 fpq <=  EPV & epw & epx  |  epv & EPW & epx  |  epv & epw & EPX  |  epv & epw & epx  ;
 FQP <=  ERW & erx & qai  |  erw & ERX & qai  |  erw & erx & QAI  |  ERW & ERX & QAI  ;
 ogp <=  ERW & erx & qai  |  erw & ERX & qai  |  erw & erx & QAI  |  erw & erx & qai  ;
 DIN <= IFN ; 
 DIO <= IFO ; 
 DIP <= IFP ; 
 CAD <= IAD ; 
 CAE <= IAE ; 
 CAF <= IAF ; 
 FMO <=  ENR & ens & ent  |  enr & ENS & ent  |  enr & ens & ENT  |  ENR & ENS & ENT  ;
 fno <=  ENR & ens & ent  |  enr & ENS & ent  |  enr & ens & ENT  |  enr & ens & ent  ;
 FOP <=  EPS & ept & epu  |  eps & EPT & epu  |  eps & ept & EPU  |  EPS & EPT & EPU  ;
 fpp <=  EPS & ept & epu  |  eps & EPT & epu  |  eps & ept & EPU  |  eps & ept & epu  ;
 FQO <=  ERT & eru & erv  |  ert & ERU & erv  |  ert & eru & ERV  |  ERT & ERU & ERV  ;
 ogo <=  ERT & eru & erv  |  ert & ERU & erv  |  ert & eru & ERV  |  ert & eru & erv  ;
 DIJ <= IFJ ; 
 DIK <= IFK ; 
 DIL <= IFL ; 
 DIM <= IFM ; 
 CAG <= IAG ; 
 CAH <= IAH ; 
 CAI <= IAI ; 
 FMN <=  ENO & enp & enq  |  eno & ENP & enq  |  eno & enp & ENQ  |  ENO & ENP & ENQ  ;
 fnn <=  ENO & enp & enq  |  eno & ENP & enq  |  eno & enp & ENQ  |  eno & enp & enq  ;
 FOO <=  EPP & epq & epr  |  epp & EPQ & epr  |  epp & epq & EPR  |  EPP & EPQ & EPR  ;
 fpo <=  EPP & epq & epr  |  epp & EPQ & epr  |  epp & epq & EPR  |  epp & epq & epr  ;
 FQN <=  ERQ & err & ers  |  erq & ERR & ers  |  erq & err & ERS  |  ERQ & ERR & ERS  ;
 ogn <=  ERQ & err & ers  |  erq & ERR & ers  |  erq & err & ERS  |  erq & err & ers  ;
 DIF <= IFFF  ; 
 DIG <= IFG ; 
 DIH <= IFH ; 
 DII <= IFE ; 
 CAJ <= IAJ ; 
 CAK <= IAK ; 
 CAL <= IAL ; 
 FMM <=  ENL & enm & enn  |  enl & ENM & enn  |  enl & enm & ENN  |  ENL & ENM & ENN  ;
 fnm <=  ENL & enm & enn  |  enl & ENM & enn  |  enl & enm & ENN  |  enl & enm & enn  ;
 FON <=  EPM & epn & epo  |  epm & EPN & epo  |  epm & epn & EPO  |  EPM & EPN & EPO  ;
 fpn <=  EPM & epn & epo  |  epm & EPN & epo  |  epm & epn & EPO  |  epm & epn & epo  ;
 FQM <=  ERN & ero & erp  |  ern & ERO & erp  |  ern & ero & ERP  |  ERN & ERO & ERP  ;
 ogm <=  ERN & ero & erp  |  ern & ERO & erp  |  ern & ero & ERP  |  ern & ero & erp  ;
 DIC <= IFC ; 
 DID <= IFD ; 
 DIE <= IFE ; 
 FAJ <=  EBC & ebd & ebe  |  ebc & EBD & ebe  |  ebc & ebd & EBE  |  EBC & EBD & EBE  ;
 fbj <=  EBC & ebd & ebe  |  ebc & EBD & ebe  |  ebc & ebd & EBE  |  ebc & ebd & ebe  ;
 FCK <=  EDD & ede & edf  |  edd & EDE & edf  |  edd & ede & EDF  |  EDD & EDE & EDF  ;
 fdk <=  EDD & ede & edf  |  edd & EDE & edf  |  edd & ede & EDF  |  edd & ede & edf  ;
 FEL <=  EFE & eff & efg  |  efe & EFF & efg  |  efe & eff & EFG  |  EFE & EFF & EFG  ;
 ffl <=  EFE & eff & efg  |  efe & EFF & efg  |  efe & eff & EFG  |  efe & eff & efg  ;
 FGK <=  EHF & ehg & ehh  |  ehf & EHG & ehh  |  ehf & ehg & EHH  |  EHF & EHG & EHH  ;
 fhk <=  EHF & ehg & ehh  |  ehf & EHG & ehh  |  ehf & ehg & EHH  |  ehf & ehg & ehh  ;
 FAI <=  EAX & eba & ebb  |  eax & EBA & ebb  |  eax & eba & EBB  |  EAX & EBA & EBB  ;
 fbi <=  EAX & eba & ebb  |  eax & EBA & ebb  |  eax & eba & EBB  |  eax & eba & ebb  ;
 FEK <=  EFB & efc & efd  |  efb & EFC & efd  |  efb & efc & EFD  |  EFB & EFC & EFD  ;
 ffk <=  EFB & efc & efd  |  efb & EFC & efd  |  efb & efc & EFD  |  efb & efc & efd  ;
 FGJ <=  EHC & ehd & ehe  |  ehc & EHD & ehe  |  ehc & ehd & EHE  |  EHC & EHD & EHE  ;
 fhj <=  EHC & ehd & ehe  |  ehc & EHD & ehe  |  ehc & ehd & EHE  |  ehc & ehd & ehe  ;
 FAH <=  EAU & eav & eaw  |  eau & EAV & eaw  |  eau & eav & EAW  |  EAU & EAV & EAW  ;
 fbh <=  EAU & eav & eaw  |  eau & EAV & eaw  |  eau & eav & EAW  |  eau & eav & eaw  ;
 FCI <=  ECV & ecw & ecx  |  ecv & ECW & ecx  |  ecv & ecw & ECX  |  ECV & ECW & ECX  ;
 fdi <=  ECV & ecw & ecx  |  ecv & ECW & ecx  |  ecv & ecw & ECX  |  ecv & ecw & ecx  ;
 FEJ <=  EEW & eex & efa  |  eew & EEX & efa  |  eew & eex & EFA  |  EEW & EEX & EFA  ;
 ffj <=  EEW & eex & efa  |  eew & EEX & efa  |  eew & eex & EFA  |  eew & eex & efa  ;
 FGI <=  EGX & eha & ehb  |  egx & EHA & ehb  |  egx & eha & EHB  |  EGX & EHA & EHB  ;
 fhi <=  EGX & eha & ehb  |  egx & EHA & ehb  |  egx & eha & EHB  |  egx & eha & ehb  ;
 FAG <=  EAR & eas & eat  |  ear & EAS & eat  |  ear & eas & EAT  |  EAR & EAS & EAT  ;
 fbg <=  EAR & eas & eat  |  ear & EAS & eat  |  ear & eas & EAT  |  ear & eas & eat  ;
 FCH <=  ECS & ect & ecu  |  ecs & ECT & ecu  |  ecs & ect & ECU  |  ECS & ECT & ECU  ;
 fdh <=  ECS & ect & ecu  |  ecs & ECT & ecu  |  ecs & ect & ECU  |  ecs & ect & ecu  ;
 FCJ <=  EDA & edb & edc  |  eda & EDB & edc  |  eda & edb & EDC  |  EDA & EDB & EDC  ;
 fdj <=  EDA & edb & edc  |  eda & EDB & edc  |  eda & edb & EDC  |  eda & edb & edc  ;
 FGH <=  EGU & egv & egw  |  egu & EGV & egw  |  egu & egv & EGW  |  EGU & EGV & EGW  ;
 fhh <=  EGU & egv & egw  |  egu & EGV & egw  |  egu & egv & EGW  |  egu & egv & egw  ;
 FIL <=  EJG & ejh & eji  |  ejg & EJH & eji  |  ejg & ejh & EJI  |  EJG & EJH & EJI  ;
 fjl <=  EJG & ejh & eji  |  ejg & EJH & eji  |  ejg & ejh & EJI  |  ejg & ejh & eji  ;
 den <= ban ; 
 deo <= bao ; 
 dep <= bap ; 
 dfa <= ifa ; 
 FKM <=  ELH & eli & elj  |  elh & ELI & elj  |  elh & eli & ELJ  |  ELH & ELI & ELJ  ;
 flm <=  ELH & eli & elj  |  elh & ELI & elj  |  elh & eli & ELJ  |  elh & eli & elj  ;
 DHK <= BAK ; 
 DHL <= BAL ; 
 CDM <= IAM ; 
 CDN <= IAN ; 
 CDO <= IAO ; 
 FII <=  EIV & eiw & eix  |  eiv & EIW & eix  |  eiv & eiw & EIX  |  EIV & EIW & EIX  ;
 fji <=  EIV & eiw & eix  |  eiv & EIW & eix  |  eiv & eiw & EIX  |  eiv & eiw & eix  ;
 FIK <=  EJD & eje & ejf  |  ejd & EJE & ejf  |  ejd & eje & EJF  |  EJD & EJE & EJF  ;
 fjk <=  EJD & eje & ejf  |  ejd & EJE & ejf  |  ejd & eje & EJF  |  ejd & eje & ejf  ;
 DEJ <= BAJ ; 
 DEK <= BAK ; 
 DEL <= BAL ; 
 DEM <= BAM ; 
 FKL <=  ELE & elf & elg  |  ele & ELF & elg  |  ele & elf & ELG  |  ELE & ELF & ELG  ;
 fll <=  ELE & elf & elg  |  ele & ELF & elg  |  ele & elf & ELG  |  ele & elf & elg  ;
 OBB <=  ICA & TSD  |  BAA & TKD  |  AAB & THD  ; 
 CDP <= IAP ; 
 CEA <= AAA ; 
 CEB <= AAB ; 
 FIJ <=  EJA & ejb & ejc  |  eja & EJB & ejc  |  eja & ejb & EJC  |  EJA & EJB & EJC  ;
 fjj <=  EJA & ejb & ejc  |  eja & EJB & ejc  |  eja & ejb & EJC  |  eja & ejb & ejc  ;
 DEF <= BAF ; 
 DEG <= BAG ; 
 DEH <= BAH ; 
 DEI <= BAI ; 
 FKK <=  ELB & elc & eld  |  elb & ELC & eld  |  elb & elc & ELD  |  ELB & ELC & ELD  ;
 flk <=  ELB & elc & eld  |  elb & ELC & eld  |  elb & elc & ELD  |  elb & elc & eld  ;
 CEC <= AAC ; 
 CED <= AAD ; 
 CEE <= AAE ; 
 CEF <= AAF & TRA |  AAF & tra ; 
 CEG <= IEA & TRA |  AAG & tra ; 
 CEH <= IEB & TRA |  AAH & tra ; 
 FEI <=  EET & eeu & eev  |  eet & EEU & eev  |  eet & eeu & EEV  |  EET & EEU & EEV  ;
 ffi <=  EET & eeu & eev  |  eet & EEU & eev  |  eet & eeu & EEV  |  eet & eeu & eev  ;
 DEB <= BAB ; 
 DEC <= BAC ; 
 DED <= BAD ; 
 DEE <= BAE ; 
 FKJ <=  EKW & ekx & ela  |  ekw & EKX & ela  |  ekw & ekx & ELA  |  EKW & EKX & ELA  ;
 flj <=  EKW & ekx & ela  |  ekw & EKX & ela  |  ekw & ekx & ELA  |  ekw & ekx & ela  ;
 AAD <=  ICD & TSB  |  BAD & TKB  |  AAD & THB  ; 
 FML <=  ENI & enj & enk  |  eni & ENJ & enk  |  eni & enj & ENK  |  ENI & ENJ & ENK  ;
 fnl <=  ENI & enj & enk  |  eni & ENJ & enk  |  eni & enj & ENK  |  eni & enj & enk  ;
 FOM <=  EPJ & epk & epl  |  epj & EPK & epl  |  epj & epk & EPL  |  EPJ & EPK & EPL  ;
 fpm <=  EPJ & epk & epl  |  epj & EPK & epl  |  epj & epk & EPL  |  epj & epk & epl  ;
 FQL <=  ERK & erl & erm  |  erk & ERL & erm  |  erk & erl & ERM  |  ERK & ERL & ERM  ;
 ogl <=  ERK & erl & erm  |  erk & ERL & erm  |  erk & erl & ERM  |  erk & erl & erm  ;
 dfb <= ifb ; 
 dfc <= ifc ; 
 dfd <= ifd ; 
 dfe <= ife ; 
 CAM <= IAM ; 
 CAN <= IAN ; 
 CAO <= IAO ; 
 FMK <=  ENF & eng & enh  |  enf & ENG & enh  |  enf & eng & ENH  |  ENF & ENG & ENH  ;
 fnk <=  ENF & eng & enh  |  enf & ENG & enh  |  enf & eng & ENH  |  enf & eng & enh  ;
 FOL <=  EPG & eph & epi  |  epg & EPH & epi  |  epg & eph & EPI  |  EPG & EPH & EPI  ;
 fpl <=  EPG & eph & epi  |  epg & EPH & epi  |  epg & eph & EPI  |  epg & eph & epi  ;
 FQK <=  ERH & eri & erj  |  erh & ERI & erj  |  erh & eri & ERJ  |  ERH & ERI & ERJ  ;
 ogk <=  ERH & eri & erj  |  erh & ERI & erj  |  erh & eri & ERJ  |  erh & eri & erj  ;
 dhn <= ban ; 
 dho <= bao ; 
 dhp <= bap ; 
 dia <= ifa ; 
 CAP <= IAP ; 
 CBA <= AAA ; 
 CBB <= AAB ; 
 FMJ <=  ENC & endd & ene  |  enc & ENDD  & ene  |  enc & endd & ENE  |  ENC & ENDD  & ENE  ;
 fnj <=  ENC & endd & ene  |  enc & ENDD  & ene  |  enc & endd & ENE  |  enc & endd & ene  ;
 FOK <=  EPD & epe & epf  |  epd & EPE & epf  |  epd & epe & EPF  |  EPD & EPE & EPF  ;
 fpk <=  EPD & epe & epf  |  epd & EPE & epf  |  epd & epe & EPF  |  epd & epe & epf  ;
 FQJ <=  ERE & erf & erg  |  ere & ERF & erg  |  ere & erf & ERG  |  ERE & ERF & ERG  ;
 ogj <=  ERE & erf & erg  |  ere & ERF & erg  |  ere & erf & ERG  |  ere & erf & erg  ;
 DHJ <= BAJ ; 
 DHM <= BAM ; 
 CBC <= AAC ; 
 CBD <= AAD ; 
 CBE <= AAE ; 
 FMI <=  EMX & ena & enb  |  emx & ENA & enb  |  emx & ena & ENB  |  EMX & ENA & ENB  ;
 fni <=  EMX & ena & enb  |  emx & ENA & enb  |  emx & ena & ENB  |  emx & ena & enb  ;
 FOJ <=  EPA & epb & epc  |  epa & EPB & epc  |  epa & epb & EPC  |  EPA & EPB & EPC  ;
 fpj <=  EPA & epb & epc  |  epa & EPB & epc  |  epa & epb & EPC  |  epa & epb & epc  ;
 FQI <=  ERB & erc & erd  |  erb & ERC & erd  |  erb & erc & ERD  |  ERB & ERC & ERD  ;
 ogi <=  ERB & erc & erd  |  erb & ERC & erd  |  erb & erc & ERD  |  erb & erc & erd  ;
 TRA <= QRA ; 
 DHG <= BAG ; 
 DHH <= BAH ; 
 DHI <= BAI ; 
 CBF <= AAF & TRA |  AAF & tra ; 
 CBG <= IEA & TRA |  AAG & tra ; 
 CBH <= IEB & TRA |  AAH & tra ; 
 HCC <=  GCF & gch & fcf  |  gcf & GCH & fcf  |  gcf & gch & FCF  |  GCF & GCH & FCF  ;
 hdc <=  GCF & gch & fcf  |  gcf & GCH & fcf  |  gcf & gch & FCF  |  gcf & gch & fcf  ;
 HCB <=  GCD & gca & fca  |  gcd & GCA & fca  |  gcd & gca & FCA  |  GCD & GCA & FCA  ;
 hdb <=  GCD & gca & fca  |  gcd & GCA & fca  |  gcd & gca & FCA  |  gcd & gca & fca  ;
 HEB <=  GEE & geb & gdd  |  gee & GEB & gdd  |  gee & geb & GDD  |  GEE & GEB & GDD  ;
 hfb <=  GEE & geb & gdd  |  gee & GEB & gdd  |  gee & geb & GDD  |  gee & geb & gdd  ;
 HGB <=  GGD & gga & gfb  |  ggd & GGA & gfb  |  ggd & gga & GFB  |  GGD & GGA & GFB  ;
 hhb <=  GGD & gga & gfb  |  ggd & GGA & gfb  |  ggd & gga & GFB  |  ggd & gga & gfb  ;
 HIH <= GHH ; 
 HAB <=  FAD & gac & gab  |  fad & GAC & gab  |  fad & gac & GAB  |  FAD & GAC & GAB  ;
 hbb <=  FAD & gac & gab  |  fad & GAC & gab  |  fad & gac & GAB  |  fad & gac & gab  ;
 HED <=  GDC & ged & gef  |  gdc & GED & gef  |  gdc & ged & GEF  |  GDC & GED & GEF  ;
 hfd <=  GDC & ged & gef  |  gdc & GED & gef  |  gdc & ged & GEF  |  gdc & ged & gef  ;
 HGD <=  GFA & gge & gff  |  gfa & GGE & gff  |  gfa & gge & GFF  |  GFA & GGE & GFF  ;
 hhd <=  GFA & gge & gff  |  gfa & GGE & gff  |  gfa & gge & GFF  |  gfa & gge & gff  ;
 HID <=  GIF & ghc & gid  |  gif & GHC & gid  |  gif & ghc & GID  |  GIF & GHC & GID  ;
 hjd <=  GIF & ghc & gid  |  gif & GHC & gid  |  gif & ghc & GID  |  gif & ghc & gid  ;
 HIB <=  GHD & gie & gib  |  ghd & GIE & gib  |  ghd & gie & GIB  |  GHD & GIE & GIB  ;
 hjb <=  GHD & gie & gib  |  ghd & GIE & gib  |  ghd & gie & GIB  |  ghd & gie & gib  ;
 HMB <=  GLG & gmg & gli  |  glg & GMG & gli  |  glg & gmg & GLI  |  GLG & GMG & GLI  ;
 hnb <=  GLG & gmg & gli  |  glg & GMG & gli  |  glg & gmg & GLI  |  glg & gmg & gli  ;
 HOB <=  GOH & gng & gni  |  goh & GNG & gni  |  goh & gng & GNI  |  GOH & GNG & GNI  ;
 hpb <=  GOH & gng & gni  |  goh & GNG & gni  |  goh & gng & GNI  |  goh & gng & gni  ;
 HKB <=  GJE & gke & gkb  |  gje & GKE & gkb  |  gje & gke & GKB  |  GJE & GKE & GKB  ;
 hlb <=  GJE & gke & gkb  |  gje & GKE & gkb  |  gje & gke & GKB  |  gje & gke & gkb  ;
 HKG <=  GJD & gkd & gka  |  gjd & GKD & gka  |  gjd & gkd & GKA  |  GJD & GKD & GKA  ;
 hlg <=  GJD & gkd & gka  |  gjd & GKD & gka  |  gjd & gkd & GKA  |  gjd & gkd & gka  ;
 HKD <=  GKF & gji & gja  |  gkf & GJI & gja  |  gkf & gji & GJA  |  GKF & GJI & GJA  ;
 hld <=  GKF & gji & gja  |  gkf & GJI & gja  |  gkf & gji & GJA  |  gkf & gji & gja  ;
 HMD <=  GLD & gmf & gma  |  gld & GMF & gma  |  gld & gmf & GMA  |  GLD & GMF & GMA  ;
 hnd <=  GLD & gmf & gma  |  gld & GMF & gma  |  gld & gmf & GMA  |  gld & gmf & gma  ;
 HOD <=  GOG & gnd & goe  |  gog & GND & goe  |  gog & gnd & GOE  |  GOG & GND & GOE  ;
 hpd <=  GOG & gnd & goe  |  gog & GND & goe  |  gog & gnd & GOE  |  gog & gnd & goe  ;
 OHH <=  GRH & gre & grb  |  grh & GRE & grb  |  grh & gre & GRB  |  GRH & GRE & GRB  ;
 oih <=  GRH & gre & grb  |  grh & GRE & grb  |  grh & gre & GRB  |  grh & gre & grb  ;
 AAB <=  ICB & TSA  |  BAB & TKA  |  AAB & THA  ; 
 OBA <=  ICA & TSC  |  BAA & TKC  |  AAA & THC  ; 
 BDA <= BCA ; 
 BDB <= BCB ; 
 BEA <= BDA ; 
 BEB <= BDB ; 
 OAB <=  ICB & TSD  |  BAA & TKD  |  AAB & THD  ; 
 HQB <=  GQG & gph & gpj  |  gqg & GPH & gpj  |  gqg & gph & GPJ  |  GQG & GPH & GPJ  ;
 ohb <=  GQG & gph & gpj  |  gqg & GPH & gpj  |  gqg & gph & GPJ  |  gqg & gph & gpj  ;
 QGA <= IGA ; 
 QHA <= IHA ; 
 QKA <= IKA ; 
 bba <= ida ; 
 bbb <= idb ; 
 BCA <= BBA ; 
 BCB <= BBB ; 
 ODA <=  IDA & TTC  |  BEA & TGC  ; 
 OEA <=  IDA & TTC  |  BEA & TGC  ; 
 OHI <=  GRI & grd & grg  |  gri & GRD & grg  |  gri & grd & GRG  |  GRI & GRD & GRG  ;
 oii <=  GRI & grd & grg  |  gri & GRD & grg  |  gri & grd & GRG  |  gri & grd & grg  ;
 OHK <= GRA ; 
 BAA <=  IDA & TTA  |  BEA & TGA  ; 
 BAB <=  IDB & TTA  |  BEB & TGA  ; 
 ODB <=  IDB & TTD  |  BEB & TGD  ; 
 OEB <=  IDB & TTD  |  BEB & TGD  ; 
 OBD <=  ICD & TSF  |  BAD & TKF  |  AAD & THF  ; 
 BAC <=  IDC & TTB  |  BEC & TGB  ; 
 BAD <=  IDD & TTB  |  BED & TGB  ; 
 ODD <=  IDD & TTF  |  BED & TGF  ; 
 OED <=  IDD & TTF  |  BED & TGF  ; 
 HQD <=  GPE & gqd & gqf  |  gpe & GQD & gqf  |  gpe & gqd & GQF  |  GPE & GQD & GQF  ;
 ohd <=  GPE & gqd & gqf  |  gpe & GQD & gqf  |  gpe & gqd & GQF  |  gpe & gqd & gqf  ;
 QRA <= IRA ; 
 QSA <= ISA ; 
 QTA <= ITA ; 
 bbc <= idc ; 
 bbd <= idd ; 
 BCC <= BBC ; 
 BCD <= BBD ; 
 ODC <=  IDC & TTE  |  BEC & TGE  ; 
 OEC <=  IDC & TTE  |  BEC & TGE  ; 
 OHJ <=  GRJ & grc & grf  |  grj & GRC & grf  |  grj & grc & GRF  |  GRJ & GRC & GRF  ;
 oij <=  GRJ & grc & grf  |  grj & GRC & grf  |  grj & grc & GRF  |  grj & grc & grf  ;
 BDC <= BCC ; 
 BDD <= BCD ; 
 BEC <= BDC ; 
 BED <= BDD ; 
 OAD <=  ICD & TSF  |  BAD & TKF  |  AAD & THF  ; 
 AAC <=  ICC & TSB  |  BAC & TKB  |  AAC & THB  ; 
 OAC <=  ICC & TSE  |  BAC & TKE  |  AAC & THE  ; 
 OBC <=  ICC & TSE  |  BAC & TKE  |  AAC & THE  ; 
 KGA <=  JGB & jga & jfa  |  jgb & JGA & jfa  |  jgb & jga & JFA  |  JGB & JGA & JFA  ;
 kha <=  JGB & jga & jfa  |  jgb & JGA & jfa  |  jgb & jga & JFA  |  jgb & jga & jfa  ;
 KIA <=  JIA & jha & jib  |  jia & JHA & jib  |  jia & jha & JIB  |  JIA & JHA & JIB  ;
 kja <=  JIA & jha & jib  |  jia & JHA & jib  |  jia & jha & JIB  |  jia & jha & jib  ;
 oqj <=  MIA & mha & nha  |  mia & MHA & nha  |  mia & mha & NHA  |  mia & mha & nha  ;
 KIC <=  JHC & jhb & jie  |  jhc & JHB & jie  |  jhc & jhb & JIE  |  JHC & JHB & JIE  ;
 kjc <=  JHC & jhb & jie  |  jhc & JHB & jie  |  jhc & jhb & JIE  |  jhc & jhb & jie  ;
 KCA <=  JBA & jca & jcb  |  jba & JCA & jcb  |  jba & jca & JCB  |  JBA & JCA & JCB  ;
 kda <=  JBA & jca & jcb  |  jba & JCA & jcb  |  jba & jca & JCB  |  jba & jca & jcb  ;
 KCB <= HCA ; 
 KGC <=  HGG & jfc & jfb  |  hgg & JFC & jfb  |  hgg & jfc & JFB  |  HGG & JFC & JFB  ;
 khc <=  HGG & jfc & jfb  |  hgg & JFC & jfb  |  hgg & jfc & JFB  |  hgg & jfc & jfb  ;
 MGB <= KGA ; 
 MIA <=  LIA & lib & lha  |  lia & LIB & lha  |  lia & lib & LHA  |  LIA & LIB & LHA  ;
 mja <=  LIA & lib & lha  |  lia & LIB & lha  |  lia & lib & LHA  |  lia & lib & lha  ;
 KKA <=  JKA & jja & jkb  |  jka & JJA & jkb  |  jka & jja & JKB  |  JKA & JJA & JKB  ;
 kla <=  JKA & jja & jkb  |  jka & JJA & jkb  |  jka & jja & JKB  |  jka & jja & jkb  ;
 KMA <=  JLA & jma & jmb  |  jla & JMA & jmb  |  jla & jma & JMB  |  JLA & JMA & JMB  ;
 kna <=  JLA & jma & jmb  |  jla & JMA & jmb  |  jla & jma & JMB  |  jla & jma & jmb  ;
 MQC <= KPA ; 
 KOA <=  JOA & jna & job  |  joa & JNA & job  |  joa & jna & JOB  |  JOA & JNA & JOB  ;
 kpa <=  JOA & jna & job  |  joa & JNA & job  |  joa & jna & JOB  |  joa & jna & job  ;
 MKA <=  KKA & kja & lja  |  kka & KJA & lja  |  kka & kja & LJA  |  KKA & KJA & LJA  ;
 mla <=  KKA & kja & lja  |  kka & KJA & lja  |  kka & kja & LJA  |  kka & kja & lja  ;
 HMG <=  GLE & gme & gmb  |  gle & GME & gmb  |  gle & gme & GMB  |  GLE & GME & GMB  ;
 hng <=  GLE & gme & gmb  |  gle & GME & gmb  |  gle & gme & GMB  |  gle & gme & gmb  ;
 KKC <=  JJB & jje & hkg  |  jjb & JJE & hkg  |  jjb & jje & HKG  |  JJB & JJE & HKG  ;
 klc <=  JJB & jje & hkg  |  jjb & JJE & hkg  |  jjb & jje & HKG  |  jjb & jje & hkg  ;
 KKE <= JJC ; 
 KMC <=  JLB & jlc & hlc  |  jlb & JLC & hlc  |  jlb & jlc & HLC  |  JLB & JLC & HLC  ;
 knc <=  JLB & jlc & hlc  |  jlb & JLC & hlc  |  jlb & jlc & HLC  |  jlb & jlc & hlc  ;
 MMC <= LMA ; 
 KOC <=  HOC & hnc & jnb  |  hoc & HNC & jnb  |  hoc & hnc & JNB  |  HOC & HNC & JNB  ;
 kpc <=  HOC & hnc & jnb  |  hoc & HNC & jnb  |  hoc & hnc & JNB  |  hoc & hnc & jnb  ;
 MOC <= LNA ; 
 OPK <=  MKA & mja & mkb  |  mka & MJA & mkb  |  mka & mja & MKB  |  MKA & MJA & MKB  ;
 oqk <=  MKA & mja & mkb  |  mka & MJA & mkb  |  mka & mja & MKB  |  mka & mja & mkb  ;
 OPM <=  MLA & nma & mlb  |  mla & NMA & mlb  |  mla & nma & MLB  |  MLA & NMA & MLB  ;
 oqm <=  MLA & nma & mlb  |  mla & NMA & mlb  |  mla & nma & MLB  |  mla & nma & mlb  ;
 MOA <=  KNC & lnb & lob  |  knc & LNB & lob  |  knc & lnb & LOB  |  KNC & LNB & LOB  ;
 mpa <=  KNC & lnb & lob  |  knc & LNB & lob  |  knc & lnb & LOB  |  knc & lnb & lob  ;
 MOB <= LOA ; 
 THA <= QHA ; 
 THC <= QHA ; 
 THE <= QHA ; 
 AAE <=  ICE & TSA  |  BAE & TKA  |  AAE & THA  ; 
 AAF <=  ICF & TSA  |  BAF & TKA  |  AAF & THA  ; 
 OAE <=  ICE & TSC  |  BAE & TKC  |  AAE & THC  ; 
 OBE <=  ICE & TSC  |  BAE & TKC  |  AAE & THC  ; 
 HOG <=  GNE & gof & goc  |  gne & GOF & goc  |  gne & gof & GOC  |  GNE & GOF & GOC  ;
 hpg <=  GNE & gof & goc  |  gne & GOF & goc  |  gne & gof & GOC  |  gne & gof & goc  ;
 HQG <=  GQE & gpf & gqb  |  gqe & GPF & gqb  |  gqe & gpf & GQB  |  GQE & GPF & GQB  ;
 ohg <=  GQE & gpf & gqb  |  gqe & GPF & gqb  |  gqe & gpf & GQB  |  gqe & gpf & gqb  ;
 BDE <= BCE ; 
 BDF <= BCF ; 
 BEE <= BDE ; 
 BEF <= BDF ; 
 OAF <=  ICF & TSD  |  BAF & TKD  |  AAF & THD  ; 
 OBF <=  ICF & TSD  |  BAF & TKD  |  AAF & THD  ; 
 bbe <= ide ; 
 bbf <= idf ; 
 BCE <= BBE ; 
 BCF <= BBF ; 
 ODE <=  IDE & TTC  |  BEE & TGC  ; 
 OEE <=  IDE & TTC  |  BEE & TGC  ; 
 KQC <=  JQE & jpb & jpc  |  jqe & JPB & jpc  |  jqe & jpb & JPC  |  JQE & JPB & JPC  ;
 okc <=  JQE & jpb & jpc  |  jqe & JPB & jpc  |  jqe & jpb & JPC  |  jqe & jpb & jpc  ;
 OKF <= JRE ; 
 TTA <= QTA ; 
 TTC <= QTA ; 
 TTE <= QTA ; 
 BAE <=  IDE & TTA  |  BEE & TGA  ; 
 BAF <=  IDF & TTA  |  BEF & TGA  ; 
 ODF <=  IDF & TTD  |  BEF & TGD  ; 
 OEF <=  IDF & TTD  |  BEF & TGD  ; 
 OCH <=  ICH & TSF  |  BAH & TKF  |  AAH & THF  ; 
 ttb <= qta ; 
 ttd <= qta ; 
 ttf <= qta ; 
 BAG <=  IDG & TTB  |  BEG & TGB  ; 
 BAH <=  IDH & TTB  |  BEH & TGB  ; 
 ODH <=  IDH & TTF  |  BEH & TGF  ; 
 OEH <=  IDH & TTF  |  BEH & TGF  ; 
 OFH <=  IDH & TTF  |  BEH & TGF  ; 
 OMB <=  LRA & lrb  |  lra & LRB  ; 
 bbg <= idg ; 
 bbh <= idh ; 
 BCG <= BBG ; 
 BCH <= BBH ; 
 ODG <=  IDG & TTE  |  BEG & TGE  ; 
 OEG <=  IDG & TTE  |  BEG & TGE  ; 
 OFG <=  IDG & TTE  |  BEG & TGE  ; 
 OKD <=  JRB & jrc & jrd  |  jrb & JRC & jrd  |  jrb & jrc & JRD  |  JRB & JRC & JRD  ;
 old <=  JRB & jrc & jrd  |  jrb & JRC & jrd  |  jrb & jrc & JRD  |  jrb & jrc & jrd  ;
 BDG <= BCG ; 
 BDH <= BCH ; 
 BEG <= BDG ; 
 BEH <= BDH ; 
 OAH <=  ICH & TSF  |  BAH & TKF  |  AAH & THF  ; 
 OBH <=  ICH & TSF  |  BAH & TKF  |  AAH & THF  ; 
 thb <= qha ; 
 thd <= qha ; 
 thf <= qha ; 
 AAG <=  ICG & TSB  |  BAG & TKB  |  AAG & THB  ; 
 AAH <=  ICH & TSB  |  BAH & TKB  |  AAH & THB  ; 
 OAG <=  ICG & TSE  |  BAG & TKE  |  AAG & THE  ; 
 OBG <=  ICG & TSE  |  BAG & TKE  |  AAG & THE  ; 
 OCG <=  ICG & TSE  |  BAG & TKE  |  AAG & THE  ; 
 OPQ <=  NQA & npa & mpa  |  nqa & NPA & mpa  |  nqa & npa & MPA  |  NQA & NPA & MPA  ;
 oqq <=  NQA & npa & mpa  |  nqa & NPA & mpa  |  nqa & npa & MPA  |  nqa & npa & mpa  ;
 OPR <= NRA ; 
 KEA <=  JEA & jeb & jda  |  jea & JEB & jda  |  jea & jeb & JDA  |  JEA & JEB & JDA  ;
 kfa <=  JEA & jeb & jda  |  jea & JEB & jda  |  jea & jeb & JDA  |  jea & jeb & jda  ;
 mfa <=  LEA & lda  |  lea & LDA  |  lea & lda  ; 
 MGA <=  LFA & lga & kfa  |  lfa & LGA & kfa  |  lfa & lga & KFA  |  LFA & LGA & KFA  ;
 mha <=  LFA & lga & kfa  |  lfa & LGA & kfa  |  lfa & lga & KFA  |  lfa & lga & kfa  ;
 KEB <=  JDB & jed & jec  |  jdb & JED & jec  |  jdb & jed & JEC  |  JDB & JED & JEC  ;
 kfb <=  JDB & jed & jec  |  jdb & JED & jec  |  jdb & jed & JEC  |  jdb & jed & jec  ;
 KGB <=  JGC & jgd & jfd  |  jgc & JGD & jfd  |  jgc & jgd & JFD  |  JGC & JGD & JFD  ;
 khb <=  JGC & jgd & jfd  |  jgc & JGD & jfd  |  jgc & jgd & JFD  |  jgc & jgd & jfd  ;
 KIB <=  JID & jhd & jic  |  jid & JHD & jic  |  jid & jhd & JIC  |  JID & JHD & JIC  ;
 kjb <=  JID & jhd & jic  |  jid & JHD & jic  |  jid & jhd & JIC  |  jid & jhd & jic  ;
 onb <=  LRA & lrb  |  lra & LRB  |  lra & lrb  ; 
 MQA <=  LPA & lqa & lpb  |  lpa & LQA & lpb  |  lpa & lqa & LPB  |  LPA & LQA & LPB  ;
 oma <=  LPA & lqa & lpb  |  lpa & LQA & lpb  |  lpa & lqa & LPB  |  lpa & lqa & lpb  ;
 MQB <= LQB ; 
 MMA <=  LLA & llb & lmb  |  lla & LLB & lmb  |  lla & llb & LMB  |  LLA & LLB & LMB  ;
 mna <=  LLA & llb & lmb  |  lla & LLB & lmb  |  lla & llb & LMB  |  lla & llb & lmb  ;
 MMB <= KLC ; 
 OPO <=  NOA & nna & mna  |  noa & NNA & mna  |  noa & nna & MNA  |  NOA & NNA & MNA  ;
 oqo <=  NOA & nna & mna  |  noa & NNA & mna  |  noa & nna & MNA  |  noa & nna & mna  ;
 MKB <=  LKA & lkb & ljb  |  lka & LKB & ljb  |  lka & lkb & LJB  |  LKA & LKB & LJB  ;
 mlb <=  LKA & lkb & ljb  |  lka & LKB & ljb  |  lka & lkb & LJB  |  lka & lkb & ljb  ;
 KKB <=  JKC & jjd & jkd  |  jkc & JJD & jkd  |  jkc & jjd & JKD  |  JKC & JJD & JKD  ;
 klb <=  JKC & jjd & jkd  |  jkc & JJD & jkd  |  jkc & jjd & JKD  |  jkc & jjd & jkd  ;
 KKD <= HJF ; 
 KMB <=  JLD & jmd & jmc  |  jld & JMD & jmc  |  jld & jmd & JMC  |  JLD & JMD & JMC  ;
 knb <=  JLD & jmd & jmc  |  jld & JMD & jmc  |  jld & jmd & JMC  |  jld & jmd & jmc  ;
 KMD <= HLF ; 
 KOB <=  JOC & jod & jnd  |  joc & JOD & jnd  |  joc & jod & JND  |  JOC & JOD & JND  ;
 kpb <=  JOC & jod & jnd  |  joc & JOD & jnd  |  joc & jod & JND  |  joc & jod & jnd  ;
 KOD <= JNC ; 
 TSA <= QSA ; 
 TSC <= QSA ; 
 TSE <= QSA ; 
 AAI <=  ICI & TSA  |  BAI & TKA  |  AAI & THA  ; 
 AAJ <=  ICJ & TSA  |  BAJ & TKA  |  AAJ & THA  ; 
 OAI <=  ICI & TSC  |  BAI & TKC  |  AAI & THC  ; 
 OBI <=  ICI & TSC  |  BAI & TKC  |  AAI & THC  ; 
 OCI <=  ICI & TSC  |  BAI & TKC  |  AAI & THC  ; 
 BDI <= BCI ; 
 BDJ <= BCJ ; 
 BEI <= BDI ; 
 BEJ <= BDJ ; 
 OAJ <=  ICJ & TSD  |  BAJ & TKD  |  AAJ & THD  ; 
 OBJ <=  ICJ & TSD  |  BAJ & TKD  |  AAJ & THD  ; 
 OCJ <=  ICJ & TSD  |  BAJ & TKD  |  AAJ & THD  ; 
 KQA <=  JPA & jqa & jqb  |  jpa & JQA & jqb  |  jpa & jqa & JQB  |  JPA & JQA & JQB  ;
 oka <=  JPA & jqa & jqb  |  jpa & JQA & jqb  |  jpa & jqa & JQB  |  jpa & jqa & jqb  ;
 OKE <= JRA ; 
 bbi <= idi ; 
 bbj <= idj ; 
 BCI <= BBI ; 
 BCJ <= BBJ ; 
 ODI <=  IDI & TTC  |  BEI & TGC  ; 
 OEI <=  IDI & TTC  |  BEI & TGC  ; 
 OFI <=  IDI & TTC  |  BEI & TGC  ; 
 BCK <= BBK ; 
 TGA <= QGA ; 
 TGC <= QGA ; 
 TGE <= QGA ; 
 BAI <=  IDI & TTA  |  BEI & TGA  ; 
 BAJ <=  IDJ & TTA  |  BEJ & TGA  ; 
 ODJ <=  IDJ & TTD  |  BEJ & TGD  ; 
 OEJ <=  IDJ & TTD  |  BEJ & TGD  ; 
 OFJ <=  IDJ & TTD  |  BEJ & TGD  ; 
 OBL <=  ICL & TSF  |  BAL & TKF  |  AAL & THF  ; 
 tgb <= qga ; 
 tgd <= qga ; 
 tgf <= qga ; 
 BAK <=  IDK & TTB  |  BEK & TGB  ; 
 BAL <=  IDL & TTB  |  BEL & TGB  ; 
 ODL <=  IDL & TTF  |  BEL & TGF  ; 
 OEL <=  IDL & TTF  |  BEL & TGF  ; 
 OFL <=  IDL & TTF  |  BEL & TGF  ; 
 KQB <=  JPD & jqd & jqc  |  jpd & JQD & jqc  |  jpd & jqd & JQC  |  JPD & JQD & JQC  ;
 okb <=  JPD & jqd & jqc  |  jpd & JQD & jqc  |  jpd & jqd & JQC  |  jpd & jqd & jqc  ;
 KQD <= HPF ; 
 bbk <= idk ; 
 bbl <= idl ; 
 BCL <= BBL ; 
 ODK <=  IDK & TTE  |  BEK & TGE  ; 
 OEK <=  IDK & TTE  |  BEK & TGE  ; 
 OFK <=  IDK & TTE  |  BEK & TGE  ; 
 BDK <= BCK ; 
 BDL <= BCL ; 
 BEK <= BDK ; 
 BEL <= BDL ; 
 OAL <=  ICL & TSF  |  BAL & TKF  |  AAL & THF  ; 
 OCL <=  ICL & TSF  |  BAL & TKF  |  AAL & THF  ; 
 tsb <= qsa ; 
 tsd <= qsa ; 
 tsf <= qsa ; 
 AAK <=  ICK & TSB  |  BAK & TKB  |  AAK & THB  ; 
 AAL <=  ICL & TSB  |  BAL & TKB  |  AAL & THB  ; 
 OAK <=  ICK & TSE  |  BAK & TKE  |  AAK & THE  ; 
 OBK <=  ICK & TSE  |  BAK & TKE  |  AAK & THE  ; 
 OCK <=  ICK & TSE  |  BAK & TKE  |  AAK & THE  ; 
 HCA <=  GCG & gbd & gba  |  gcg & GBD & gba  |  gcg & gbd & GBA  |  GCG & GBD & GBA  ;
 hda <=  GCG & gbd & gba  |  gcg & GBD & gba  |  gcg & gbd & GBA  |  gcg & gbd & gba  ;
 HEA <=  GDG & geh & gda  |  gdg & GEH & gda  |  gdg & geh & GDA  |  GDG & GEH & GDA  ;
 hfa <=  GDG & geh & gda  |  gdg & GEH & gda  |  gdg & geh & GDA  |  gdg & geh & gda  ;
 HGA <=  GFH & ggg & gfe  |  gfh & GGG & gfe  |  gfh & ggg & GFE  |  GFH & GGG & GFE  ;
 hha <=  GFH & ggg & gfe  |  gfh & GGG & gfe  |  gfh & ggg & GFE  |  gfh & ggg & gfe  ;
 HIA <=  GIH & ghg & gha  |  gih & GHG & gha  |  gih & ghg & GHA  |  GIH & GHG & GHA  ;
 hja <=  GIH & ghg & gha  |  gih & GHG & gha  |  gih & ghg & GHA  |  gih & ghg & gha  ;
 HEC <=  GEG & gei & gdh  |  geg & GEI & gdh  |  geg & gei & GDH  |  GEG & GEI & GDH  ;
 hfc <=  GEG & gei & gdh  |  geg & GEI & gdh  |  geg & gei & GDH  |  geg & gei & gdh  ;
 HGC <=  GFG & ggf & ggh  |  gfg & GGF & ggh  |  gfg & ggf & GGH  |  GFG & GGF & GGH  ;
 hhc <=  GFG & ggf & ggh  |  gfg & GGF & ggh  |  gfg & ggf & GGH  |  gfg & ggf & ggh  ;
 HIC <=  GII & gig & ghf  |  gii & GIG & ghf  |  gii & gig & GHF  |  GII & GIG & GHF  ;
 hjc <=  GII & gig & ghf  |  gii & GIG & ghf  |  gii & gig & GHF  |  gii & gig & ghf  ;
 HIG <= FIA ; 
 HCD <=  GBC & gcc & gce  |  gbc & GCC & gce  |  gbc & gcc & GCE  |  GBC & GCC & GCE  ;
 hdd <=  GBC & gcc & gce  |  gbc & GCC & gce  |  gbc & gcc & GCE  |  gbc & gcc & gce  ;
 HEG <= GDF ; 
 HGG <=  GFI & gfd & ggc  |  gfi & GFD & ggc  |  gfi & gfd & GGC  |  GFI & GFD & GGC  ;
 hhg <=  GFI & gfd & ggc  |  gfi & GFD & ggc  |  gfi & gfd & GGC  |  gfi & gfd & ggc  ;
 HAA <=  FAE & gad & gaa  |  fae & GAD & gaa  |  fae & gad & GAA  |  FAE & GAD & GAA  ;
 hba <=  FAE & gad & gaa  |  fae & GAD & gaa  |  fae & gad & GAA  |  fae & gad & gaa  ;
 HCE <=  GCI & gbb & gcb  |  gci & GBB & gcb  |  gci & gbb & GCB  |  GCI & GBB & GCB  ;
 hde <=  GCI & gbb & gcb  |  gci & GBB & gcb  |  gci & gbb & GCB  |  gci & gbb & gcb  ;
 HEE <=  GEA & gde & gej  |  gea & GDE & gej  |  gea & gde & GEJ  |  GEA & GDE & GEJ  ;
 hfe <=  GEA & gde & gej  |  gea & GDE & gej  |  gea & gde & GEJ  |  gea & gde & gej  ;
 HIE <=  GIJ & gia & ghe  |  gij & GIA & ghe  |  gij & gia & GHE  |  GIJ & GIA & GHE  ;
 hje <=  GIJ & gia & ghe  |  gij & GIA & ghe  |  gij & gia & GHE  |  gij & gia & ghe  ;
 HGE <=  FGA & fgf & ggi  |  fga & FGF & ggi  |  fga & fgf & GGI  |  FGA & FGF & GGI  ;
 hhe <=  FGA & fgf & ggi  |  fga & FGF & ggi  |  fga & fgf & GGI  |  fga & fgf & ggi  ;
 HEF <=  GDB & gdi & gec  |  gdb & GDI & gec  |  gdb & gdi & GEC  |  GDB & GDI & GEC  ;
 hff <=  GDB & gdi & gec  |  gdb & GDI & gec  |  gdb & gdi & GEC  |  gdb & gdi & gec  ;
 HGF <=  GFJ & gfc & ggb  |  gfj & GFC & ggb  |  gfj & gfc & GGB  |  GFJ & GFC & GGB  ;
 hhf <=  GFJ & gfc & ggb  |  gfj & GFC & ggb  |  gfj & gfc & GGB  |  gfj & gfc & ggb  ;
 HIF <=  GHI & ghb & gic  |  ghi & GHB & gic  |  ghi & ghb & GIC  |  GHI & GHB & GIC  ;
 hjf <=  GHI & ghb & gic  |  ghi & GHB & gic  |  ghi & ghb & GIC  |  ghi & ghb & gic  ;
 HKA <=  GJH & gkh & gjb  |  gjh & GKH & gjb  |  gjh & gkh & GJB  |  GJH & GKH & GJB  ;
 hla <=  GJH & gkh & gjb  |  gjh & GKH & gjb  |  gjh & gkh & GJB  |  gjh & gkh & gjb  ;
 HMA <=  GLH & gmh & glb  |  glh & GMH & glb  |  glh & gmh & GLB  |  GLH & GMH & GLB  ;
 hna <=  GLH & gmh & glb  |  glh & GMH & glb  |  glh & gmh & GLB  |  glh & gmh & glb  ;
 HOA <=  GOI & gnh & gnb  |  goi & GNH & gnb  |  goi & gnh & GNB  |  GOI & GNH & GNB  ;
 hpa <=  GOI & gnh & gnb  |  goi & GNH & gnb  |  goi & gnh & GNB  |  goi & gnh & gnb  ;
 HKC <=  GKI & gjg & gkg  |  gki & GJG & gkg  |  gki & gjg & GKG  |  GKI & GJG & GKG  ;
 hlc <=  GKI & gjg & gkg  |  gki & GJG & gkg  |  gki & gjg & GKG  |  gki & gjg & gkg  ;
 HMC <=  GMI & gla & gmd  |  gmi & GLA & gmd  |  gmi & gla & GMD  |  GMI & GLA & GMD  ;
 hnc <=  GMI & gla & gmd  |  gmi & GLA & gmd  |  gmi & gla & GMD  |  gmi & gla & gmd  ;
 HOC <=  GOJ & gna & gob  |  goj & GNA & gob  |  goj & gna & GOB  |  GOJ & GNA & GOB  ;
 hpc <=  GOJ & gna & gob  |  goj & GNA & gob  |  goj & gna & GOB  |  goj & gna & gob  ;
 HOE <=  GOK & gnf & goa  |  gok & GNF & goa  |  gok & gnf & GOA  |  GOK & GNF & GOA  ;
 hpe <=  GOK & gnf & goa  |  gok & GNF & goa  |  gok & gnf & GOA  |  gok & gnf & goa  ;
 HKE <=  GKJ & gjf & fkb  |  gkj & GJF & fkb  |  gkj & gjf & FKB  |  GKJ & GJF & FKB  ;
 hle <=  GKJ & gjf & fkb  |  gkj & GJF & fkb  |  gkj & gjf & FKB  |  gkj & gjf & fkb  ;
 HKH <= FKA ; 
 HME <=  GLF & gmj & fma  |  glf & GMJ & fma  |  glf & gmj & FMA  |  GLF & GMJ & FMA  ;
 hne <=  GLF & gmj & fma  |  glf & GMJ & fma  |  glf & gmj & FMA  |  glf & gmj & fma  ;
 HKF <=  GJJ & gjc & gkc  |  gjj & GJC & gkc  |  gjj & gjc & GKC  |  GJJ & GJC & GKC  ;
 hlf <=  GJJ & gjc & gkc  |  gjj & GJC & gkc  |  gjj & gjc & GKC  |  gjj & gjc & gkc  ;
 HMF <=  GLC & glj & gmc  |  glc & GLJ & gmc  |  glc & glj & GMC  |  GLC & GLJ & GMC  ;
 hnf <=  GLC & glj & gmc  |  glc & GLJ & gmc  |  glc & glj & GMC  |  glc & glj & gmc  ;
 HOF <=  GNC & god & gnj  |  gnc & GOD & gnj  |  gnc & god & GNJ  |  GNC & GOD & GNJ  ;
 hpf <=  GNC & god & gnj  |  gnc & GOD & gnj  |  gnc & god & GNJ  |  gnc & god & gnj  ;
 HQA <=  GQH & gpi & gpc  |  gqh & GPI & gpc  |  gqh & gpi & GPC  |  GQH & GPI & GPC  ;
 oha <=  GQH & gpi & gpc  |  gqh & GPI & gpc  |  gqh & gpi & GPC  |  gqh & gpi & gpc  ;
 TKA <= QKA ; 
 TKE <= QKA ; 
 AAM <=  ICM & TSA  |  BAM & TKA  |  AAM & THA  ; 
 AAN <=  ICN & TSA  |  BAN & TKA  |  AAN & THA  ; 
 OAM <=  ICM & TSC  |  BAM & TKC  |  AAM & THC  ; 
 OBM <=  ICM & TSC  |  BAM & TKC  |  AAM & THC  ; 
 OCM <=  ICM & TSC  |  BAM & TKC  |  AAM & THC  ; 
 BDM <= BCM ; 
 BDN <= BCN ; 
 BEM <= BDM ; 
 BEN <= BDN ; 
 OAN <=  ICN & TSD  |  BAN & TKD  |  AAN & THD  ; 
 OBN <=  ICN & TSD  |  BAN & TKD  |  AAN & THD  ; 
 OCN <=  ICN & TSD  |  BAN & TKD  |  AAN & THD  ; 
 OCP <=  ICP & TSF  |  BAP & TKF  |  AAP & THF  ; 
 bbm <= idm ; 
 bbn <= idn ; 
 BCM <= BBM ; 
 BCN <= BBN ; 
 ODM <=  IDM & TTC  |  BEM & TGC  ; 
 OEM <=  IDM & TTC  |  BEM & TGC  ; 
 OFM <=  IDM & TTC  |  BEM & TGC  ; 
 BCO <= BBO ; 
 bbp <= idp ; 
 HQC <=  GQI & gpb & gqa  |  gqi & GPB & gqa  |  gqi & gpb & GQA  |  GQI & GPB & GQA  ;
 ohc <=  GQI & gpb & gqa  |  gqi & GPB & gqa  |  gqi & gpb & GQA  |  gqi & gpb & gqa  ;
 HQH <= FPB ; 
 BAM <=  IDM & TTA  |  BEM & TGA  ; 
 BAN <=  IDN & TTA  |  BEN & TGA  ; 
 ODN <=  IDN & TTD  |  BEN & TGD  ; 
 OEN <=  IDN & TTD  |  BEN & TGD  ; 
 OFN <=  IDN & TTD  |  BEN & TGD  ; 
 BAO <=  IDO & TTB  |  BEO & TGB  ; 
 BAP <=  IDP & TTB  |  BEP & TGB  ; 
 ODP <=  IDP & TTF  |  BEP & TGF  ; 
 OEP <=  IDP & TTF  |  BEP & TGF  ; 
 OFP <=  IDP & TTF  |  BEP & TGF  ; 
 bbo <= ido ; 
 BCP <= BBP ; 
 ODO <=  IDO & TTE  |  BEO & TGE  ; 
 OEO <=  IDO & TTE  |  BEO & TGE  ; 
 OFO <=  IDO & TTE  |  BEO & TGE  ; 
 HQE <=  GQJ & gpg & gpa  |  gqj & GPG & gpa  |  gqj & gpg & GPA  |  GQJ & GPG & GPA  ;
 ohe <=  GQJ & gpg & gpa  |  gqj & GPG & gpa  |  gqj & gpg & GPA  |  gqj & gpg & gpa  ;
 HQI <= FQA ; 
 BDO <= BCO ; 
 BDP <= BCP ; 
 BEO <= BDO ; 
 BEP <= BDP ; 
 OAP <=  ICP & TSF  |  BAP & TKF  |  AAP & THF  ; 
 OBP <=  ICP & TSF  |  BAP & TKF  |  AAP & THF  ; 
 HQF <=  GPD & gqc & gpk  |  gpd & GQC & gpk  |  gpd & gqc & GPK  |  GPD & GQC & GPK  ;
 ohf <=  GPD & gqc & gpk  |  gpd & GQC & gpk  |  gpd & gqc & GPK  |  gpd & gqc & gpk  ;
 tkb <= qka ; 
 TKC <= QKA ; 
 tkd <= qka ; 
 tkf <= qka ; 
 AAO <=  ICO & TSB  |  BAO & TKB  |  AAO & THB  ; 
 AAP <=  ICP & TSB  |  BAP & TKB  |  AAP & THB  ; 
 OAO <=  ICO & TSE  |  BAO & TKE  |  AAO & THE  ; 
 OBO <=  ICO & TSE  |  BAO & TKE  |  AAO & THE  ; 
 OCO <=  ICO & TSE  |  BAO & TKE  |  AAO & THE  ; 
 FAF <=  EAO & eap & eaq  |  eao & EAP & eaq  |  eao & eap & EAQ  |  EAO & EAP & EAQ  ;
 fbf <=  EAO & eap & eaq  |  eao & EAP & eaq  |  eao & eap & EAQ  |  eao & eap & eaq  ;
 FCG <=  ECP & ecq & ecr  |  ecp & ECQ & ecr  |  ecp & ecq & ECR  |  ECP & ECQ & ECR  ;
 fdg <=  ECP & ecq & ecr  |  ecp & ECQ & ecr  |  ecp & ecq & ECR  |  ecp & ecq & ecr  ;
 FCA <= QAB ; 
 FEH <=  EEQ & eer & ees  |  eeq & EER & ees  |  eeq & eer & EES  |  EEQ & EER & EES  ;
 ffh <=  EEQ & eer & ees  |  eeq & EER & ees  |  eeq & eer & EES  |  eeq & eer & ees  ;
 FGG <=  EGR & egs & egt  |  egr & EGS & egt  |  egr & egs & EGT  |  EGR & EGS & EGT  ;
 fhg <=  EGR & egs & egt  |  egr & EGS & egt  |  egr & egs & EGT  |  egr & egs & egt  ;
 FAE <=  EAL & eam & ean  |  eal & EAM & ean  |  eal & eam & EAN  |  EAL & EAM & EAN  ;
 fbe <=  EAL & eam & ean  |  eal & EAM & ean  |  eal & eam & EAN  |  eal & eam & ean  ;
 FCF <=  ECM & ecn & eco  |  ecm & ECN & eco  |  ecm & ecn & ECO  |  ECM & ECN & ECO  ;
 fdf <=  ECM & ecn & eco  |  ecm & ECN & eco  |  ecm & ecn & ECO  |  ecm & ecn & eco  ;
 FEB <= QAC ; 
 FEG <=  EEN & eeo & eep  |  een & EEO & eep  |  een & eeo & EEP  |  EEN & EEO & EEP  ;
 ffg <=  EEN & eeo & eep  |  een & EEO & eep  |  een & eeo & EEP  |  een & eeo & eep  ;
 FGF <=  EGO & egp & egq  |  ego & EGP & egq  |  ego & egp & EGQ  |  EGO & EGP & EGQ  ;
 fhf <=  EGO & egp & egq  |  ego & EGP & egq  |  ego & egp & EGQ  |  ego & egp & egq  ;
 FAD <=  EAI & eaj & eak  |  eai & EAJ & eak  |  eai & eaj & EAK  |  EAI & EAJ & EAK  ;
 fbd <=  EAI & eaj & eak  |  eai & EAJ & eak  |  eai & eaj & EAK  |  eai & eaj & eak  ;
 FCE <=  ECJ & eck & ecl  |  ecj & ECK & ecl  |  ecj & eck & ECL  |  ECJ & ECK & ECL  ;
 fde <=  ECJ & eck & ecl  |  ecj & ECK & ecl  |  ecj & eck & ECL  |  ecj & eck & ecl  ;
 FEF <=  EEK & eel & eem  |  eek & EEL & eem  |  eek & eel & EEM  |  EEK & EEL & EEM  ;
 fff <=  EEK & eel & eem  |  eek & EEL & eem  |  eek & eel & EEM  |  eek & eel & eem  ;
 FGE <=  EGL & egm & egn  |  egl & EGM & egn  |  egl & egm & EGN  |  EGL & EGM & EGN  ;
 fhe <=  EGL & egm & egn  |  egl & EGM & egn  |  egl & egm & EGN  |  egl & egm & egn  ;
 FAC <=  EAF & eag & eah  |  eaf & EAG & eah  |  eaf & eag & EAH  |  EAF & EAG & EAH  ;
 fbc <=  EAF & eag & eah  |  eaf & EAG & eah  |  eaf & eag & EAH  |  eaf & eag & eah  ;
 FCD <=  ECG & ech & eci  |  ecg & ECH & eci  |  ecg & ech & ECI  |  ECG & ECH & ECI  ;
 fdd <=  ECG & ech & eci  |  ecg & ECH & eci  |  ecg & ech & ECI  |  ecg & ech & eci  ;
 FEE <=  EEH & eei & eej  |  eeh & EEI & eej  |  eeh & eei & EEJ  |  EEH & EEI & EEJ  ;
 ffe <=  EEH & eei & eej  |  eeh & EEI & eej  |  eeh & eei & EEJ  |  eeh & eei & eej  ;
 FGD <=  EGI & egj & egk  |  egi & EGJ & egk  |  egi & egj & EGK  |  EGI & EGJ & EGK  ;
 fhd <=  EGI & egj & egk  |  egi & EGJ & egk  |  egi & egj & EGK  |  egi & egj & egk  ;
 OAA <=  ICA & TSC  |  BAA & TKC  |  AAA & THC  ; 
 CEI <= IEC & TRC |  AAI & trc ; 
 CEJ <= IED & TRC |  AAJ & trc ; 
 CEK <= IEE & TRC |  AAK & trc ; 
 FIH <=  EIS & eit & eiu  |  eis & EIT & eiu  |  eis & eit & EIU  |  EIS & EIT & EIU  ;
 fjh <=  EIS & eit & eiu  |  eis & EIT & eiu  |  eis & eit & EIU  |  eis & eit & eiu  ;
 AAA <=  ICA & TSA  |  BAA & TKA  |  AAA & THA  ; 
 dbb <= bab ; 
 dbc <= bac ; 
 dbd <= bad ; 
 dbe <= bae ; 
 FKI <=  EKT & eku & ekv  |  ekt & EKU & ekv  |  ekt & eku & EKV  |  EKT & EKU & EKV  ;
 fli <=  EKT & eku & ekv  |  ekt & EKU & ekv  |  ekt & eku & EKV  |  ekt & eku & ekv  ;
 DAF <= IBF ; 
 DAG <= IBG ; 
 CEL <= IEF & TRC |  AAL & trc ; 
 CEM <= IEG & TRC |  AAM & trc ; 
 CEN <= IEH & TRC |  AAN & trc ; 
 FIG <=  EIP & eiq & eir  |  eip & EIQ & eir  |  eip & eiq & EIR  |  EIP & EIQ & EIR  ;
 fjg <=  EIP & eiq & eir  |  eip & EIQ & eir  |  eip & eiq & EIR  |  eip & eiq & eir  ;
 DAN <= IBN ; 
 DAO <= IBO ; 
 DAP <= IBP ; 
 DBA <= BAA ; 
 FKH <=  EKQ & ekr & eks  |  ekq & EKR & eks  |  ekq & ekr & EKS  |  EKQ & EKR & EKS  ;
 flh <=  EKQ & ekr & eks  |  ekq & EKR & eks  |  ekq & ekr & EKS  |  ekq & ekr & eks  ;
 CEO <= IEI & TRC |  AAO & trc ; 
 CEP <= IEJ & TRC |  AAP & trc ; 
 CFA <= IEK & TRC |  IEK & trc ; 
 FIF <=  EIM & ein & eio  |  eim & EIN & eio  |  eim & ein & EIO  |  EIM & EIN & EIO  ;
 fjf <=  EIM & ein & eio  |  eim & EIN & eio  |  eim & ein & EIO  |  eim & ein & eio  ;
 DAM <= IBM ; 
 DAJ <= IBJ ; 
 DAL <= IBL ; 
 DAK <= IBK ; 
 FKG <=  EKN & eko & ekp  |  ekn & EKO & ekp  |  ekn & eko & EKP  |  EKN & EKO & EKP  ;
 flg <=  EKN & eko & ekp  |  ekn & EKO & ekp  |  ekn & eko & EKP  |  ekn & eko & ekp  ;
 trc <= qra ; 
 CFB <= IEL ; 
 CFC <= IEM ; 
 CFD <= IEN ; 
 FIE <=  EIJ & eik & eil  |  eij & EIK & eil  |  eij & eik & EIL  |  EIJ & EIK & EIL  ;
 fje <=  EIJ & eik & eil  |  eij & EIK & eil  |  eij & eik & EIL  |  eij & eik & eil  ;
 FQF <=  EQQ & eqr & eqs  |  eqq & EQR & eqs  |  eqq & eqr & EQS  |  EQQ & EQR & EQS  ;
 ogf <=  EQQ & eqr & eqs  |  eqq & EQR & eqs  |  eqq & eqr & EQS  |  eqq & eqr & eqs  ;
 DAH <= IBH ; 
 DAI <= IBI ; 
 FKF <=  EKK & ekl & ekm  |  ekk & EKL & ekm  |  ekk & ekl & EKM  |  EKK & EKL & EKM  ;
 flf <=  EKK & ekl & ekm  |  ekk & EKL & ekm  |  ekk & ekl & EKM  |  ekk & ekl & ekm  ;
 CBI <= IEC & TRB |  AAI & trb ; 
 CBJ <= IED & TRB |  AAJ & trb ; 
 CBK <= IEE & TRB |  AAK & trb ; 
 FMH <=  EMU & emv & emw  |  emu & EMV & emw  |  emu & emv & EMW  |  EMU & EMV & EMW  ;
 fnh <=  EMU & emv & emw  |  emu & EMV & emw  |  emu & emv & EMW  |  emu & emv & emw  ;
 FOI <=  EOV & eow & eox  |  eov & EOW & eox  |  eov & eow & EOX  |  EOV & EOW & EOX  ;
 fpi <=  EOV & eow & eox  |  eov & EOW & eox  |  eov & eow & EOX  |  eov & eow & eox  ;
 FQH <=  EQW & eqx & era  |  eqw & EQX & era  |  eqw & eqx & ERA  |  EQW & EQX & ERA  ;
 ogh <=  EQW & eqx & era  |  eqw & EQX & era  |  eqw & eqx & ERA  |  eqw & eqx & era  ;
 dbf <= baf ; 
 dbg <= bag ; 
 dbh <= bah ; 
 dbi <= bai ; 
 CBL <= IEF & TRB |  AAL & trb ; 
 CBM <= IEG & TRB |  AAM & trb ; 
 CBN <= IEH & TRB |  AAN & trb ; 
 FMG <=  EMR & ems & emt  |  emr & EMS & emt  |  emr & ems & EMT  |  EMR & EMS & EMT  ;
 fng <=  EMR & ems & emt  |  emr & EMS & emt  |  emr & ems & EMT  |  emr & ems & emt  ;
 FOH <=  EOS & eot & eou  |  eos & EOT & eou  |  eos & eot & EOU  |  EOS & EOT & EOU  ;
 fph <=  EOS & eot & eou  |  eos & EOT & eou  |  eos & eot & EOU  |  eos & eot & eou  ;
 FQG <=  EQT & equ & eqv  |  eqt & EQU & eqv  |  eqt & equ & EQV  |  EQT & EQU & EQV  ;
 ogg <=  EQT & equ & eqv  |  eqt & EQU & eqv  |  eqt & equ & EQV  |  eqt & equ & eqv  ;
 dhb <= bab ; 
 dhc <= bac ; 
 dhd <= bad ; 
 dhe <= bae ; 
 CBO <= IEI & TRB |  AAO & trb ; 
 CBP <= IEJ & TRB |  AAP & trb ; 
 CCA <= IEK & TRB |  IEK & trb ; 
 FMF <=  EMO & emp & emq  |  emo & EMP & emq  |  emo & emp & EMQ  |  EMO & EMP & EMQ  ;
 fnf <=  EMO & emp & emq  |  emo & EMP & emq  |  emo & emp & EMQ  |  emo & emp & emq  ;
 FOG <=  EOP & eoq & eor  |  eop & EOQ & eor  |  eop & eoq & EOR  |  EOP & EOQ & EOR  ;
 fpg <=  EOP & eoq & eor  |  eop & EOQ & eor  |  eop & eoq & EOR  |  eop & eoq & eor  ;
 TRB <= QRA ; 
 DGN <= IBN ; 
 DGO <= IBO ; 
 DGP <= IBP ; 
 DHA <= BAA ; 
 CCB <= IEL ; 
 CCC <= IEM ; 
 CCD <= IEN ; 
 FME <=  EML & emm & emn  |  eml & EMM & emn  |  eml & emm & EMN  |  EML & EMM & EMN  ;
 fne <=  EML & emm & emn  |  eml & EMM & emn  |  eml & emm & EMN  |  eml & emm & emn  ;
 FOF <=  EOM & eon & eoo  |  eom & EON & eoo  |  eom & eon & EOO  |  EOM & EON & EOO  ;
 fpf <=  EOM & eon & eoo  |  eom & EON & eoo  |  eom & eon & EOO  |  eom & eon & eoo  ;
 FQE <=  EQN & eqo & eqp  |  eqn & EQO & eqp  |  eqn & eqo & EQP  |  EQN & EQO & EQP  ;
 oge <=  EQN & eqo & eqp  |  eqn & EQO & eqp  |  eqn & eqo & EQP  |  eqn & eqo & eqp  ;
 DGK <= IBK ; 
 DGL <= IBL ; 
 DGM <= IBM ; 
 FAB <=  EAC & ead & eae  |  eac & EAD & eae  |  eac & ead & EAE  |  EAC & EAD & EAE  ;
 fbb <=  EAC & ead & eae  |  eac & EAD & eae  |  eac & ead & EAE  |  eac & ead & eae  ;
 FCC <=  ECD & ece & ecf  |  ecd & ECE & ecf  |  ecd & ece & ECF  |  ECD & ECE & ECF  ;
 fdc <=  ECD & ece & ecf  |  ecd & ECE & ecf  |  ecd & ece & ECF  |  ecd & ece & ecf  ;
 FED <=  EEE & eef & eeg  |  eee & EEF & eeg  |  eee & eef & EEG  |  EEE & EEF & EEG  ;
 ffd <=  EEE & eef & eeg  |  eee & EEF & eeg  |  eee & eef & EEG  |  eee & eef & eeg  ;
 FGC <=  EGF & egg & egh  |  egf & EGG & egh  |  egf & egg & EGH  |  EGF & EGG & EGH  ;
 fhc <=  EGF & egg & egh  |  egf & EGG & egh  |  egf & egg & EGH  |  egf & egg & egh  ;
 FAA <=  QAA & eaa & eab  |  qaa & EAA & eab  |  qaa & eaa & EAB  |  QAA & EAA & EAB  ;
 fba <=  QAA & eaa & eab  |  qaa & EAA & eab  |  qaa & eaa & EAB  |  qaa & eaa & eab  ;
 TAM <= QMM ; 
 TAR <= QMR ; 
 TAS <= QMS ; 
 FEC <=  EEB & eec & eed  |  eeb & EEC & eed  |  eeb & eec & EED  |  EEB & EEC & EED  ;
 ffc <=  EEB & eec & eed  |  eeb & EEC & eed  |  eeb & eec & EED  |  eeb & eec & eed  ;
 FGB <=  EGC & egd & ege  |  egc & EGD & ege  |  egc & egd & EGE  |  EGC & EGD & EGE  ;
 fhb <=  EGC & egd & ege  |  egc & EGD & ege  |  egc & egd & EGE  |  egc & egd & ege  ;
 FGA <=  QAD & ega & egb  |  qad & EGA & egb  |  qad & ega & EGB  |  QAD & EGA & EGB  ;
 fha <=  QAD & ega & egb  |  qad & EGA & egb  |  qad & ega & EGB  |  qad & ega & egb  ;
 FEA <= EEA ; 
 QAA <=  TAM  ; 
 QAB <=  TAR  |  TAS  ; 
 FCB <=  ECA & ecb & ecc  |  eca & ECB & ecc  |  eca & ecb & ECC  |  ECA & ECB & ECC  ;
 fdb <=  ECA & ecb & ecc  |  eca & ECB & ecc  |  eca & ecb & ECC  |  eca & ecb & ecc  ;
 FID <=  EIG & eih & eii  |  eig & EIH & eii  |  eig & eih & EII  |  EIG & EIH & EII  ;
 fjd <=  EIG & eih & eii  |  eig & EIH & eii  |  eig & eih & EII  |  eig & eih & eii  ;
 ddf <= ibf ; 
 ddg <= ibg ; 
 ddh <= ibh ; 
 ddi <= ibi ; 
 FKE <=  EKH & eki & ekj  |  ekh & EKI & ekj  |  ekh & eki & EKJ  |  EKH & EKI & EKJ  ;
 fle <=  EKH & eki & ekj  |  ekh & EKI & ekj  |  ekh & eki & EKJ  |  ekh & eki & ekj  ;
 CFE <= IEO ; 
 CFF <= IEP ; 
 CFG <= IEQ ; 
 FIC <=  EID & eie & eif  |  eid & EIE & eif  |  eid & eie & EIF  |  EID & EIE & EIF  ;
 fjc <=  EID & eie & eif  |  eid & EIE & eif  |  eid & eie & EIF  |  eid & eie & eif  ;
 DDB <= IBB ; 
 DDC <= IBC ; 
 DDD <= IBD ; 
 DDE <= IBE ; 
 FKD <=  EKE & ekf & ekg  |  eke & EKF & ekg  |  eke & ekf & EKG  |  EKE & EKF & EKG  ;
 fld <=  EKE & ekf & ekg  |  eke & EKF & ekg  |  eke & ekf & EKG  |  eke & ekf & ekg  ;
 FKB <= QAF ; 
 CFH <= IER ; 
 CFI <= IES ; 
 CFJ <= IET ; 
 FIB <=  EIA & eib & eic  |  eia & EIB & eic  |  eia & eib & EIC  |  EIA & EIB & EIC  ;
 fjb <=  EIA & eib & eic  |  eia & EIB & eic  |  eia & eib & EIC  |  eia & eib & eic  ;
 FIA <= QAE ; 
 DDA <= IBA ; 
 FKC <=  EKB & ekc & ekd  |  ekb & EKC & ekd  |  ekb & ekc & EKD  |  EKB & EKC & EKD  ;
 flc <=  EKB & ekc & ekd  |  ekb & EKC & ekd  |  ekb & ekc & EKD  |  ekb & ekc & ekd  ;
 CFK <= IEU ; 
 CFL <= IEV ; 
 CFM <= IEW ; 
 QAE <=  TAR  ; 
 QAF <=  TAM  |  TAR  ; 
 QAI <=  TAR  |  TAS  ; 
 FKA <= EKA ; 
 QAC <=  TAS  ; 
 QAD <=  TAM  ; 
 QAG <=  TAM  |  TAS  ; 
 QAH <=  TAR  ; 
 FMD <=  EMI & emj & emk  |  emi & EMJ & emk  |  emi & emj & EMK  |  EMI & EMJ & EMK  ;
 fnd <=  EMI & emj & emk  |  emi & EMJ & emk  |  emi & emj & EMK  |  emi & emj & emk  ;
 FOE <=  EOJ & eok & eol  |  eoj & EOK & eol  |  eoj & eok & EOL  |  EOJ & EOK & EOL  ;
 fpe <=  EOJ & eok & eol  |  eoj & EOK & eol  |  eoj & eok & EOL  |  eoj & eok & eol  ;
 FQD <=  EQK & eql & eqm  |  eqk & EQL & eqm  |  eqk & eql & EQM  |  EQK & EQL & EQM  ;
 ogd <=  EQK & eql & eqm  |  eqk & EQL & eqm  |  eqk & eql & EQM  |  eqk & eql & eqm  ;
 ddj <= ibj ; 
 ddk <= ibk ; 
 ddl <= ibl ; 
 ddm <= ibm ; 
 CCE <= IEO ; 
 CCF <= IEP ; 
 CCG <= IEQ ; 
 FMC <=  EMF & emg & emh  |  emf & EMG & emh  |  emf & emg & EMH  |  EMF & EMG & EMH  ;
 fnc <=  EMF & emg & emh  |  emf & EMG & emh  |  emf & emg & EMH  |  emf & emg & emh  ;
 FOD <=  EOG & eoh & eoi  |  eog & EOH & eoi  |  eog & eoh & EOI  |  EOG & EOH & EOI  ;
 fpd <=  EOG & eoh & eoi  |  eog & EOH & eoi  |  eog & eoh & EOI  |  eog & eoh & eoi  ;
 FQC <=  EQH & eqi & eqj  |  eqh & EQI & eqj  |  eqh & eqi & EQJ  |  EQH & EQI & EQJ  ;
 ogc <=  EQH & eqi & eqj  |  eqh & EQI & eqj  |  eqh & eqi & EQJ  |  eqh & eqi & eqj  ;
 dgf <= ibf ; 
 dgg <= ibg ; 
 dgh <= ibh ; 
 dgi <= ibi ; 
 CCH <= IER ; 
 CCI <= IES ; 
 CCJ <= IET ; 
 FMB <=  EMC & emd & eme  |  emc & EMD & eme  |  emc & emd & EME  |  EMC & EMD & EME  ;
 fnb <=  EMC & emd & eme  |  emc & EMD & eme  |  emc & emd & EME  |  emc & emd & eme  ;
 FOC <=  EOD & eoe & eof  |  eod & EOE & eof  |  eod & eoe & EOF  |  EOD & EOE & EOF  ;
 fpc <=  EOD & eoe & eof  |  eod & EOE & eof  |  eod & eoe & EOF  |  eod & eoe & eof  ;
 FQB <=  EQE & eqf & eqg  |  eqe & EQF & eqg  |  eqe & eqf & EQG  |  EQE & EQF & EQG  ;
 ogb <=  EQE & eqf & eqg  |  eqe & EQF & eqg  |  eqe & eqf & EQG  |  eqe & eqf & eqg  ;
 DGB <= IBB ; 
 DGC <= IBC ; 
 DGD <= IBD ; 
 DGE <= IBE ; 
 CCK <= IEU ; 
 CCL <= IEV ; 
 CCM <= IEW ; 
 FMA <=  QAG & ema & emb  |  qag & EMA & emb  |  qag & ema & EMB  |  QAG & EMA & EMB  ;
 fna <=  QAG & ema & emb  |  qag & EMA & emb  |  qag & ema & EMB  |  qag & ema & emb  ;
 FOB <=  EOA & eob & eoc  |  eoa & EOB & eoc  |  eoa & eob & EOC  |  EOA & EOB & EOC  ;
 fpb <=  EOA & eob & eoc  |  eoa & EOB & eoc  |  eoa & eob & EOC  |  eoa & eob & eoc  ;
 FOA <= QAH ; 
 FQA <=  EQB & eqc & eqd  |  eqb & EQC & eqd  |  eqb & eqc & EQD  |  EQB & EQC & EQD  ;
 oga <=  EQB & eqc & eqd  |  eqb & EQC & eqd  |  eqb & eqc & EQD  |  eqb & eqc & eqd  ;
 DGA <= IBA ; 
 QMM <= IMM ; 
 QMR <= IMR ; 
 QMS <= IMS ; 
 CCN <= IEX ; 
 CCO <= IEY ; 
 CCP <= IEZ ; 
end 
endmodule;
