module mb( IZZ,
 IBA, 
 IBB, 
 IBC, 
 IBD, 
 IBE, 
 IBF, 
 IBG, 
 IBH, 
 IBI, 
 IBJ, 
 IBK, 
 IBL, 
 IBM, 
 IBN, 
 IBO, 
 IBP, 
 ICA, 
 ICB, 
 ICC, 
 ICD, 
 ICE, 
 ICF, 
 ICG, 
 ICH, 
 ICI, 
 ICJ, 
 ICK, 
 ICL, 
 ICM, 
 ICN, 
 ICO, 
 ICP, 
 IDA, 
 IDB, 
 IDC, 
 IDD, 
 IDE, 
 IDF, 
 IDG, 
 IDH, 
 IDI, 
 IDJ, 
 IDK, 
 IDL, 
 IDM, 
 IDN, 
 IDO, 
 IDP, 
 IEA, 
 IEB, 
 IEC, 
 IED, 
 IEE, 
 IEF, 
 IEG, 
 IEH, 
 IEI, 
 IEJ, 
 IEK, 
 IEL, 
 IEM, 
 IEN, 
 IEO, 
 IEP, 
 IEQ, 
 IER, 
 IES, 
 IET, 
 IEU, 
 IEV, 
 IEW, 
 IEX, 
 IEY, 
 IEZ, 
 IFA, 
 IFB, 
 IFC, 
 IFD, 
 IFE, 
 IFFF , 
 IFG, 
 IFH, 
 IFI, 
 IFJ, 
 IFK, 
 IFL, 
 IFM, 
 IFN, 
 IFO, 
 IFP, 
 IGA, 
 IGB, 
 IGC, 
 IGD, 
 IGE, 
 IGF, 
 IGG, 
 IGH, 
 IGI, 
 IGJ, 
 IGK, 
 IGL, 
 IGM, 
 IGN, 
 IGO, 
 IGP, 
 IHA, 
 IIA, 
 IKA, 
 ILA, 
 ILB, 
 ILC, 
 ILD, 
 ILE, 
 ILF, 
 ILG, 
 ILH, 
 ILI, 
 ILJ, 
 ILK, 
 ILL, 
 ILM, 
 ILN, 
 ILO, 
 ILP, 
 IMA, 
 IMB, 
 IMC, 
 IMD, 
 IME, 
 IMF, 
 IMG, 
 IMH, 
 IMI, 
 IMJ, 
 IMK, 
 IML, 
 IMM, 
 IMN, 
 INA, 
 INB, 
 INC, 
 IND, 
 INE, 
 INF, 
 ING, 
 IOA, 
 IOB, 
 IOC, 
 IRA, 
 ISA, 
 ITA, 
 ITB, 
 OAA, 
 OAB, 
 OAC, 
 OAD, 
 OAE, 
 OAF, 
 OAG, 
 OAH, 
 OAI, 
 OAJ, 
 OAK, 
 OAL, 
 OAM, 
 OAN, 
 OAO, 
 OAP, 
 OBL, 
 OBM, 
 OBN, 
 OBO, 
 OBP, 
 OCA, 
 OCB, 
 OCC, 
 OCD, 
 OCE, 
 OCF, 
 OCG, 
 OCH, 
 OCI, 
 OCJ, 
 OCK, 
 OCL, 
 OCM, 
 OCN, 
 OCO, 
 OCP, 
 ODL, 
 ODM, 
 ODN, 
 ODO, 
 ODP, 
 OGA, 
 OGB, 
 OGC, 
 OGD, 
 OGE, 
 OGF, 
 OGG, 
 OGH, 
 OGI, 
 OGJ, 
 OGK, 
 OGL, 
 OGM, 
 OHA, 
 OHB, 
 OHC, 
 OHD, 
 OHE, 
 OHF, 
 OHG, 
 OHH, 
 OHI, 
 OHJ, 
 OKA, 
 OKB, 
 OKC, 
 OKD, 
 OKE, 
 OLD, 
 OMA, 
 OMB, 
 OPA, 
 OPB, 
 OPC, 
 OPD, 
 OPE, 
 OPF, 
 OPG, 
 OPH, 
 OPI, 
 OPK, 
 OPM, 
 OPO, 
 OPQ, 
 OPR, 
 OQA, 
 OQC, 
 OQE, 
 OQI, 
 OQK, 
 OQM, 
 OQO, 
OQQ ); 
    
 input IZZ; 
 input IBA; 
 input IBB; 
 input IBC; 
 input IBD; 
 input IBE; 
 input IBF; 
 input IBG; 
 input IBH; 
 input IBI; 
 input IBJ; 
 input IBK; 
 input IBL; 
 input IBM; 
 input IBN; 
 input IBO; 
 input IBP; 
 input ICA; 
 input ICB; 
 input ICC; 
 input ICD; 
 input ICE; 
 input ICF; 
 input ICG; 
 input ICH; 
 input ICI; 
 input ICJ; 
 input ICK; 
 input ICL; 
 input ICM; 
 input ICN; 
 input ICO; 
 input ICP; 
 input IDA; 
 input IDB; 
 input IDC; 
 input IDD; 
 input IDE; 
 input IDF; 
 input IDG; 
 input IDH; 
 input IDI; 
 input IDJ; 
 input IDK; 
 input IDL; 
 input IDM; 
 input IDN; 
 input IDO; 
 input IDP; 
 input IEA; 
 input IEB; 
 input IEC; 
 input IED; 
 input IEE; 
 input IEF; 
 input IEG; 
 input IEH; 
 input IEI; 
 input IEJ; 
 input IEK; 
 input IEL; 
 input IEM; 
 input IEN; 
 input IEO; 
 input IEP; 
 input IEQ; 
 input IER; 
 input IES; 
 input IET; 
 input IEU; 
 input IEV; 
 input IEW; 
 input IEX; 
 input IEY; 
 input IEZ; 
 input IFA; 
 input IFB; 
 input IFC; 
 input IFD; 
 input IFE; 
 input IFFF ; 
 input IFG; 
 input IFH; 
 input IFI; 
 input IFJ; 
 input IFK; 
 input IFL; 
 input IFM; 
 input IFN; 
 input IFO; 
 input IFP; 
 input IGA; 
 input IGB; 
 input IGC; 
 input IGD; 
 input IGE; 
 input IGF; 
 input IGG; 
 input IGH; 
 input IGI; 
 input IGJ; 
 input IGK; 
 input IGL; 
 input IGM; 
 input IGN; 
 input IGO; 
 input IGP; 
 input IHA; 
 input IIA; 
 input IKA; 
 input ILA; 
 input ILB; 
 input ILC; 
 input ILD; 
 input ILE; 
 input ILF; 
 input ILG; 
 input ILH; 
 input ILI; 
 input ILJ; 
 input ILK; 
 input ILL; 
 input ILM; 
 input ILN; 
 input ILO; 
 input ILP; 
 input IMA; 
 input IMB; 
 input IMC; 
 input IMD; 
 input IME; 
 input IMF; 
 input IMG; 
 input IMH; 
 input IMI; 
 input IMJ; 
 input IMK; 
 input IML; 
 input IMM; 
 input IMN; 
 input INA; 
 input INB; 
 input INC; 
 input IND; 
 input INE; 
 input INF; 
 input ING; 
 input IOA; 
 input IOB; 
 input IOC; 
 input IRA; 
 input ISA; 
 input ITA; 
 input ITB; 
 output OAA; 
 output OAB; 
 output OAC; 
 output OAD; 
 output OAE; 
 output OAF; 
 output OAG; 
 output OAH; 
 output OAI; 
 output OAJ; 
 output OAK; 
 output OAL; 
 output OAM; 
 output OAN; 
 output OAO; 
 output OAP; 
 output OBL; 
 output OBM; 
 output OBN; 
 output OBO; 
 output OBP; 
 output OCA; 
 output OCB; 
 output OCC; 
 output OCD; 
 output OCE; 
 output OCF; 
 output OCG; 
 output OCH; 
 output OCI; 
 output OCJ; 
 output OCK; 
 output OCL; 
 output OCM; 
 output OCN; 
 output OCO; 
 output OCP; 
 output ODL; 
 output ODM; 
 output ODN; 
 output ODO; 
 output ODP; 
 output OGA; 
 output OGB; 
 output OGC; 
 output OGD; 
 output OGE; 
 output OGF; 
 output OGG; 
 output OGH; 
 output OGI; 
 output OGJ; 
 output OGK; 
 output OGL; 
 output OGM; 
 output OHA; 
 output OHB; 
 output OHC; 
 output OHD; 
 output OHE; 
 output OHF; 
 output OHG; 
 output OHH; 
 output OHI; 
 output OHJ; 
 output OKA; 
 output OKB; 
 output OKC; 
 output OKD; 
 output OKE; 
 output OLD; 
 output OMA; 
 output OMB; 
 output OPA; 
 output OPB; 
 output OPC; 
 output OPD; 
 output OPE; 
 output OPF; 
 output OPG; 
 output OPH; 
 output OPI; 
 output OPK; 
 output OPM; 
 output OPO; 
 output OPQ; 
 output OPR; 
 output OQA; 
 output OQC; 
 output OQE; 
 output OQI; 
 output OQK; 
 output OQM; 
 output OQO; 
 output OQQ; 
  
  
reg  AAA ;
reg  AAB ;
reg  AAC ;
reg  AAD ;
reg  AAE ;
reg  AAF ;
reg  AAG ;
reg  AAH ;
reg  AAI ;
reg  AAJ ;
reg  AAK ;
reg  AAL ;
reg  AAM ;
reg  AAN ;
reg  AAO ;
reg  AAP ;
reg  BAA ;
reg  BAB ;
reg  BAC ;
reg  BAD ;
reg  BAE ;
reg  BAF ;
reg  BAG ;
reg  BAH ;
reg  BAI ;
reg  BAJ ;
reg  BAK ;
reg  BAL ;
reg  BAM ;
reg  BAN ;
reg  BAO ;
reg  BAP ;
reg  bba ;
reg  bbb ;
reg  bbc ;
reg  bbd ;
reg  bbe ;
reg  bbf ;
reg  bbg ;
reg  bbh ;
reg  bbi ;
reg  bbj ;
reg  bbk ;
reg  bbl ;
reg  bbm ;
reg  bbn ;
reg  bbo ;
reg  bbp ;
reg  BCA ;
reg  BCB ;
reg  BCC ;
reg  BCD ;
reg  BCE ;
reg  BCF ;
reg  BCG ;
reg  BCH ;
reg  BCI ;
reg  BCJ ;
reg  BCK ;
reg  BCL ;
reg  BCM ;
reg  BCN ;
reg  BCO ;
reg  BCP ;
reg  BDA ;
reg  BDB ;
reg  BDC ;
reg  BDD ;
reg  BDE ;
reg  BDF ;
reg  BDG ;
reg  BDH ;
reg  BDI ;
reg  BDJ ;
reg  BDK ;
reg  BDL ;
reg  BDM ;
reg  BDN ;
reg  BDO ;
reg  BDP ;
reg  BEA ;
reg  BEB ;
reg  BEC ;
reg  BED ;
reg  BEE ;
reg  BEF ;
reg  BEG ;
reg  BEH ;
reg  BEI ;
reg  BEJ ;
reg  BEK ;
reg  BEL ;
reg  BEM ;
reg  BEN ;
reg  BEO ;
reg  BEP ;
reg  CAC ;
reg  CAD ;
reg  CAE ;
reg  CAF ;
reg  CAG ;
reg  CAH ;
reg  CAI ;
reg  CAJ ;
reg  CAK ;
reg  CAL ;
reg  CAM ;
reg  CAN ;
reg  CAO ;
reg  CAP ;
reg  CBA ;
reg  CBB ;
reg  CBC ;
reg  CBD ;
reg  CBE ;
reg  CBF ;
reg  CBG ;
reg  CBH ;
reg  CBI ;
reg  CBJ ;
reg  CBK ;
reg  CBL ;
reg  CBM ;
reg  CBN ;
reg  CBO ;
reg  CBP ;
reg  CCA ;
reg  CCB ;
reg  CCC ;
reg  CCD ;
reg  CCE ;
reg  CCF ;
reg  CCG ;
reg  CCH ;
reg  CCI ;
reg  CCJ ;
reg  CCK ;
reg  CCL ;
reg  CCM ;
reg  CCN ;
reg  CCO ;
reg  CCP ;
reg  CDC ;
reg  CDD ;
reg  CDE ;
reg  CDF ;
reg  CDG ;
reg  CDH ;
reg  CDI ;
reg  CDJ ;
reg  CDK ;
reg  CDL ;
reg  CDM ;
reg  CDN ;
reg  CDO ;
reg  CDP ;
reg  CEA ;
reg  CEB ;
reg  CEC ;
reg  CED ;
reg  CEE ;
reg  CEF ;
reg  CEG ;
reg  CEH ;
reg  CEI ;
reg  CEJ ;
reg  CEK ;
reg  CEL ;
reg  CEM ;
reg  CEN ;
reg  CEO ;
reg  CEP ;
reg  CFA ;
reg  CFB ;
reg  CFC ;
reg  CFD ;
reg  CFE ;
reg  CFF ;
reg  CFG ;
reg  CFH ;
reg  CFI ;
reg  CFJ ;
reg  CFK ;
reg  CFL ;
reg  CFM ;
reg  CFN ;
reg  CFO ;
reg  CFP ;
reg  DAC ;
reg  DAD ;
reg  DAE ;
reg  DAF ;
reg  DAG ;
reg  DAH ;
reg  DAI ;
reg  DAJ ;
reg  DAK ;
reg  DAL ;
reg  DAM ;
reg  DAN ;
reg  DAO ;
reg  DAP ;
reg  DBA ;
reg  DBB ;
reg  DBC ;
reg  DBD ;
reg  DBE ;
reg  DBF ;
reg  DBG ;
reg  DBH ;
reg  DBI ;
reg  DBJ ;
reg  DBK ;
reg  DBL ;
reg  DBM ;
reg  DBN ;
reg  DBO ;
reg  DBP ;
reg  DCA ;
reg  DCB ;
reg  DCC ;
reg  DCD ;
reg  DCE ;
reg  DCF ;
reg  DCG ;
reg  DCH ;
reg  DCI ;
reg  DCJ ;
reg  DCK ;
reg  DCL ;
reg  DCM ;
reg  DCN ;
reg  DCO ;
reg  DCP ;
reg  ddf ;
reg  ddg ;
reg  ddh ;
reg  ddi ;
reg  ddj ;
reg  ddk ;
reg  ddl ;
reg  ddm ;
reg  ddn ;
reg  ddo ;
reg  ddp ;
reg  dea ;
reg  deb ;
reg  dec ;
reg  ded ;
reg  dee ;
reg  def ;
reg  deg ;
reg  deh ;
reg  dei ;
reg  dej ;
reg  dek ;
reg  del ;
reg  dem ;
reg  den ;
reg  deo ;
reg  dep ;
reg  dfa ;
reg  dfb ;
reg  dfc ;
reg  dfd ;
reg  dfe ;
reg  dff ;
reg  dfg ;
reg  dfh ;
reg  dfi ;
reg  dfj ;
reg  dfk ;
reg  dfl ;
reg  dfm ;
reg  dfn ;
reg  dfo ;
reg  dfp ;
reg  DGA ;
reg  DGB ;
reg  DGC ;
reg  DGD ;
reg  DGE ;
reg  DGF ;
reg  DGG ;
reg  DGH ;
reg  DGI ;
reg  DGJ ;
reg  DGK ;
reg  DGL ;
reg  DGM ;
reg  DGN ;
reg  DGO ;
reg  DGP ;
reg  DHA ;
reg  DHB ;
reg  DHC ;
reg  DHD ;
reg  DHE ;
reg  DHF ;
reg  DHG ;
reg  DHH ;
reg  DHI ;
reg  DHJ ;
reg  DHK ;
reg  DHL ;
reg  DHM ;
reg  DHN ;
reg  DHO ;
reg  DHP ;
reg  FAA ;
reg  FAB ;
reg  FAC ;
reg  FAD ;
reg  FAE ;
reg  FAF ;
reg  FAG ;
reg  FAH ;
reg  FAI ;
reg  FAJ ;
reg  FAK ;
reg  FAL ;
reg  FAM ;
reg  FAN ;
reg  FAO ;
reg  FAP ;
reg  FAQ ;
reg  fba ;
reg  fbb ;
reg  fbc ;
reg  fbd ;
reg  fbe ;
reg  fbf ;
reg  fbg ;
reg  fbh ;
reg  fbi ;
reg  fbj ;
reg  fbk ;
reg  fbl ;
reg  fbm ;
reg  fbn ;
reg  fbo ;
reg  FCA ;
reg  FCB ;
reg  FCC ;
reg  FCD ;
reg  FCE ;
reg  FCF ;
reg  FCG ;
reg  FCH ;
reg  FCI ;
reg  FCJ ;
reg  FCK ;
reg  FCL ;
reg  FCM ;
reg  FCN ;
reg  FCO ;
reg  FCP ;
reg  fda ;
reg  fdb ;
reg  fdc ;
reg  fdd ;
reg  fde ;
reg  fdf ;
reg  fdg ;
reg  fdh ;
reg  fdi ;
reg  fdj ;
reg  fdk ;
reg  fdl ;
reg  fdm ;
reg  fdn ;
reg  fdo ;
reg  FEA ;
reg  FEB ;
reg  FEC ;
reg  FED ;
reg  FEE ;
reg  FEF ;
reg  FEG ;
reg  FEH ;
reg  FEI ;
reg  FEJ ;
reg  FEK ;
reg  FEL ;
reg  FEM ;
reg  FEN ;
reg  FEO ;
reg  ffa ;
reg  ffb ;
reg  ffc ;
reg  ffd ;
reg  ffe ;
reg  fff ;
reg  ffg ;
reg  ffh ;
reg  ffi ;
reg  ffj ;
reg  ffk ;
reg  ffl ;
reg  ffm ;
reg  ffn ;
reg  ffo ;
reg  FGA ;
reg  FGB ;
reg  FGC ;
reg  FGD ;
reg  FGE ;
reg  FGF ;
reg  FGG ;
reg  FGH ;
reg  FGI ;
reg  FGJ ;
reg  FGK ;
reg  FGL ;
reg  FGM ;
reg  FGN ;
reg  FGO ;
reg  FGP ;
reg  fha ;
reg  fhb ;
reg  fhc ;
reg  fhd ;
reg  fhe ;
reg  fhf ;
reg  fhg ;
reg  fhh ;
reg  fhi ;
reg  fhj ;
reg  fhk ;
reg  fhl ;
reg  fhm ;
reg  fhn ;
reg  FIA ;
reg  FIB ;
reg  FIC ;
reg  FID ;
reg  FIE ;
reg  FIF ;
reg  FIG ;
reg  FIH ;
reg  FII ;
reg  FIJ ;
reg  FIK ;
reg  FIL ;
reg  FIM ;
reg  FIN ;
reg  FIO ;
reg  fja ;
reg  fjb ;
reg  fjc ;
reg  fjd ;
reg  fje ;
reg  fjf ;
reg  fjg ;
reg  fjh ;
reg  fji ;
reg  fjj ;
reg  fjk ;
reg  fjl ;
reg  fjm ;
reg  fjn ;
reg  FKA ;
reg  FKB ;
reg  FKC ;
reg  FKD ;
reg  FKE ;
reg  FKF ;
reg  FKG ;
reg  FKH ;
reg  FKI ;
reg  FKJ ;
reg  FKK ;
reg  FKL ;
reg  FKM ;
reg  FKN ;
reg  fla ;
reg  flb ;
reg  flc ;
reg  fld ;
reg  fle ;
reg  flf ;
reg  flg ;
reg  flh ;
reg  fli ;
reg  flj ;
reg  flk ;
reg  fll ;
reg  flm ;
reg  fln ;
reg  FMA ;
reg  FMB ;
reg  FMC ;
reg  FMD ;
reg  FME ;
reg  FMF ;
reg  FMG ;
reg  FMH ;
reg  FMI ;
reg  FMJ ;
reg  FMK ;
reg  FML ;
reg  FMM ;
reg  FMN ;
reg  FMO ;
reg  fna ;
reg  fnb ;
reg  fnc ;
reg  fnd ;
reg  fne ;
reg  fnf ;
reg  fng ;
reg  fnh ;
reg  fni ;
reg  fnj ;
reg  fnk ;
reg  fnl ;
reg  fnm ;
reg  FOA ;
reg  FOB ;
reg  FOC ;
reg  FOD ;
reg  FOE ;
reg  FOF ;
reg  FOG ;
reg  FOH ;
reg  FOI ;
reg  FOJ ;
reg  FOK ;
reg  FOL ;
reg  FOM ;
reg  FON ;
reg  fpa ;
reg  fpb ;
reg  fpc ;
reg  fpd ;
reg  fpe ;
reg  fpf ;
reg  fpg ;
reg  fph ;
reg  fpi ;
reg  fpj ;
reg  fpk ;
reg  fpl ;
reg  fpm ;
reg  FQA ;
reg  FQB ;
reg  FQC ;
reg  FQD ;
reg  FQE ;
reg  FQF ;
reg  FQG ;
reg  FQH ;
reg  FQI ;
reg  FQJ ;
reg  FQK ;
reg  FQL ;
reg  FQM ;
reg  HAA ;
reg  HAB ;
reg  HAC ;
reg  HAD ;
reg  HAF ;
reg  HAG ;
reg  HAH ;
reg  HAI ;
reg  hba ;
reg  hbb ;
reg  hbc ;
reg  hbd ;
reg  hbf ;
reg  hbg ;
reg  HCA ;
reg  HCB ;
reg  HCC ;
reg  HCD ;
reg  HCE ;
reg  HCF ;
reg  hda ;
reg  hdb ;
reg  hdc ;
reg  hdd ;
reg  hde ;
reg  HEA ;
reg  HEB ;
reg  HEC ;
reg  HED ;
reg  HEE ;
reg  HEF ;
reg  HEG ;
reg  HEH ;
reg  hfa ;
reg  hfb ;
reg  hfc ;
reg  hfd ;
reg  hfe ;
reg  hff ;
reg  HGA ;
reg  HGB ;
reg  HGC ;
reg  HGD ;
reg  HGE ;
reg  HGF ;
reg  HGG ;
reg  hha ;
reg  hhb ;
reg  hhc ;
reg  hhd ;
reg  hhe ;
reg  hhf ;
reg  hhg ;
reg  HIA ;
reg  HIB ;
reg  HIC ;
reg  HID ;
reg  HIE ;
reg  HIF ;
reg  HIG ;
reg  hja ;
reg  hjb ;
reg  hjc ;
reg  hjd ;
reg  hje ;
reg  hjf ;
reg  hjg ;
reg  HKA ;
reg  HKB ;
reg  HKC ;
reg  HKD ;
reg  HKE ;
reg  HKF ;
reg  HKG ;
reg  hla ;
reg  hlb ;
reg  hlc ;
reg  hld ;
reg  hle ;
reg  hlf ;
reg  HMA ;
reg  HMB ;
reg  HMC ;
reg  HMD ;
reg  HME ;
reg  HMF ;
reg  HMG ;
reg  HMH ;
reg  hna ;
reg  hnb ;
reg  hnc ;
reg  hnd ;
reg  hne ;
reg  hnf ;
reg  HOA ;
reg  HOB ;
reg  HOC ;
reg  HOD ;
reg  HOE ;
reg  HOF ;
reg  hpa ;
reg  hpb ;
reg  hpc ;
reg  hpd ;
reg  hpe ;
reg  hpf ;
reg  HQA ;
reg  HQB ;
reg  HQC ;
reg  HQD ;
reg  HQE ;
reg  HQF ;
reg  HQG ;
reg  KAA ;
reg  KAB ;
reg  KAC ;
reg  KAD ;
reg  KAE ;
reg  KAF ;
reg  kba ;
reg  kbb ;
reg  kbc ;
reg  kbd ;
reg  KCA ;
reg  KCB ;
reg  KCC ;
reg  KCD ;
reg  KCE ;
reg  kda ;
reg  kdb ;
reg  kdc ;
reg  KEA ;
reg  KEB ;
reg  KEC ;
reg  kfa ;
reg  kfb ;
reg  kfc ;
reg  KGA ;
reg  KGB ;
reg  KGC ;
reg  kha ;
reg  khb ;
reg  khc ;
reg  KIA ;
reg  KIB ;
reg  KIC ;
reg  KID ;
reg  kja ;
reg  kjb ;
reg  kjc ;
reg  KKA ;
reg  KKB ;
reg  KKC ;
reg  KKD ;
reg  kla ;
reg  klb ;
reg  klc ;
reg  KMA ;
reg  KMB ;
reg  KMC ;
reg  KMD ;
reg  kna ;
reg  knb ;
reg  knc ;
reg  KOA ;
reg  KOB ;
reg  KOC ;
reg  KOD ;
reg  kpa ;
reg  kpb ;
reg  KQA ;
reg  KQB ;
reg  KQC ;
reg  MAA ;
reg  MAB ;
reg  MAC ;
reg  MAD ;
reg  mba ;
reg  mbb ;
reg  MCA ;
reg  MCB ;
reg  mda ;
reg  mdb ;
reg  MEA ;
reg  MEB ;
reg  MEC ;
reg  mfa ;
reg  MGA ;
reg  MGB ;
reg  mha ;
reg  MIA ;
reg  MIB ;
reg  MIC ;
reg  mja ;
reg  MKA ;
reg  MKB ;
reg  MKC ;
reg  mla ;
reg  MMA ;
reg  MMB ;
reg  MMC ;
reg  mna ;
reg  MOA ;
reg  MOB ;
reg  MOC ;
reg  mpa ;
reg  MQA ;
reg  MQB ;
reg  MQC ;
reg  OAA ;
reg  OAB ;
reg  OAC ;
reg  OAD ;
reg  OAE ;
reg  OAF ;
reg  OAG ;
reg  OAH ;
reg  OAI ;
reg  OAJ ;
reg  OAK ;
reg  OAL ;
reg  OAM ;
reg  OAN ;
reg  OAO ;
reg  OAP ;
reg  OBA ;
reg  OBB ;
reg  OBC ;
reg  OBD ;
reg  OBE ;
reg  OBF ;
reg  OBG ;
reg  OBH ;
reg  OBI ;
reg  OBJ ;
reg  OBK ;
reg  OBL ;
reg  OBM ;
reg  OBN ;
reg  OBO ;
reg  OBP ;
reg  oca ;
reg  ocb ;
reg  occ ;
reg  ocd ;
reg  oce ;
reg  ocf ;
reg  ocg ;
reg  och ;
reg  oci ;
reg  ocj ;
reg  ock ;
reg  ocl ;
reg  ocm ;
reg  ocn ;
reg  oco ;
reg  ocp ;
reg  oda ;
reg  odb ;
reg  odc ;
reg  odd ;
reg  ode ;
reg  odf ;
reg  odg ;
reg  odh ;
reg  odi ;
reg  odj ;
reg  odk ;
reg  odl ;
reg  odm ;
reg  odn ;
reg  odo ;
reg  odp ;
reg  oga ;
reg  ogb ;
reg  ogc ;
reg  ogd ;
reg  oge ;
reg  ogf ;
reg  ogg ;
reg  ogh ;
reg  ogi ;
reg  ogj ;
reg  ogk ;
reg  ogl ;
reg  ogm ;
reg  oha ;
reg  ohb ;
reg  ohc ;
reg  ohd ;
reg  ohe ;
reg  ohf ;
reg  OHG ;
reg  OHH ;
reg  OHI ;
reg  OHJ ;
reg  oig ;
reg  oih ;
reg  oka ;
reg  okb ;
reg  okc ;
reg  OKD ;
reg  OKE ;
reg  old ;
reg  oma ;
reg  OMB ;
reg  OPA ;
reg  OPB ;
reg  OPC ;
reg  OPD ;
reg  OPE ;
reg  OPF ;
reg  OPG ;
reg  OPH ;
reg  OPI ;
reg  OPK ;
reg  OPM ;
reg  OPO ;
reg  OPQ ;
reg  OPR ;
reg  oqa ;
reg  oqc ;
reg  oqe ;
reg  oqi ;
reg  oqk ;
reg  oqm ;
reg  oqo ;
reg  oqq ;
reg  QAA ;
reg  QGA ;
reg  QHA ;
reg  QIA ;
reg  QIB ;
reg  QIC ;
reg  QID ;
reg  QIE ;
reg  QKA ;
reg  QTA ;
reg  QTB ;
reg  TGA ;
reg  TGB ;
reg  TGC ;
reg  THA ;
reg  THB ;
reg  THC ;
reg  THD ;
reg  THE ;
reg  THF ;
reg  TKA ;
reg  TKB ;
reg  TKC ;
reg  TKD ;
reg  TKE ;
reg  TKF ;
reg  TRA ;
reg  TRB ;
reg  TSA ;
reg  TSB ;
reg  TSC ;
reg  TSD ;
reg  TSE ;
reg  TSF ;
reg  TTA ;
reg  TTB ;
reg  TTC ;
wire  aaa ;
wire  aab ;
wire  aac ;
wire  aad ;
wire  aae ;
wire  aaf ;
wire  aag ;
wire  aah ;
wire  aai ;
wire  aaj ;
wire  aak ;
wire  aal ;
wire  aam ;
wire  aan ;
wire  aao ;
wire  aap ;
wire  baa ;
wire  bab ;
wire  bac ;
wire  bad ;
wire  bae ;
wire  baf ;
wire  bag ;
wire  bah ;
wire  bai ;
wire  baj ;
wire  bak ;
wire  bal ;
wire  bam ;
wire  ban ;
wire  bao ;
wire  bap ;
wire  BBA ;
wire  BBB ;
wire  BBC ;
wire  BBD ;
wire  BBE ;
wire  BBF ;
wire  BBG ;
wire  BBH ;
wire  BBI ;
wire  BBJ ;
wire  BBK ;
wire  BBL ;
wire  BBM ;
wire  BBN ;
wire  BBO ;
wire  BBP ;
wire  bca ;
wire  bcb ;
wire  bcc ;
wire  bcd ;
wire  bce ;
wire  bcf ;
wire  bcg ;
wire  bch ;
wire  bci ;
wire  bcj ;
wire  bck ;
wire  bcl ;
wire  bcm ;
wire  bcn ;
wire  bco ;
wire  bcp ;
wire  bda ;
wire  bdb ;
wire  bdc ;
wire  bdd ;
wire  bde ;
wire  bdf ;
wire  bdg ;
wire  bdh ;
wire  bdi ;
wire  bdj ;
wire  bdk ;
wire  bdl ;
wire  bdm ;
wire  bdn ;
wire  bdo ;
wire  bdp ;
wire  bea ;
wire  beb ;
wire  bec ;
wire  bed ;
wire  bee ;
wire  bef ;
wire  beg ;
wire  beh ;
wire  bei ;
wire  bej ;
wire  bek ;
wire  bel ;
wire  bem ;
wire  ben ;
wire  beo ;
wire  bep ;
wire  cac ;
wire  cad ;
wire  cae ;
wire  caf ;
wire  cag ;
wire  cah ;
wire  cai ;
wire  caj ;
wire  cak ;
wire  cal ;
wire  cam ;
wire  can ;
wire  cao ;
wire  cap ;
wire  cba ;
wire  cbb ;
wire  cbc ;
wire  cbd ;
wire  cbe ;
wire  cbf ;
wire  cbg ;
wire  cbh ;
wire  cbi ;
wire  cbj ;
wire  cbk ;
wire  cbl ;
wire  cbm ;
wire  cbn ;
wire  cbo ;
wire  cbp ;
wire  cca ;
wire  ccb ;
wire  ccc ;
wire  ccd ;
wire  cce ;
wire  ccf ;
wire  ccg ;
wire  cch ;
wire  cci ;
wire  ccj ;
wire  cck ;
wire  ccl ;
wire  ccm ;
wire  ccn ;
wire  cco ;
wire  ccp ;
wire  cdc ;
wire  cdd ;
wire  cde ;
wire  cdf ;
wire  cdg ;
wire  cdh ;
wire  cdi ;
wire  cdj ;
wire  cdk ;
wire  cdl ;
wire  cdm ;
wire  cdn ;
wire  cdo ;
wire  cdp ;
wire  cea ;
wire  ceb ;
wire  cec ;
wire  ced ;
wire  cee ;
wire  cef ;
wire  ceg ;
wire  ceh ;
wire  cei ;
wire  cej ;
wire  cek ;
wire  cel ;
wire  cem ;
wire  cen ;
wire  ceo ;
wire  cep ;
wire  cfa ;
wire  cfb ;
wire  cfc ;
wire  cfd ;
wire  cfe ;
wire  cff ;
wire  cfg ;
wire  cfh ;
wire  cfi ;
wire  cfj ;
wire  cfk ;
wire  cfl ;
wire  cfm ;
wire  cfn ;
wire  cfo ;
wire  cfp ;
wire  dac ;
wire  dad ;
wire  dae ;
wire  daf ;
wire  dag ;
wire  dah ;
wire  dai ;
wire  daj ;
wire  dak ;
wire  dal ;
wire  dam ;
wire  dan ;
wire  dao ;
wire  dap ;
wire  dba ;
wire  dbb ;
wire  dbc ;
wire  dbd ;
wire  dbe ;
wire  dbf ;
wire  dbg ;
wire  dbh ;
wire  dbi ;
wire  dbj ;
wire  dbk ;
wire  dbl ;
wire  dbm ;
wire  dbn ;
wire  dbo ;
wire  dbp ;
wire  dca ;
wire  dcb ;
wire  dcc ;
wire  dcd ;
wire  dce ;
wire  dcf ;
wire  dcg ;
wire  dch ;
wire  dci ;
wire  dcj ;
wire  dck ;
wire  dcl ;
wire  dcm ;
wire  dcn ;
wire  dco ;
wire  dcp ;
wire  DDF ;
wire  DDG ;
wire  DDH ;
wire  DDI ;
wire  DDJ ;
wire  DDK ;
wire  DDL ;
wire  DDM ;
wire  DDN ;
wire  DDO ;
wire  DDP ;
wire  DEA ;
wire  DEB ;
wire  DEC ;
wire  DED ;
wire  DEE ;
wire  DEF ;
wire  DEG ;
wire  DEH ;
wire  DEI ;
wire  DEJ ;
wire  DEK ;
wire  DEL ;
wire  DEM ;
wire  DEN ;
wire  DEO ;
wire  DEP ;
wire  DFA ;
wire  DFB ;
wire  DFC ;
wire  DFD ;
wire  DFE ;
wire  DFF ;
wire  DFG ;
wire  DFH ;
wire  DFI ;
wire  DFJ ;
wire  DFK ;
wire  DFL ;
wire  DFM ;
wire  DFN ;
wire  DFO ;
wire  DFP ;
wire  dga ;
wire  dgb ;
wire  dgc ;
wire  dgd ;
wire  dge ;
wire  dgf ;
wire  dgg ;
wire  dgh ;
wire  dgi ;
wire  dgj ;
wire  dgk ;
wire  dgl ;
wire  dgm ;
wire  dgn ;
wire  dgo ;
wire  dgp ;
wire  dha ;
wire  dhb ;
wire  dhc ;
wire  dhd ;
wire  dhe ;
wire  dhf ;
wire  dhg ;
wire  dhh ;
wire  dhi ;
wire  dhj ;
wire  dhk ;
wire  dhl ;
wire  dhm ;
wire  dhn ;
wire  dho ;
wire  dhp ;
wire  eac ;
wire  EAC ;
wire  ead ;
wire  EAD ;
wire  eae ;
wire  EAE ;
wire  eaf ;
wire  EAF ;
wire  eag ;
wire  EAG ;
wire  eah ;
wire  EAH ;
wire  eai ;
wire  EAI ;
wire  eaj ;
wire  EAJ ;
wire  eak ;
wire  EAK ;
wire  eal ;
wire  EAL ;
wire  eam ;
wire  EAM ;
wire  ean ;
wire  EAN ;
wire  eao ;
wire  EAO ;
wire  eap ;
wire  EAP ;
wire  eaq ;
wire  EAQ ;
wire  ear ;
wire  EAR ;
wire  eas ;
wire  EAS ;
wire  eat ;
wire  EAT ;
wire  eau ;
wire  EAU ;
wire  eav ;
wire  EAV ;
wire  eaw ;
wire  EAW ;
wire  eax ;
wire  EAX ;
wire  eba ;
wire  EBA ;
wire  ebb ;
wire  EBB ;
wire  ebc ;
wire  EBC ;
wire  ebd ;
wire  EBD ;
wire  ebe ;
wire  EBE ;
wire  ebf ;
wire  EBF ;
wire  ebg ;
wire  EBG ;
wire  ebh ;
wire  EBH ;
wire  ebi ;
wire  EBI ;
wire  ebj ;
wire  EBJ ;
wire  ebk ;
wire  EBK ;
wire  ebl ;
wire  EBL ;
wire  ebm ;
wire  EBM ;
wire  ebn ;
wire  EBN ;
wire  ebo ;
wire  EBO ;
wire  ebp ;
wire  EBP ;
wire  ebq ;
wire  EBQ ;
wire  ebr ;
wire  EBR ;
wire  ebs ;
wire  EBS ;
wire  ebt ;
wire  EBT ;
wire  ebu ;
wire  EBU ;
wire  ebv ;
wire  EBV ;
wire  ebw ;
wire  EBW ;
wire  ebx ;
wire  EBX ;
wire  ecd ;
wire  ECD ;
wire  ece ;
wire  ECE ;
wire  ecf ;
wire  ECF ;
wire  ecg ;
wire  ECG ;
wire  ech ;
wire  ECH ;
wire  eci ;
wire  ECI ;
wire  ecj ;
wire  ECJ ;
wire  eck ;
wire  ECK ;
wire  ecl ;
wire  ECL ;
wire  ecm ;
wire  ECM ;
wire  ecn ;
wire  ECN ;
wire  eco ;
wire  ECO ;
wire  ecp ;
wire  ECP ;
wire  ecq ;
wire  ECQ ;
wire  ecr ;
wire  ECR ;
wire  ecs ;
wire  ECS ;
wire  ect ;
wire  ECT ;
wire  ecu ;
wire  ECU ;
wire  ecv ;
wire  ECV ;
wire  ecw ;
wire  ECW ;
wire  ecx ;
wire  ECX ;
wire  eda ;
wire  EDA ;
wire  edb ;
wire  EDB ;
wire  edc ;
wire  EDC ;
wire  edd ;
wire  EDD ;
wire  ede ;
wire  EDE ;
wire  edf ;
wire  EDF ;
wire  edg ;
wire  EDG ;
wire  edh ;
wire  EDH ;
wire  edi ;
wire  EDI ;
wire  edj ;
wire  EDJ ;
wire  edk ;
wire  EDK ;
wire  edl ;
wire  EDL ;
wire  edm ;
wire  EDM ;
wire  edn ;
wire  EDN ;
wire  edo ;
wire  EDO ;
wire  edp ;
wire  EDP ;
wire  edq ;
wire  EDQ ;
wire  edr ;
wire  EDR ;
wire  eds ;
wire  EDS ;
wire  edt ;
wire  EDT ;
wire  edu ;
wire  EDU ;
wire  edv ;
wire  EDV ;
wire  edw ;
wire  EDW ;
wire  edx ;
wire  EDX ;
wire  eee ;
wire  EEE ;
wire  eef ;
wire  EEF ;
wire  eeg ;
wire  EEG ;
wire  eeh ;
wire  EEH ;
wire  eei ;
wire  EEI ;
wire  eej ;
wire  EEJ ;
wire  eek ;
wire  EEK ;
wire  eel ;
wire  EEL ;
wire  eem ;
wire  EEM ;
wire  een ;
wire  EEN ;
wire  eeo ;
wire  EEO ;
wire  eep ;
wire  EEP ;
wire  eeq ;
wire  EEQ ;
wire  eer ;
wire  EER ;
wire  ees ;
wire  EES ;
wire  eet ;
wire  EET ;
wire  eeu ;
wire  EEU ;
wire  eev ;
wire  EEV ;
wire  eew ;
wire  EEW ;
wire  eex ;
wire  EEX ;
wire  efa ;
wire  EFA ;
wire  efb ;
wire  EFB ;
wire  efc ;
wire  EFC ;
wire  efd ;
wire  EFD ;
wire  efe ;
wire  EFE ;
wire  eff ;
wire  EFF ;
wire  efg ;
wire  EFG ;
wire  efh ;
wire  EFH ;
wire  efi ;
wire  EFI ;
wire  efj ;
wire  EFJ ;
wire  efk ;
wire  EFK ;
wire  efl ;
wire  EFL ;
wire  efm ;
wire  EFM ;
wire  efn ;
wire  EFN ;
wire  efo ;
wire  EFO ;
wire  efp ;
wire  EFP ;
wire  efq ;
wire  EFQ ;
wire  efr ;
wire  EFR ;
wire  efs ;
wire  EFS ;
wire  eft ;
wire  EFT ;
wire  efu ;
wire  EFU ;
wire  efv ;
wire  EFV ;
wire  efw ;
wire  EFW ;
wire  efx ;
wire  EFX ;
wire  egf ;
wire  EGF ;
wire  egg ;
wire  EGG ;
wire  egh ;
wire  EGH ;
wire  egi ;
wire  EGI ;
wire  egj ;
wire  EGJ ;
wire  egk ;
wire  EGK ;
wire  egl ;
wire  EGL ;
wire  egm ;
wire  EGM ;
wire  egn ;
wire  EGN ;
wire  ego ;
wire  EGO ;
wire  egp ;
wire  EGP ;
wire  egq ;
wire  EGQ ;
wire  egr ;
wire  EGR ;
wire  egs ;
wire  EGS ;
wire  egt ;
wire  EGT ;
wire  egu ;
wire  EGU ;
wire  egv ;
wire  EGV ;
wire  egw ;
wire  EGW ;
wire  egx ;
wire  EGX ;
wire  eha ;
wire  EHA ;
wire  ehb ;
wire  EHB ;
wire  ehc ;
wire  EHC ;
wire  ehd ;
wire  EHD ;
wire  ehe ;
wire  EHE ;
wire  ehf ;
wire  EHF ;
wire  ehg ;
wire  EHG ;
wire  ehh ;
wire  EHH ;
wire  ehi ;
wire  EHI ;
wire  ehj ;
wire  EHJ ;
wire  ehk ;
wire  EHK ;
wire  ehl ;
wire  EHL ;
wire  ehm ;
wire  EHM ;
wire  ehn ;
wire  EHN ;
wire  eho ;
wire  EHO ;
wire  ehp ;
wire  EHP ;
wire  ehq ;
wire  EHQ ;
wire  ehr ;
wire  EHR ;
wire  ehs ;
wire  EHS ;
wire  eht ;
wire  EHT ;
wire  ehu ;
wire  EHU ;
wire  ehv ;
wire  EHV ;
wire  ehw ;
wire  EHW ;
wire  ehx ;
wire  EHX ;
wire  eig ;
wire  EIG ;
wire  eih ;
wire  EIH ;
wire  eii ;
wire  EII ;
wire  eij ;
wire  EIJ ;
wire  eik ;
wire  EIK ;
wire  eil ;
wire  EIL ;
wire  eim ;
wire  EIM ;
wire  ein ;
wire  EIN ;
wire  eio ;
wire  EIO ;
wire  eip ;
wire  EIP ;
wire  eiq ;
wire  EIQ ;
wire  eir ;
wire  EIR ;
wire  eis ;
wire  EIS ;
wire  eit ;
wire  EIT ;
wire  eiu ;
wire  EIU ;
wire  eiv ;
wire  EIV ;
wire  eiw ;
wire  EIW ;
wire  eix ;
wire  EIX ;
wire  eja ;
wire  EJA ;
wire  ejb ;
wire  EJB ;
wire  ejc ;
wire  EJC ;
wire  ejd ;
wire  EJD ;
wire  eje ;
wire  EJE ;
wire  ejf ;
wire  EJF ;
wire  ejg ;
wire  EJG ;
wire  ejh ;
wire  EJH ;
wire  eji ;
wire  EJI ;
wire  ejj ;
wire  EJJ ;
wire  ejk ;
wire  EJK ;
wire  ejl ;
wire  EJL ;
wire  ejm ;
wire  EJM ;
wire  ejn ;
wire  EJN ;
wire  ejo ;
wire  EJO ;
wire  ejp ;
wire  EJP ;
wire  ejq ;
wire  EJQ ;
wire  ejr ;
wire  EJR ;
wire  ejs ;
wire  EJS ;
wire  ejt ;
wire  EJT ;
wire  eju ;
wire  EJU ;
wire  ejv ;
wire  EJV ;
wire  ejw ;
wire  EJW ;
wire  ejx ;
wire  EJX ;
wire  ekh ;
wire  EKH ;
wire  eki ;
wire  EKI ;
wire  ekj ;
wire  EKJ ;
wire  ekk ;
wire  EKK ;
wire  ekl ;
wire  EKL ;
wire  ekm ;
wire  EKM ;
wire  ekn ;
wire  EKN ;
wire  eko ;
wire  EKO ;
wire  ekp ;
wire  EKP ;
wire  ekq ;
wire  EKQ ;
wire  ekr ;
wire  EKR ;
wire  eks ;
wire  EKS ;
wire  ekt ;
wire  EKT ;
wire  eku ;
wire  EKU ;
wire  ekv ;
wire  EKV ;
wire  ekw ;
wire  EKW ;
wire  ekx ;
wire  EKX ;
wire  ela ;
wire  ELA ;
wire  elb ;
wire  ELB ;
wire  elc ;
wire  ELC ;
wire  eld ;
wire  ELD ;
wire  ele ;
wire  ELE ;
wire  elf ;
wire  ELF ;
wire  elg ;
wire  ELG ;
wire  elh ;
wire  ELH ;
wire  eli ;
wire  ELI ;
wire  elj ;
wire  ELJ ;
wire  elk ;
wire  ELK ;
wire  ell ;
wire  ELL ;
wire  elm ;
wire  ELM ;
wire  eln ;
wire  ELN ;
wire  elo ;
wire  ELO ;
wire  elp ;
wire  ELP ;
wire  elq ;
wire  ELQ ;
wire  elr ;
wire  ELR ;
wire  els ;
wire  ELS ;
wire  elt ;
wire  ELT ;
wire  elu ;
wire  ELU ;
wire  elv ;
wire  ELV ;
wire  elw ;
wire  ELW ;
wire  elx ;
wire  ELX ;
wire  emi ;
wire  EMI ;
wire  emj ;
wire  EMJ ;
wire  emk ;
wire  EMK ;
wire  eml ;
wire  EML ;
wire  emm ;
wire  EMM ;
wire  emn ;
wire  EMN ;
wire  emo ;
wire  EMO ;
wire  emp ;
wire  EMP ;
wire  emq ;
wire  EMQ ;
wire  emr ;
wire  EMR ;
wire  ems ;
wire  EMS ;
wire  emt ;
wire  EMT ;
wire  emu ;
wire  EMU ;
wire  emv ;
wire  EMV ;
wire  emw ;
wire  EMW ;
wire  emx ;
wire  EMX ;
wire  ena ;
wire  ENA ;
wire  enb ;
wire  ENB ;
wire  enc ;
wire  ENC ;
wire  endd ;
wire  ENDD  ;
wire  ene ;
wire  ENE ;
wire  enf ;
wire  ENF ;
wire  eng ;
wire  ENG ;
wire  enh ;
wire  ENH ;
wire  eni ;
wire  ENI ;
wire  enj ;
wire  ENJ ;
wire  enk ;
wire  ENK ;
wire  enl ;
wire  ENL ;
wire  enm ;
wire  ENM ;
wire  enn ;
wire  ENN ;
wire  eno ;
wire  ENO ;
wire  enp ;
wire  ENP ;
wire  enq ;
wire  ENQ ;
wire  enr ;
wire  ENR ;
wire  ens ;
wire  ENS ;
wire  ent ;
wire  ENT ;
wire  enu ;
wire  ENU ;
wire  env ;
wire  ENV ;
wire  enw ;
wire  ENW ;
wire  enx ;
wire  ENX ;
wire  eoj ;
wire  EOJ ;
wire  eok ;
wire  EOK ;
wire  eol ;
wire  EOL ;
wire  eom ;
wire  EOM ;
wire  eon ;
wire  EON ;
wire  eoo ;
wire  EOO ;
wire  eop ;
wire  EOP ;
wire  eoq ;
wire  EOQ ;
wire  eor ;
wire  EOR ;
wire  eos ;
wire  EOS ;
wire  eot ;
wire  EOT ;
wire  eou ;
wire  EOU ;
wire  eov ;
wire  EOV ;
wire  eow ;
wire  EOW ;
wire  eox ;
wire  EOX ;
wire  epa ;
wire  EPA ;
wire  epb ;
wire  EPB ;
wire  epc ;
wire  EPC ;
wire  epd ;
wire  EPD ;
wire  epe ;
wire  EPE ;
wire  epf ;
wire  EPF ;
wire  epg ;
wire  EPG ;
wire  eph ;
wire  EPH ;
wire  epi ;
wire  EPI ;
wire  epj ;
wire  EPJ ;
wire  epk ;
wire  EPK ;
wire  epl ;
wire  EPL ;
wire  epm ;
wire  EPM ;
wire  epn ;
wire  EPN ;
wire  epo ;
wire  EPO ;
wire  epp ;
wire  EPP ;
wire  epq ;
wire  EPQ ;
wire  epr ;
wire  EPR ;
wire  eps ;
wire  EPS ;
wire  ept ;
wire  EPT ;
wire  epu ;
wire  EPU ;
wire  epv ;
wire  EPV ;
wire  epw ;
wire  EPW ;
wire  epx ;
wire  EPX ;
wire  eqk ;
wire  EQK ;
wire  eql ;
wire  EQL ;
wire  eqm ;
wire  EQM ;
wire  eqn ;
wire  EQN ;
wire  eqo ;
wire  EQO ;
wire  eqp ;
wire  EQP ;
wire  eqq ;
wire  EQQ ;
wire  eqr ;
wire  EQR ;
wire  eqs ;
wire  EQS ;
wire  eqt ;
wire  EQT ;
wire  equ ;
wire  EQU ;
wire  eqv ;
wire  EQV ;
wire  eqw ;
wire  EQW ;
wire  eqx ;
wire  EQX ;
wire  era ;
wire  ERA ;
wire  erb ;
wire  ERB ;
wire  erc ;
wire  ERC ;
wire  erd ;
wire  ERD ;
wire  ere ;
wire  ERE ;
wire  erf ;
wire  ERF ;
wire  erg ;
wire  ERG ;
wire  erh ;
wire  ERH ;
wire  eri ;
wire  ERI ;
wire  erj ;
wire  ERJ ;
wire  erk ;
wire  ERK ;
wire  erl ;
wire  ERL ;
wire  erm ;
wire  ERM ;
wire  ern ;
wire  ERN ;
wire  ero ;
wire  ERO ;
wire  erp ;
wire  ERP ;
wire  erq ;
wire  ERQ ;
wire  err ;
wire  ERR ;
wire  ers ;
wire  ERS ;
wire  ert ;
wire  ERT ;
wire  eru ;
wire  ERU ;
wire  erv ;
wire  ERV ;
wire  erw ;
wire  ERW ;
wire  erx ;
wire  ERX ;
wire  faa ;
wire  fab ;
wire  fac ;
wire  fad ;
wire  fae ;
wire  faf ;
wire  fag ;
wire  fah ;
wire  fai ;
wire  faj ;
wire  fak ;
wire  fal ;
wire  fam ;
wire  fan ;
wire  fao ;
wire  fap ;
wire  faq ;
wire  FBA ;
wire  FBB ;
wire  FBC ;
wire  FBD ;
wire  FBE ;
wire  FBF ;
wire  FBG ;
wire  FBH ;
wire  FBI ;
wire  FBJ ;
wire  FBK ;
wire  FBL ;
wire  FBM ;
wire  FBN ;
wire  FBO ;
wire  fca ;
wire  fcb ;
wire  fcc ;
wire  fcd ;
wire  fce ;
wire  fcf ;
wire  fcg ;
wire  fch ;
wire  fci ;
wire  fcj ;
wire  fck ;
wire  fcl ;
wire  fcm ;
wire  fcn ;
wire  fco ;
wire  fcp ;
wire  FDA ;
wire  FDB ;
wire  FDC ;
wire  FDD ;
wire  FDE ;
wire  FDF ;
wire  FDG ;
wire  FDH ;
wire  FDI ;
wire  FDJ ;
wire  FDK ;
wire  FDL ;
wire  FDM ;
wire  FDN ;
wire  FDO ;
wire  fea ;
wire  feb ;
wire  fec ;
wire  fed ;
wire  fee ;
wire  fef ;
wire  feg ;
wire  feh ;
wire  fei ;
wire  fej ;
wire  fek ;
wire  fel ;
wire  fem ;
wire  fen ;
wire  feo ;
wire  FFA ;
wire  FFB ;
wire  FFC ;
wire  FFD ;
wire  FFE ;
wire  FFF ;
wire  FFG ;
wire  FFH ;
wire  FFI ;
wire  FFJ ;
wire  FFK ;
wire  FFL ;
wire  FFM ;
wire  FFN ;
wire  FFO ;
wire  fga ;
wire  fgb ;
wire  fgc ;
wire  fgd ;
wire  fge ;
wire  fgf ;
wire  fgg ;
wire  fgh ;
wire  fgi ;
wire  fgj ;
wire  fgk ;
wire  fgl ;
wire  fgm ;
wire  fgn ;
wire  fgo ;
wire  fgp ;
wire  FHA ;
wire  FHB ;
wire  FHC ;
wire  FHD ;
wire  FHE ;
wire  FHF ;
wire  FHG ;
wire  FHH ;
wire  FHI ;
wire  FHJ ;
wire  FHK ;
wire  FHL ;
wire  FHM ;
wire  FHN ;
wire  fia ;
wire  fib ;
wire  fic ;
wire  fid ;
wire  fie ;
wire  fif ;
wire  fig ;
wire  fih ;
wire  fii ;
wire  fij ;
wire  fik ;
wire  fil ;
wire  fim ;
wire  fin ;
wire  fio ;
wire  FJA ;
wire  FJB ;
wire  FJC ;
wire  FJD ;
wire  FJE ;
wire  FJF ;
wire  FJG ;
wire  FJH ;
wire  FJI ;
wire  FJJ ;
wire  FJK ;
wire  FJL ;
wire  FJM ;
wire  FJN ;
wire  fka ;
wire  fkb ;
wire  fkc ;
wire  fkd ;
wire  fke ;
wire  fkf ;
wire  fkg ;
wire  fkh ;
wire  fki ;
wire  fkj ;
wire  fkk ;
wire  fkl ;
wire  fkm ;
wire  fkn ;
wire  FLA ;
wire  FLB ;
wire  FLC ;
wire  FLD ;
wire  FLE ;
wire  FLF ;
wire  FLG ;
wire  FLH ;
wire  FLI ;
wire  FLJ ;
wire  FLK ;
wire  FLL ;
wire  FLM ;
wire  FLN ;
wire  fma ;
wire  fmb ;
wire  fmc ;
wire  fmd ;
wire  fme ;
wire  fmf ;
wire  fmg ;
wire  fmh ;
wire  fmi ;
wire  fmj ;
wire  fmk ;
wire  fml ;
wire  fmm ;
wire  fmn ;
wire  fmo ;
wire  FNA ;
wire  FNB ;
wire  FNC ;
wire  FND ;
wire  FNE ;
wire  FNF ;
wire  FNG ;
wire  FNH ;
wire  FNI ;
wire  FNJ ;
wire  FNK ;
wire  FNL ;
wire  FNM ;
wire  foa ;
wire  fob ;
wire  foc ;
wire  fod ;
wire  foe ;
wire  fof ;
wire  fog ;
wire  foh ;
wire  foi ;
wire  foj ;
wire  fok ;
wire  fol ;
wire  fom ;
wire  fon ;
wire  FPA ;
wire  FPB ;
wire  FPC ;
wire  FPD ;
wire  FPE ;
wire  FPF ;
wire  FPG ;
wire  FPH ;
wire  FPI ;
wire  FPJ ;
wire  FPK ;
wire  FPL ;
wire  FPM ;
wire  fqa ;
wire  fqb ;
wire  fqc ;
wire  fqd ;
wire  fqe ;
wire  fqf ;
wire  fqg ;
wire  fqh ;
wire  fqi ;
wire  fqj ;
wire  fqk ;
wire  fql ;
wire  fqm ;
wire  gaa ;
wire  GAA ;
wire  gab ;
wire  GAB ;
wire  gac ;
wire  GAC ;
wire  gad ;
wire  GAD ;
wire  gae ;
wire  GAE ;
wire  gba ;
wire  GBA ;
wire  gbb ;
wire  GBB ;
wire  gbc ;
wire  GBC ;
wire  gbd ;
wire  GBD ;
wire  gbe ;
wire  GBE ;
wire  gca ;
wire  GCA ;
wire  gcb ;
wire  GCB ;
wire  gcc ;
wire  GCC ;
wire  gcd ;
wire  GCD ;
wire  gce ;
wire  GCE ;
wire  gcf ;
wire  GCF ;
wire  gcg ;
wire  GCG ;
wire  gch ;
wire  GCH ;
wire  gci ;
wire  GCI ;
wire  gcj ;
wire  GCJ ;
wire  gda ;
wire  GDA ;
wire  gdb ;
wire  GDB ;
wire  gdc ;
wire  GDC ;
wire  gdd ;
wire  GDD ;
wire  gde ;
wire  GDE ;
wire  gdf ;
wire  GDF ;
wire  gdg ;
wire  GDG ;
wire  gdh ;
wire  GDH ;
wire  gdi ;
wire  GDI ;
wire  gdj ;
wire  GDJ ;
wire  gea ;
wire  GEA ;
wire  geb ;
wire  GEB ;
wire  gec ;
wire  GEC ;
wire  ged ;
wire  GED ;
wire  gee ;
wire  GEE ;
wire  gef ;
wire  GEF ;
wire  geg ;
wire  GEG ;
wire  geh ;
wire  GEH ;
wire  gei ;
wire  GEI ;
wire  gej ;
wire  GEJ ;
wire  gfa ;
wire  GFA ;
wire  gfb ;
wire  GFB ;
wire  gfc ;
wire  GFC ;
wire  gfd ;
wire  GFD ;
wire  gfe ;
wire  GFE ;
wire  gff ;
wire  GFF ;
wire  gfg ;
wire  GFG ;
wire  gfh ;
wire  GFH ;
wire  gfi ;
wire  GFI ;
wire  gfj ;
wire  GFJ ;
wire  gga ;
wire  GGA ;
wire  ggb ;
wire  GGB ;
wire  ggc ;
wire  GGC ;
wire  ggd ;
wire  GGD ;
wire  gge ;
wire  GGE ;
wire  ggf ;
wire  GGF ;
wire  ggg ;
wire  GGG ;
wire  ggh ;
wire  GGH ;
wire  ggi ;
wire  GGI ;
wire  ggj ;
wire  GGJ ;
wire  gha ;
wire  GHA ;
wire  ghb ;
wire  GHB ;
wire  ghc ;
wire  GHC ;
wire  ghd ;
wire  GHD ;
wire  ghe ;
wire  GHE ;
wire  ghf ;
wire  GHF ;
wire  ghg ;
wire  GHG ;
wire  ghh ;
wire  GHH ;
wire  ghi ;
wire  GHI ;
wire  ghj ;
wire  GHJ ;
wire  gia ;
wire  GIA ;
wire  gib ;
wire  GIB ;
wire  gic ;
wire  GIC ;
wire  gid ;
wire  GID ;
wire  gie ;
wire  GIE ;
wire  gif ;
wire  GIF ;
wire  gig ;
wire  GIG ;
wire  gih ;
wire  GIH ;
wire  gii ;
wire  GII ;
wire  gja ;
wire  GJA ;
wire  gjb ;
wire  GJB ;
wire  gjc ;
wire  GJC ;
wire  gjd ;
wire  GJD ;
wire  gje ;
wire  GJE ;
wire  gjf ;
wire  GJF ;
wire  gjg ;
wire  GJG ;
wire  gjh ;
wire  GJH ;
wire  gji ;
wire  GJI ;
wire  gka ;
wire  GKA ;
wire  gkb ;
wire  GKB ;
wire  gkc ;
wire  GKC ;
wire  gkd ;
wire  GKD ;
wire  gke ;
wire  GKE ;
wire  gkf ;
wire  GKF ;
wire  gkg ;
wire  GKG ;
wire  gkh ;
wire  GKH ;
wire  gki ;
wire  GKI ;
wire  gla ;
wire  GLA ;
wire  glb ;
wire  GLB ;
wire  glc ;
wire  GLC ;
wire  gld ;
wire  GLD ;
wire  gle ;
wire  GLE ;
wire  glf ;
wire  GLF ;
wire  glg ;
wire  GLG ;
wire  glh ;
wire  GLH ;
wire  gli ;
wire  GLI ;
wire  gma ;
wire  GMA ;
wire  gmb ;
wire  GMB ;
wire  gmc ;
wire  GMC ;
wire  gmd ;
wire  GMD ;
wire  gme ;
wire  GME ;
wire  gmf ;
wire  GMF ;
wire  gmg ;
wire  GMG ;
wire  gmh ;
wire  GMH ;
wire  gmi ;
wire  GMI ;
wire  gna ;
wire  GNA ;
wire  gnb ;
wire  GNB ;
wire  gnc ;
wire  GNC ;
wire  gnd ;
wire  GND ;
wire  gne ;
wire  GNE ;
wire  gnf ;
wire  GNF ;
wire  gng ;
wire  GNG ;
wire  gnh ;
wire  GNH ;
wire  gni ;
wire  GNI ;
wire  goa ;
wire  GOA ;
wire  gob ;
wire  GOB ;
wire  goc ;
wire  GOC ;
wire  god ;
wire  GOD ;
wire  goe ;
wire  GOE ;
wire  gof ;
wire  GOF ;
wire  gog ;
wire  GOG ;
wire  goh ;
wire  GOH ;
wire  goi ;
wire  GOI ;
wire  gpa ;
wire  GPA ;
wire  gpb ;
wire  GPB ;
wire  gpc ;
wire  GPC ;
wire  gpd ;
wire  GPD ;
wire  gpe ;
wire  GPE ;
wire  gpf ;
wire  GPF ;
wire  gpg ;
wire  GPG ;
wire  gph ;
wire  GPH ;
wire  gpi ;
wire  GPI ;
wire  gqa ;
wire  GQA ;
wire  gqb ;
wire  GQB ;
wire  gqc ;
wire  GQC ;
wire  gqd ;
wire  GQD ;
wire  gqe ;
wire  GQE ;
wire  gqf ;
wire  GQF ;
wire  gqg ;
wire  GQG ;
wire  gqh ;
wire  GQH ;
wire  gra ;
wire  GRA ;
wire  grb ;
wire  GRB ;
wire  grc ;
wire  GRC ;
wire  grd ;
wire  GRD ;
wire  gre ;
wire  GRE ;
wire  grf ;
wire  GRF ;
wire  grg ;
wire  GRG ;
wire  grh ;
wire  GRH ;
wire  haa ;
wire  hab ;
wire  hac ;
wire  had ;
wire  hae ;
wire  HAE ;
wire  haf ;
wire  hag ;
wire  hah ;
wire  hai ;
wire  HBA ;
wire  HBB ;
wire  HBC ;
wire  HBD ;
wire  hbe ;
wire  HBE ;
wire  HBF ;
wire  HBG ;
wire  hca ;
wire  hcb ;
wire  hcc ;
wire  hcd ;
wire  hce ;
wire  hcf ;
wire  HDA ;
wire  HDB ;
wire  HDC ;
wire  HDD ;
wire  HDE ;
wire  hea ;
wire  heb ;
wire  hec ;
wire  hed ;
wire  hee ;
wire  hef ;
wire  heg ;
wire  heh ;
wire  HFA ;
wire  HFB ;
wire  HFC ;
wire  HFD ;
wire  HFE ;
wire  HFF ;
wire  hga ;
wire  hgb ;
wire  hgc ;
wire  hgd ;
wire  hge ;
wire  hgf ;
wire  hgg ;
wire  HHA ;
wire  HHB ;
wire  HHC ;
wire  HHD ;
wire  HHE ;
wire  HHF ;
wire  HHG ;
wire  hia ;
wire  hib ;
wire  hic ;
wire  hid ;
wire  hie ;
wire  hif ;
wire  hig ;
wire  HJA ;
wire  HJB ;
wire  HJC ;
wire  HJD ;
wire  HJE ;
wire  HJF ;
wire  HJG ;
wire  hka ;
wire  hkb ;
wire  hkc ;
wire  hkd ;
wire  hke ;
wire  hkf ;
wire  hkg ;
wire  HLA ;
wire  HLB ;
wire  HLC ;
wire  HLD ;
wire  HLE ;
wire  HLF ;
wire  hma ;
wire  hmb ;
wire  hmc ;
wire  hmd ;
wire  hme ;
wire  hmf ;
wire  hmg ;
wire  hmh ;
wire  HNA ;
wire  HNB ;
wire  HNC ;
wire  HND ;
wire  HNE ;
wire  HNF ;
wire  hoa ;
wire  hob ;
wire  hoc ;
wire  hod ;
wire  hoe ;
wire  hof ;
wire  HPA ;
wire  HPB ;
wire  HPC ;
wire  HPD ;
wire  HPE ;
wire  HPF ;
wire  hqa ;
wire  hqb ;
wire  hqc ;
wire  hqd ;
wire  hqe ;
wire  hqf ;
wire  hqg ;
wire  iba ;
wire  ibb ;
wire  ibc ;
wire  ibd ;
wire  ibe ;
wire  ibf ;
wire  ibg ;
wire  ibh ;
wire  ibi ;
wire  ibj ;
wire  ibk ;
wire  ibl ;
wire  ibm ;
wire  ibn ;
wire  ibo ;
wire  ibp ;
wire  ica ;
wire  icb ;
wire  icc ;
wire  icd ;
wire  ice ;
wire  icf ;
wire  icg ;
wire  ich ;
wire  ici ;
wire  icj ;
wire  ick ;
wire  icl ;
wire  icm ;
wire  icn ;
wire  ico ;
wire  icp ;
wire  ida ;
wire  idb ;
wire  idc ;
wire  idd ;
wire  ide ;
wire  idf ;
wire  idg ;
wire  idh ;
wire  idi ;
wire  idj ;
wire  idk ;
wire  idl ;
wire  idm ;
wire  idn ;
wire  ido ;
wire  idp ;
wire  iea ;
wire  ieb ;
wire  iec ;
wire  ied ;
wire  iee ;
wire  ief ;
wire  ieg ;
wire  ieh ;
wire  iei ;
wire  iej ;
wire  iek ;
wire  iel ;
wire  iem ;
wire  ien ;
wire  ieo ;
wire  iep ;
wire  ieq ;
wire  ier ;
wire  ies ;
wire  iet ;
wire  ieu ;
wire  iev ;
wire  iew ;
wire  iex ;
wire  iey ;
wire  iez ;
wire  ifa ;
wire  ifb ;
wire  ifc ;
wire  ifd ;
wire  ife ;
wire  ifff  ;
wire  ifg ;
wire  ifh ;
wire  ifi ;
wire  ifj ;
wire  ifk ;
wire  ifl ;
wire  ifm ;
wire  ifn ;
wire  ifo ;
wire  ifp ;
wire  iga ;
wire  igb ;
wire  igc ;
wire  igd ;
wire  ige ;
wire  igf ;
wire  igg ;
wire  igh ;
wire  igi ;
wire  igj ;
wire  igk ;
wire  igl ;
wire  igm ;
wire  ign ;
wire  igo ;
wire  igp ;
wire  iha ;
wire  iia ;
wire  ika ;
wire  ila ;
wire  ilb ;
wire  ilc ;
wire  ild ;
wire  ile ;
wire  ilf ;
wire  ilg ;
wire  ilh ;
wire  ili ;
wire  ilj ;
wire  ilk ;
wire  ill ;
wire  ilm ;
wire  iln ;
wire  ilo ;
wire  ilp ;
wire  ima ;
wire  imb ;
wire  imc ;
wire  imd ;
wire  ime ;
wire  imf ;
wire  img ;
wire  imh ;
wire  imi ;
wire  imj ;
wire  imk ;
wire  iml ;
wire  imm ;
wire  imn ;
wire  ina ;
wire  inb ;
wire  inc ;
wire  ind ;
wire  ine ;
wire  inf ;
wire  ing ;
wire  ioa ;
wire  iob ;
wire  ioc ;
wire  ira ;
wire  isa ;
wire  ita ;
wire  itb ;
wire  jaa ;
wire  JAA ;
wire  jab ;
wire  JAB ;
wire  jac ;
wire  JAC ;
wire  jba ;
wire  JBA ;
wire  jbb ;
wire  JBB ;
wire  jbc ;
wire  JBC ;
wire  jca ;
wire  JCA ;
wire  jcb ;
wire  JCB ;
wire  jcc ;
wire  JCC ;
wire  jcd ;
wire  JCD ;
wire  jda ;
wire  JDA ;
wire  jdb ;
wire  JDB ;
wire  jdc ;
wire  JDC ;
wire  jdd ;
wire  JDD ;
wire  jea ;
wire  JEA ;
wire  jeb ;
wire  JEB ;
wire  jec ;
wire  JEC ;
wire  jed ;
wire  JED ;
wire  jfa ;
wire  JFA ;
wire  jfb ;
wire  JFB ;
wire  jfc ;
wire  JFC ;
wire  jfd ;
wire  JFD ;
wire  jga ;
wire  JGA ;
wire  jgb ;
wire  JGB ;
wire  jgc ;
wire  JGC ;
wire  jgd ;
wire  JGD ;
wire  jha ;
wire  JHA ;
wire  jhb ;
wire  JHB ;
wire  jhc ;
wire  JHC ;
wire  jhd ;
wire  JHD ;
wire  jia ;
wire  JIA ;
wire  jib ;
wire  JIB ;
wire  jic ;
wire  JIC ;
wire  jid ;
wire  JID ;
wire  jja ;
wire  JJA ;
wire  jjb ;
wire  JJB ;
wire  jjc ;
wire  JJC ;
wire  jjd ;
wire  JJD ;
wire  jka ;
wire  JKA ;
wire  jkb ;
wire  JKB ;
wire  jkc ;
wire  JKC ;
wire  jkd ;
wire  JKD ;
wire  jla ;
wire  JLA ;
wire  jlb ;
wire  JLB ;
wire  jlc ;
wire  JLC ;
wire  jld ;
wire  JLD ;
wire  jma ;
wire  JMA ;
wire  jmb ;
wire  JMB ;
wire  jmc ;
wire  JMC ;
wire  jmd ;
wire  JMD ;
wire  jna ;
wire  JNA ;
wire  jnb ;
wire  JNB ;
wire  jnc ;
wire  JNC ;
wire  jnd ;
wire  JND ;
wire  joa ;
wire  JOA ;
wire  job ;
wire  JOB ;
wire  joc ;
wire  JOC ;
wire  jod ;
wire  JOD ;
wire  jpa ;
wire  JPA ;
wire  jpb ;
wire  JPB ;
wire  jpc ;
wire  JPC ;
wire  jpd ;
wire  JPD ;
wire  jqa ;
wire  JQA ;
wire  jqb ;
wire  JQB ;
wire  jqc ;
wire  JQC ;
wire  jqd ;
wire  JQD ;
wire  jra ;
wire  JRA ;
wire  jrb ;
wire  JRB ;
wire  jrc ;
wire  JRC ;
wire  jrd ;
wire  JRD ;
wire  kaa ;
wire  kab ;
wire  kac ;
wire  kad ;
wire  kae ;
wire  kaf ;
wire  KBA ;
wire  KBB ;
wire  KBC ;
wire  KBD ;
wire  kca ;
wire  kcb ;
wire  kcc ;
wire  kcd ;
wire  kce ;
wire  KDA ;
wire  KDB ;
wire  KDC ;
wire  kea ;
wire  keb ;
wire  kec ;
wire  KFA ;
wire  KFB ;
wire  KFC ;
wire  kga ;
wire  kgb ;
wire  kgc ;
wire  KHA ;
wire  KHB ;
wire  KHC ;
wire  kia ;
wire  kib ;
wire  kic ;
wire  kid ;
wire  KJA ;
wire  KJB ;
wire  KJC ;
wire  kka ;
wire  kkb ;
wire  kkc ;
wire  kkd ;
wire  KLA ;
wire  KLB ;
wire  KLC ;
wire  kma ;
wire  kmb ;
wire  kmc ;
wire  kmd ;
wire  KNA ;
wire  KNB ;
wire  KNC ;
wire  koa ;
wire  kob ;
wire  koc ;
wire  kod ;
wire  KPA ;
wire  KPB ;
wire  kqa ;
wire  kqb ;
wire  kqc ;
wire  laa ;
wire  LAA ;
wire  lab ;
wire  LAB ;
wire  lba ;
wire  LBA ;
wire  lbb ;
wire  LBB ;
wire  lca ;
wire  LCA ;
wire  lcb ;
wire  LCB ;
wire  lcc ;
wire  LCC ;
wire  lda ;
wire  LDA ;
wire  ldb ;
wire  LDB ;
wire  ldc ;
wire  LDC ;
wire  lea ;
wire  LEA ;
wire  leb ;
wire  LEB ;
wire  lfa ;
wire  LFA ;
wire  lfb ;
wire  LFB ;
wire  lga ;
wire  LGA ;
wire  lgb ;
wire  LGB ;
wire  lha ;
wire  LHA ;
wire  lhb ;
wire  LHB ;
wire  lia ;
wire  LIA ;
wire  lib ;
wire  LIB ;
wire  lja ;
wire  LJA ;
wire  ljb ;
wire  LJB ;
wire  lka ;
wire  LKA ;
wire  lkb ;
wire  LKB ;
wire  lla ;
wire  LLA ;
wire  llb ;
wire  LLB ;
wire  lma ;
wire  LMA ;
wire  lmb ;
wire  LMB ;
wire  lna ;
wire  LNA ;
wire  lnb ;
wire  LNB ;
wire  loa ;
wire  LOA ;
wire  lob ;
wire  LOB ;
wire  lpa ;
wire  LPA ;
wire  lpb ;
wire  LPB ;
wire  lqa ;
wire  LQA ;
wire  lra ;
wire  LRA ;
wire  maa ;
wire  mab ;
wire  mac ;
wire  mad ;
wire  MBA ;
wire  MBB ;
wire  mca ;
wire  mcb ;
wire  MDA ;
wire  MDB ;
wire  mea ;
wire  meb ;
wire  mec ;
wire  MFA ;
wire  mga ;
wire  mgb ;
wire  MHA ;
wire  mia ;
wire  mib ;
wire  mic ;
wire  MJA ;
wire  mka ;
wire  mkb ;
wire  mkc ;
wire  MLA ;
wire  mma ;
wire  mmb ;
wire  mmc ;
wire  MNA ;
wire  moa ;
wire  mob ;
wire  moc ;
wire  MPA ;
wire  mqa ;
wire  mqb ;
wire  mqc ;
wire  naa ;
wire  NAA ;
wire  nba ;
wire  NBA ;
wire  nca ;
wire  NCA ;
wire  nda ;
wire  NDA ;
wire  nea ;
wire  NEA ;
wire  nfa ;
wire  NFA ;
wire  nga ;
wire  NGA ;
wire  nha ;
wire  NHA ;
wire  nia ;
wire  NIA ;
wire  nja ;
wire  NJA ;
wire  nka ;
wire  NKA ;
wire  nla ;
wire  NLA ;
wire  nma ;
wire  NMA ;
wire  nna ;
wire  NNA ;
wire  noa ;
wire  NOA ;
wire  npa ;
wire  NPA ;
wire  nqa ;
wire  NQA ;
wire  nra ;
wire  NRA ;
wire  oaa ;
wire  oab ;
wire  oac ;
wire  oad ;
wire  oae ;
wire  oaf ;
wire  oag ;
wire  oah ;
wire  oai ;
wire  oaj ;
wire  oak ;
wire  oal ;
wire  oam ;
wire  oan ;
wire  oao ;
wire  oap ;
wire  oba ;
wire  obb ;
wire  obc ;
wire  obd ;
wire  obe ;
wire  obf ;
wire  obg ;
wire  obh ;
wire  obi ;
wire  obj ;
wire  obk ;
wire  obl ;
wire  obm ;
wire  obn ;
wire  obo ;
wire  obp ;
wire  OCA ;
wire  OCB ;
wire  OCC ;
wire  OCD ;
wire  OCE ;
wire  OCF ;
wire  OCG ;
wire  OCH ;
wire  OCI ;
wire  OCJ ;
wire  OCK ;
wire  OCL ;
wire  OCM ;
wire  OCN ;
wire  OCO ;
wire  OCP ;
wire  ODA ;
wire  ODB ;
wire  ODC ;
wire  ODD ;
wire  ODE ;
wire  ODF ;
wire  ODG ;
wire  ODH ;
wire  ODI ;
wire  ODJ ;
wire  ODK ;
wire  ODL ;
wire  ODM ;
wire  ODN ;
wire  ODO ;
wire  ODP ;
wire  OGA ;
wire  OGB ;
wire  OGC ;
wire  OGD ;
wire  OGE ;
wire  OGF ;
wire  OGG ;
wire  OGH ;
wire  OGI ;
wire  OGJ ;
wire  OGK ;
wire  OGL ;
wire  OGM ;
wire  OHA ;
wire  OHB ;
wire  OHC ;
wire  OHD ;
wire  OHE ;
wire  OHF ;
wire  ohg ;
wire  ohh ;
wire  ohi ;
wire  ohj ;
wire  OIG ;
wire  OIH ;
wire  OKA ;
wire  OKB ;
wire  OKC ;
wire  okd ;
wire  oke ;
wire  OLD ;
wire  OMA ;
wire  omb ;
wire  opa ;
wire  opb ;
wire  opc ;
wire  opd ;
wire  ope ;
wire  opf ;
wire  opg ;
wire  oph ;
wire  opi ;
wire  opk ;
wire  opm ;
wire  opo ;
wire  opq ;
wire  opr ;
wire  OQA ;
wire  OQC ;
wire  OQE ;
wire  OQI ;
wire  OQK ;
wire  OQM ;
wire  OQO ;
wire  OQQ ;
wire  qaa ;
wire  qga ;
wire  qha ;
wire  qia ;
wire  qib ;
wire  qic ;
wire  qid ;
wire  qie ;
wire  qka ;
wire  qta ;
wire  qtb ;
wire  tga ;
wire  tgb ;
wire  tgc ;
wire  tha ;
wire  thb ;
wire  thc ;
wire  thd ;
wire  the ;
wire  thf ;
wire  tka ;
wire  tkb ;
wire  tkc ;
wire  tkd ;
wire  tke ;
wire  tkf ;
wire  tra ;
wire  trb ;
wire  tsa ;
wire  tsb ;
wire  tsc ;
wire  tsd ;
wire  tse ;
wire  tsf ;
wire  tta ;
wire  ttb ;
wire  ttc ;
wire  ZZI ;
wire  ZZO ;
assign ZZI = 1'b1;
assign ZZO = 1'b0;
assign fae = ~FAE;  //complement 
assign FBE = ~fbe;  //complement 
assign faf = ~FAF;  //complement 
assign FBF = ~fbf;  //complement 
assign fag = ~FAG;  //complement 
assign FBG = ~fbg;  //complement 
assign fah = ~FAH;  //complement 
assign FBH = ~fbh;  //complement 
assign aab = ~AAB;  //complement 
assign fab = ~FAB;  //complement 
assign FBB = ~fbb;  //complement 
assign fac = ~FAC;  //complement 
assign FBC = ~fbc;  //complement 
assign fad = ~FAD;  //complement 
assign FBD = ~fbd;  //complement 
assign fcd = ~FCD;  //complement 
assign FDD = ~fdd;  //complement 
assign fce = ~FCE;  //complement 
assign FDE = ~fde;  //complement 
assign fcf = ~FCF;  //complement 
assign FDF = ~fdf;  //complement 
assign fcg = ~FCG;  //complement 
assign FDG = ~fdg;  //complement 
assign aac = ~AAC;  //complement 
assign fca = ~FCA;  //complement 
assign FDA = ~fda;  //complement 
assign fcb = ~FCB;  //complement 
assign FDB = ~fdb;  //complement 
assign fcc = ~FCC;  //complement 
assign FDC = ~fdc;  //complement 
assign aad = ~AAD;  //complement 
assign aae = ~AAE;  //complement 
assign aaf = ~AAF;  //complement 
assign aag = ~AAG;  //complement 
assign fec = ~FEC;  //complement 
assign FFC = ~ffc;  //complement 
assign fed = ~FED;  //complement 
assign FFD = ~ffd;  //complement 
assign fee = ~FEE;  //complement 
assign FFE = ~ffe;  //complement 
assign fef = ~FEF;  //complement 
assign FFF = ~fff;  //complement 
assign ODA = ~oda;  //complement 
assign ODB = ~odb;  //complement 
assign ODC = ~odc;  //complement 
assign ODD = ~odd;  //complement 
assign ODE = ~ode;  //complement 
assign ODF = ~odf;  //complement 
assign ODG = ~odg;  //complement 
assign ODH = ~odh;  //complement 
assign fea = ~FEA;  //complement 
assign FFA = ~ffa;  //complement 
assign feb = ~FEB;  //complement 
assign FFB = ~ffb;  //complement 
assign ODI = ~odi;  //complement 
assign ODJ = ~odj;  //complement 
assign ODK = ~odk;  //complement 
assign ODL = ~odl;  //complement 
assign ODM = ~odm;  //complement 
assign ODN = ~odn;  //complement 
assign ODO = ~odo;  //complement 
assign ODP = ~odp;  //complement 
assign aaa = ~AAA;  //complement 
assign fam = ~FAM;  //complement 
assign FBM = ~fbm;  //complement 
assign qha = ~QHA;  //complement 
assign tha = ~THA;  //complement 
assign thb = ~THB;  //complement 
assign thc = ~THC;  //complement 
assign fan = ~FAN;  //complement 
assign FBN = ~fbn;  //complement 
assign faq = ~FAQ;  //complement 
assign fao = ~FAO;  //complement 
assign FBO = ~fbo;  //complement 
assign fap = ~FAP;  //complement 
assign faj = ~FAJ;  //complement 
assign FBJ = ~fbj;  //complement 
assign thd = ~THD;  //complement 
assign the = ~THE;  //complement 
assign thf = ~THF;  //complement 
assign fak = ~FAK;  //complement 
assign FBK = ~fbk;  //complement 
assign fal = ~FAL;  //complement 
assign FBL = ~fbl;  //complement 
assign fcn = ~FCN;  //complement 
assign FDN = ~fdn;  //complement 
assign fco = ~FCO;  //complement 
assign FDO = ~fdo;  //complement 
assign fcp = ~FCP;  //complement 
assign faa = ~FAA;  //complement 
assign FBA = ~fba;  //complement 
assign fai = ~FAI;  //complement 
assign FBI = ~fbi;  //complement 
assign fck = ~FCK;  //complement 
assign FDK = ~fdk;  //complement 
assign fcl = ~FCL;  //complement 
assign FDL = ~fdl;  //complement 
assign fcm = ~FCM;  //complement 
assign FDM = ~fdm;  //complement 
assign fch = ~FCH;  //complement 
assign FDH = ~fdh;  //complement 
assign fci = ~FCI;  //complement 
assign FDI = ~fdi;  //complement 
assign fcj = ~FCJ;  //complement 
assign FDJ = ~fdj;  //complement 
assign fem = ~FEM;  //complement 
assign FFM = ~ffm;  //complement 
assign tsa = ~TSA;  //complement 
assign tsb = ~TSB;  //complement 
assign tsc = ~TSC;  //complement 
assign tsd = ~TSD;  //complement 
assign fen = ~FEN;  //complement 
assign FFN = ~ffn;  //complement 
assign feo = ~FEO;  //complement 
assign FFO = ~ffo;  //complement 
assign fej = ~FEJ;  //complement 
assign FFJ = ~ffj;  //complement 
assign tra = ~TRA;  //complement 
assign trb = ~TRB;  //complement 
assign qtb = ~QTB;  //complement 
assign fek = ~FEK;  //complement 
assign FFK = ~ffk;  //complement 
assign fel = ~FEL;  //complement 
assign FFL = ~ffl;  //complement 
assign feg = ~FEG;  //complement 
assign FFG = ~ffg;  //complement 
assign mqc = ~MQC;  //complement 
assign moc = ~MOC;  //complement 
assign mmc = ~MMC;  //complement 
assign omb = ~OMB;  //complement 
assign feh = ~FEH;  //complement 
assign FFH = ~ffh;  //complement 
assign fei = ~FEI;  //complement 
assign FFI = ~ffi;  //complement 
assign ERI =  CBJ & DFA  ; 
assign eri = ~ERI;  //complement 
assign EMJ =  CCO & DGJ  ; 
assign emj = ~EMJ;  //complement 
assign dha = ~DHA;  //complement 
assign dhb = ~DHB;  //complement 
assign dhc = ~DHC;  //complement 
assign dhd = ~DHD;  //complement 
assign cac = ~CAC;  //complement 
assign cdc = ~CDC;  //complement 
assign cad = ~CAD;  //complement 
assign cdd = ~CDD;  //complement 
assign EMI =  CCP & DGI  ; 
assign emi = ~EMI;  //complement 
assign EOJ =  CCP & DGJ  ; 
assign eoj = ~EOJ;  //complement 
assign EBX =  CAC & DCP  ; 
assign ebx = ~EBX;  //complement 
assign EBW =  CAD & DCO  ; 
assign ebw = ~EBW;  //complement 
assign EDX =  CAD & DCP  ; 
assign edx = ~EDX;  //complement 
assign dhe = ~DHE;  //complement 
assign dhf = ~DHF;  //complement 
assign dhg = ~DHG;  //complement 
assign dhh = ~DHH;  //complement 
assign cae = ~CAE;  //complement 
assign cde = ~CDE;  //complement 
assign cah = ~CAH;  //complement 
assign qaa = ~QAA;  //complement 
assign EDW =  CAE & DCO  ; 
assign edw = ~EDW;  //complement 
assign ELV =  CAJ & DCN  ; 
assign elv = ~ELV;  //complement 
assign ELU =  CAK & DCM  ; 
assign elu = ~ELU;  //complement 
assign ENV =  CAK & DCN  ; 
assign env = ~ENV;  //complement 
assign ELT =  CAL & DCL  ; 
assign elt = ~ELT;  //complement 
assign ENU =  CAL & DCM  ; 
assign enu = ~ENU;  //complement 
assign dhi = ~DHI;  //complement 
assign dhj = ~DHJ;  //complement 
assign dhk = ~DHK;  //complement 
assign dhl = ~DHL;  //complement 
assign cag = ~CAG;  //complement 
assign cdg = ~CDG;  //complement 
assign tse = ~TSE;  //complement 
assign ELS =  CAM & DCK  ; 
assign els = ~ELS;  //complement 
assign ENT =  CAM & DCL  ; 
assign ent = ~ENT;  //complement 
assign ELR =  CAN & DCJ  ; 
assign elr = ~ELR;  //complement 
assign ENS =  CAN & DCK  ; 
assign ens = ~ENS;  //complement 
assign ELQ =  CAO & DCI  ; 
assign elq = ~ELQ;  //complement 
assign ENR =  CAO & DCJ  ; 
assign enr = ~ENR;  //complement 
assign dga = ~DGA;  //complement 
assign dgb = ~DGB;  //complement 
assign dgc = ~DGC;  //complement 
assign dgd = ~DGD;  //complement 
assign dac = ~DAC;  //complement 
assign dad = ~DAD;  //complement 
assign dae = ~DAE;  //complement 
assign daf = ~DAF;  //complement 
assign ELP =  CAP & DCH  ; 
assign elp = ~ELP;  //complement 
assign ENQ =  CAP & DCI  ; 
assign enq = ~ENQ;  //complement 
assign EBJ =  CBA & DCB  ; 
assign ebj = ~EBJ;  //complement 
assign ELO =  CBA & DCG  ; 
assign elo = ~ELO;  //complement 
assign ENP =  CBA & DCH  ; 
assign enp = ~ENP;  //complement 
assign ELN =  CBB & DCF  ; 
assign eln = ~ELN;  //complement 
assign dhm = ~DHM;  //complement 
assign dhn = ~DHN;  //complement 
assign dho = ~DHO;  //complement 
assign dhp = ~DHP;  //complement 
assign dah = ~DAH;  //complement 
assign DDH = ~ddh;  //complement 
assign dag = ~DAG;  //complement 
assign DDG = ~ddg;  //complement 
assign ENO =  CBB & DCG  ; 
assign eno = ~ENO;  //complement 
assign ELM =  CBC & DCE  ; 
assign elm = ~ELM;  //complement 
assign ENN =  CBC & DCF  ; 
assign enn = ~ENN;  //complement 
assign ELL =  CBD & DCD  ; 
assign ell = ~ELL;  //complement 
assign ENM =  CBD & DCE  ; 
assign enm = ~ENM;  //complement 
assign EHJ =  CBD & DFB  ; 
assign ehj = ~EHJ;  //complement 
assign DDF = ~ddf;  //complement 
assign cdh = ~CDH;  //complement 
assign tsf = ~TSF;  //complement 
assign dai = ~DAI;  //complement 
assign DDI = ~ddi;  //complement 
assign daj = ~DAJ;  //complement 
assign DDJ = ~ddj;  //complement 
assign ELK =  CBE & DCC  ; 
assign elk = ~ELK;  //complement 
assign ENL =  CBE & DCD  ; 
assign enl = ~ENL;  //complement 
assign EIU =  CCB & DBE  ; 
assign eiu = ~EIU;  //complement 
assign ENK =  CBF & DCC  ; 
assign enk = ~ENK;  //complement 
assign EHH =  CBF & DEP  ; 
assign ehh = ~EHH;  //complement 
assign mkc = ~MKC;  //complement 
assign mic = ~MIC;  //complement 
assign meb = ~MEB;  //complement 
assign mec = ~MEC;  //complement 
assign dak = ~DAK;  //complement 
assign DDK = ~ddk;  //complement 
assign dal = ~DAL;  //complement 
assign DDL = ~ddl;  //complement 
assign ELI =  CBG & DCA  ; 
assign eli = ~ELI;  //complement 
assign ENJ =  CBG & DCB  ; 
assign enj = ~ENJ;  //complement 
assign EHG =  CBG & DEO  ; 
assign ehg = ~EHG;  //complement 
assign ELH =  CBH & DBP  ; 
assign elh = ~ELH;  //complement 
assign ENI =  CBH & DCA  ; 
assign eni = ~ENI;  //complement 
assign EHF =  CBH & DEN  ; 
assign ehf = ~EHF;  //complement 
assign dao = ~DAO;  //complement 
assign DDO = ~ddo;  //complement 
assign dap = ~DAP;  //complement 
assign DDP = ~ddp;  //complement 
assign dam = ~DAM;  //complement 
assign DDM = ~ddm;  //complement 
assign dan = ~DAN;  //complement 
assign DDN = ~ddn;  //complement 
assign fgb = ~FGB;  //complement 
assign FHB = ~fhb;  //complement 
assign fgc = ~FGC;  //complement 
assign FHC = ~fhc;  //complement 
assign fgd = ~FGD;  //complement 
assign FHD = ~fhd;  //complement 
assign fge = ~FGE;  //complement 
assign FHE = ~fhe;  //complement 
assign fic = ~FIC;  //complement 
assign FJC = ~fjc;  //complement 
assign fid = ~FID;  //complement 
assign FJD = ~fjd;  //complement 
assign fie = ~FIE;  //complement 
assign FJE = ~fje;  //complement 
assign fga = ~FGA;  //complement 
assign FHA = ~fha;  //complement 
assign fib = ~FIB;  //complement 
assign FJB = ~fjb;  //complement 
assign fkh = ~FKH;  //complement 
assign FLH = ~flh;  //complement 
assign fia = ~FIA;  //complement 
assign FJA = ~fja;  //complement 
assign fkg = ~FKG;  //complement 
assign FLG = ~flg;  //complement 
assign aal = ~AAL;  //complement 
assign fkc = ~FKC;  //complement 
assign FLC = ~flc;  //complement 
assign fkd = ~FKD;  //complement 
assign FLD = ~fld;  //complement 
assign fke = ~FKE;  //complement 
assign FLE = ~fle;  //complement 
assign fkf = ~FKF;  //complement 
assign FLF = ~flf;  //complement 
assign aam = ~AAM;  //complement 
assign aan = ~AAN;  //complement 
assign fka = ~FKA;  //complement 
assign FLA = ~fla;  //complement 
assign fkb = ~FKB;  //complement 
assign FLB = ~flb;  //complement 
assign OCA = ~oca;  //complement 
assign OCB = ~ocb;  //complement 
assign OCC = ~occ;  //complement 
assign OCD = ~ocd;  //complement 
assign OCE = ~oce;  //complement 
assign OCF = ~ocf;  //complement 
assign OCG = ~ocg;  //complement 
assign OCH = ~och;  //complement 
assign OCI = ~oci;  //complement 
assign OCJ = ~ocj;  //complement 
assign OCK = ~ock;  //complement 
assign OCL = ~ocl;  //complement 
assign OCM = ~ocm;  //complement 
assign OCN = ~ocn;  //complement 
assign OCO = ~oco;  //complement 
assign OCP = ~ocp;  //complement 
assign aah = ~AAH;  //complement 
assign aai = ~AAI;  //complement 
assign aaj = ~AAJ;  //complement 
assign aak = ~AAK;  //complement 
assign fgl = ~FGL;  //complement 
assign FHL = ~fhl;  //complement 
assign fgp = ~FGP;  //complement 
assign fgm = ~FGM;  //complement 
assign FHM = ~fhm;  //complement 
assign fgo = ~FGO;  //complement 
assign fgn = ~FGN;  //complement 
assign FHN = ~fhn;  //complement 
assign fgi = ~FGI;  //complement 
assign FHI = ~fhi;  //complement 
assign fgj = ~FGJ;  //complement 
assign FHJ = ~fhj;  //complement 
assign fgk = ~FGK;  //complement 
assign FHK = ~fhk;  //complement 
assign fgf = ~FGF;  //complement 
assign FHF = ~fhf;  //complement 
assign fgg = ~FGG;  //complement 
assign FHG = ~fhg;  //complement 
assign fgh = ~FGH;  //complement 
assign FHH = ~fhh;  //complement 
assign fil = ~FIL;  //complement 
assign FJL = ~fjl;  //complement 
assign fim = ~FIM;  //complement 
assign FJM = ~fjm;  //complement 
assign fin = ~FIN;  //complement 
assign FJN = ~fjn;  //complement 
assign fio = ~FIO;  //complement 
assign fii = ~FII;  //complement 
assign FJI = ~fji;  //complement 
assign fij = ~FIJ;  //complement 
assign FJJ = ~fjj;  //complement 
assign fik = ~FIK;  //complement 
assign FJK = ~fjk;  //complement 
assign fif = ~FIF;  //complement 
assign FJF = ~fjf;  //complement 
assign fig = ~FIG;  //complement 
assign FJG = ~fjg;  //complement 
assign fih = ~FIH;  //complement 
assign FJH = ~fjh;  //complement 
assign fkl = ~FKL;  //complement 
assign FLL = ~fll;  //complement 
assign qie = ~QIE;  //complement 
assign fkm = ~FKM;  //complement 
assign FLM = ~flm;  //complement 
assign fkn = ~FKN;  //complement 
assign FLN = ~fln;  //complement 
assign fki = ~FKI;  //complement 
assign FLI = ~fli;  //complement 
assign qia = ~QIA;  //complement 
assign qib = ~QIB;  //complement 
assign qic = ~QIC;  //complement 
assign qid = ~QID;  //complement 
assign fkj = ~FKJ;  //complement 
assign FLJ = ~flj;  //complement 
assign fkk = ~FKK;  //complement 
assign FLK = ~flk;  //complement 
assign EPJ =  CBH & DFB  ; 
assign epj = ~EPJ;  //complement 
assign ELG =  CBI & DBO  ; 
assign elg = ~ELG;  //complement 
assign EHE =  CBI & DEM  ; 
assign ehe = ~EHE;  //complement 
assign EPI =  CBI & DFA  ; 
assign epi = ~EPI;  //complement 
assign ERJ =  CBI & DFB  ; 
assign erj = ~ERJ;  //complement 
assign ELF =  CBJ & DBN  ; 
assign elf = ~ELF;  //complement 
assign cai = ~CAI;  //complement 
assign cdi = ~CDI;  //complement 
assign caj = ~CAJ;  //complement 
assign cdj = ~CDJ;  //complement 
assign EHD =  CBJ & DEL  ; 
assign ehd = ~EHD;  //complement 
assign ELE =  CBK & DBM  ; 
assign ele = ~ELE;  //complement 
assign EHC =  CBK & DEK  ; 
assign ehc = ~EHC;  //complement 
assign ELD =  CBL & DBL  ; 
assign eld = ~ELD;  //complement 
assign EHB =  CBL & DEJ  ; 
assign ehb = ~EHB;  //complement 
assign ELC =  CBM & DBK  ; 
assign elc = ~ELC;  //complement 
assign cak = ~CAK;  //complement 
assign cdk = ~CDK;  //complement 
assign cal = ~CAL;  //complement 
assign cdl = ~CDL;  //complement 
assign EHA =  CBM & DEI  ; 
assign eha = ~EHA;  //complement 
assign ELB =  CBN & DBJ  ; 
assign elb = ~ELB;  //complement 
assign EGX =  CBN & DEH  ; 
assign egx = ~EGX;  //complement 
assign ELA =  CBO & DBI  ; 
assign ela = ~ELA;  //complement 
assign EGW =  CBO & DEG  ; 
assign egw = ~EGW;  //complement 
assign cam = ~CAM;  //complement 
assign cdm = ~CDM;  //complement 
assign can = ~CAN;  //complement 
assign cdn = ~CDN;  //complement 
assign EKX =  CBP & DBH  ; 
assign ekx = ~EKX;  //complement 
assign EGV =  CBP & DEF  ; 
assign egv = ~EGV;  //complement 
assign EKW =  CCA & DBG  ; 
assign ekw = ~EKW;  //complement 
assign EGU =  CCA & DEE  ; 
assign egu = ~EGU;  //complement 
assign EKV =  CCB & DBF  ; 
assign ekv = ~EKV;  //complement 
assign EGT =  CCB & DED  ; 
assign egt = ~EGT;  //complement 
assign dba = ~DBA;  //complement 
assign DEA = ~dea;  //complement 
assign dbb = ~DBB;  //complement 
assign DEB = ~deb;  //complement 
assign EKU =  CCC & DBE  ; 
assign eku = ~EKU;  //complement 
assign EGS =  CCC & DEC  ; 
assign egs = ~EGS;  //complement 
assign EKT =  CCD & DBD  ; 
assign ekt = ~EKT;  //complement 
assign EGR =  CCD & DEB  ; 
assign egr = ~EGR;  //complement 
assign dbc = ~DBC;  //complement 
assign DEC = ~dec;  //complement 
assign dbd = ~DBD;  //complement 
assign DED = ~ded;  //complement 
assign EIR =  CCE & DBB  ; 
assign eir = ~EIR;  //complement 
assign EKS =  CCE & DBC  ; 
assign eks = ~EKS;  //complement 
assign EGQ =  CCE & DEA  ; 
assign egq = ~EGQ;  //complement 
assign EKR =  CCF & DBB  ; 
assign ekr = ~EKR;  //complement 
assign EGP =  CCF & DDP  ; 
assign egp = ~EGP;  //complement 
assign dgi = ~DGI;  //complement 
assign dgj = ~DGJ;  //complement 
assign dgk = ~DGK;  //complement 
assign dgl = ~DGL;  //complement 
assign dbe = ~DBE;  //complement 
assign DEE = ~dee;  //complement 
assign dbf = ~DBF;  //complement 
assign DEF = ~def;  //complement 
assign dge = ~DGE;  //complement 
assign dgf = ~DGF;  //complement 
assign dgg = ~DGG;  //complement 
assign dgh = ~DGH;  //complement 
assign dbg = ~DBG;  //complement 
assign DEG = ~deg;  //complement 
assign dbh = ~DBH;  //complement 
assign DEH = ~deh;  //complement 
assign fql = ~FQL;  //complement 
assign OGL = ~ogl;  //complement 
assign fqm = ~FQM;  //complement 
assign OGM = ~ogm;  //complement 
assign foa = ~FOA;  //complement 
assign FPA = ~fpa;  //complement 
assign fob = ~FOB;  //complement 
assign FPB = ~fpb;  //complement 
assign fqh = ~FQH;  //complement 
assign OGH = ~ogh;  //complement 
assign fqi = ~FQI;  //complement 
assign OGI = ~ogi;  //complement 
assign fqj = ~FQJ;  //complement 
assign OGJ = ~ogj;  //complement 
assign fqk = ~FQK;  //complement 
assign OGK = ~ogk;  //complement 
assign fqd = ~FQD;  //complement 
assign OGD = ~ogd;  //complement 
assign fqe = ~FQE;  //complement 
assign OGE = ~oge;  //complement 
assign fqf = ~FQF;  //complement 
assign OGF = ~ogf;  //complement 
assign fqg = ~FQG;  //complement 
assign OGG = ~ogg;  //complement 
assign fqa = ~FQA;  //complement 
assign OGA = ~oga;  //complement 
assign bac = ~BAC;  //complement 
assign fqb = ~FQB;  //complement 
assign OGB = ~ogb;  //complement 
assign fqc = ~FQC;  //complement 
assign OGC = ~ogc;  //complement 
assign bad = ~BAD;  //complement 
assign bae = ~BAE;  //complement 
assign baf = ~BAF;  //complement 
assign bag = ~BAG;  //complement 
assign bah = ~BAH;  //complement 
assign bai = ~BAI;  //complement 
assign baj = ~BAJ;  //complement 
assign bak = ~BAK;  //complement 
assign aao = ~AAO;  //complement 
assign aap = ~AAP;  //complement 
assign baa = ~BAA;  //complement 
assign bab = ~BAB;  //complement 
assign fmk = ~FMK;  //complement 
assign FNK = ~fnk;  //complement 
assign fml = ~FML;  //complement 
assign FNL = ~fnl;  //complement 
assign fmo = ~FMO;  //complement 
assign fmm = ~FMM;  //complement 
assign FNM = ~fnm;  //complement 
assign fmn = ~FMN;  //complement 
assign fmh = ~FMH;  //complement 
assign FNH = ~fnh;  //complement 
assign fmi = ~FMI;  //complement 
assign FNI = ~fni;  //complement 
assign fmj = ~FMJ;  //complement 
assign FNJ = ~fnj;  //complement 
assign fme = ~FME;  //complement 
assign FNE = ~fne;  //complement 
assign fmf = ~FMF;  //complement 
assign FNF = ~fnf;  //complement 
assign fmg = ~FMG;  //complement 
assign FNG = ~fng;  //complement 
assign fmb = ~FMB;  //complement 
assign FNB = ~fnb;  //complement 
assign fmc = ~FMC;  //complement 
assign FNC = ~fnc;  //complement 
assign fmd = ~FMD;  //complement 
assign FND = ~fnd;  //complement 
assign fol = ~FOL;  //complement 
assign FPL = ~fpl;  //complement 
assign fom = ~FOM;  //complement 
assign FPM = ~fpm;  //complement 
assign fon = ~FON;  //complement 
assign fma = ~FMA;  //complement 
assign FNA = ~fna;  //complement 
assign foi = ~FOI;  //complement 
assign FPI = ~fpi;  //complement 
assign foj = ~FOJ;  //complement 
assign FPJ = ~fpj;  //complement 
assign fok = ~FOK;  //complement 
assign FPK = ~fpk;  //complement 
assign fof = ~FOF;  //complement 
assign FPF = ~fpf;  //complement 
assign fog = ~FOG;  //complement 
assign FPG = ~fpg;  //complement 
assign foh = ~FOH;  //complement 
assign FPH = ~fph;  //complement 
assign foc = ~FOC;  //complement 
assign FPC = ~fpc;  //complement 
assign fod = ~FOD;  //complement 
assign FPD = ~fpd;  //complement 
assign foe = ~FOE;  //complement 
assign FPE = ~fpe;  //complement 
assign EAL =  CCG & DAL  ; 
assign eal = ~EAL;  //complement 
assign EKQ =  CCG & DBA  ; 
assign ekq = ~EKQ;  //complement 
assign EGO =  CCG & DDO  ; 
assign ego = ~EGO;  //complement 
assign EKP =  CCH & DAP  ; 
assign ekp = ~EKP;  //complement 
assign EGN =  CCH & DDN  ; 
assign egn = ~EGN;  //complement 
assign bap = ~BAP;  //complement 
assign cao = ~CAO;  //complement 
assign cdo = ~CDO;  //complement 
assign caf = ~CAF;  //complement 
assign cdf = ~CDF;  //complement 
assign EKO =  CCI & DAO  ; 
assign eko = ~EKO;  //complement 
assign EGM =  CCI & DDM  ; 
assign egm = ~EGM;  //complement 
assign EGL =  CCJ & DDL  ; 
assign egl = ~EGL;  //complement 
assign EKM =  CCK & DAM  ; 
assign ekm = ~EKM;  //complement 
assign EGK =  CCK & DDK  ; 
assign egk = ~EGK;  //complement 
assign cap = ~CAP;  //complement 
assign cdp = ~CDP;  //complement 
assign cba = ~CBA;  //complement 
assign cea = ~CEA;  //complement 
assign cbb = ~CBB;  //complement 
assign ceb = ~CEB;  //complement 
assign EGJ =  CCL & DDJ  ; 
assign egj = ~EGJ;  //complement 
assign EAF =  CCM & DAF  ; 
assign eaf = ~EAF;  //complement 
assign EKK =  CCM & DAK  ; 
assign ekk = ~EKK;  //complement 
assign EGI =  CCM & DDI  ; 
assign egi = ~EGI;  //complement 
assign EAE =  CCN & DAE  ; 
assign eae = ~EAE;  //complement 
assign ECF =  CCN & DAF  ; 
assign ecf = ~ECF;  //complement 
assign cbc = ~CBC;  //complement 
assign cec = ~CEC;  //complement 
assign cbd = ~CBD;  //complement 
assign ced = ~CED;  //complement 
assign EKJ =  CCN & DAJ  ; 
assign ekj = ~EKJ;  //complement 
assign EGH =  CCN & DDH  ; 
assign egh = ~EGH;  //complement 
assign EAD =  CCO & DAD  ; 
assign ead = ~EAD;  //complement 
assign ECE =  CCO & DAE  ; 
assign ece = ~ECE;  //complement 
assign EEF =  CCO & DAF  ; 
assign eef = ~EEF;  //complement 
assign EKI =  CCO & DAI  ; 
assign eki = ~EKI;  //complement 
assign EGG =  CCO & DDG  ; 
assign egg = ~EGG;  //complement 
assign EAC =  CCP & DAC  ; 
assign eac = ~EAC;  //complement 
assign ECD =  CCP & DAD  ; 
assign ecd = ~ECD;  //complement 
assign EEE =  CCP & DAE  ; 
assign eee = ~EEE;  //complement 
assign EKH =  CCP & DAH  ; 
assign ekh = ~EKH;  //complement 
assign EGF =  CCP & DDF  ; 
assign egf = ~EGF;  //complement 
assign EIG =  CCP & DAG  ; 
assign eig = ~EIG;  //complement 
assign dbi = ~DBI;  //complement 
assign DEI = ~dei;  //complement 
assign dbj = ~DBJ;  //complement 
assign DEJ = ~dej;  //complement 
assign EAG =  CCL & DAG  ; 
assign eag = ~EAG;  //complement 
assign ECG =  CCM & DAG  ; 
assign ecg = ~ECG;  //complement 
assign EEG =  CCN & DAG  ; 
assign eeg = ~EEG;  //complement 
assign EAH = DAH & CCK ; 
assign eah = ~EAH ; //complement 
assign ECH = DAH & CCL ; 
assign ech = ~ECH ;  //complement 
assign EEH = DAH & CCM ; 
assign eeh = ~EEH ;  //complement 
assign EIH = DAH & CCO; 
assign eih = ~EIH; 
assign dgm = ~DGM;  //complement 
assign dgn = ~DGN;  //complement 
assign dgo = ~DGO;  //complement 
assign dgp = ~DGP;  //complement 
assign dbk = ~DBK;  //complement 
assign DEK = ~dek;  //complement 
assign dbl = ~DBL;  //complement 
assign DEL = ~del;  //complement 
assign EAI = DAI & CCJ ; 
assign eai = ~EAI ; //complement 
assign ECI = DAI & CCK ; 
assign eci = ~ECI ;  //complement 
assign EEI = DAI & CCL ; 
assign eei = ~EEI ;  //complement 
assign EII = DAI & CCN; 
assign eii = ~EII; 
assign EAJ = DAJ & CCI ; 
assign eaj = ~EAJ ; //complement 
assign ECJ = DAJ & CCJ ; 
assign ecj = ~ECJ ;  //complement 
assign EEJ = DAJ & CCK ; 
assign eej = ~EEJ ;  //complement 
assign EIJ = DAJ & CCM; 
assign eij = ~EIJ; 
assign bal = ~BAL;  //complement 
assign dbm = ~DBM;  //complement 
assign DEM = ~dem;  //complement 
assign dbn = ~DBN;  //complement 
assign DEN = ~den;  //complement 
assign bam = ~BAM;  //complement 
assign ban = ~BAN;  //complement 
assign bao = ~BAO;  //complement 
assign dbo = ~DBO;  //complement 
assign DEO = ~deo;  //complement 
assign dbp = ~DBP;  //complement 
assign DEP = ~dep;  //complement 
assign GEB =  FDD & fdl & fdh  |  fdd & FDL & fdh  |  fdd & fdl & FDH  |  FDD & FDL & FDH  ; 
assign geb = ~GEB; //complement 
assign gfb =  FDD & fdl & fdh  |  fdd & FDL & fdh  |  fdd & fdl & FDH  |  fdd & fdl & fdh  ; 
assign GFB = ~gfb;  //complement 
assign GEH =  FDC & fdj & fdn  |  fdc & FDJ & fdn  |  fdc & fdj & FDN  |  FDC & FDJ & FDN  ; 
assign geh = ~GEH; //complement 
assign gfh =  FDC & fdj & fdn  |  fdc & FDJ & fdn  |  fdc & fdj & FDN  |  fdc & fdj & fdn  ; 
assign GFH = ~gfh;  //complement 
assign GED =  FDA & fde & fdm  |  fda & FDE & fdm  |  fda & fde & FDM  |  FDA & FDE & FDM  ; 
assign ged = ~GED; //complement 
assign gfd =  FDA & fde & fdm  |  fda & FDE & fdm  |  fda & fde & FDM  |  fda & fde & fdm  ; 
assign GFD = ~gfd;  //complement 
assign GCI =  FCO & fcg & fck  |  fco & FCG & fck  |  fco & fcg & FCK  |  FCO & FCG & FCK  ; 
assign gci = ~GCI; //complement 
assign gdi =  FCO & fcg & fck  |  fco & FCG & fck  |  fco & fcg & FCK  |  fco & fcg & fck  ; 
assign GDI = ~gdi;  //complement 
assign GEA =  FED & fea & fel  |  fed & FEA & fel  |  fed & fea & FEL  |  FED & FEA & FEL  ; 
assign gea = ~GEA; //complement 
assign gfa =  FED & fea & fel  |  fed & FEA & fel  |  fed & fea & FEL  |  fed & fea & fel  ; 
assign GFA = ~gfa;  //complement 
assign GEE =  FEB & fef & fei  |  feb & FEF & fei  |  feb & fef & FEI  |  FEB & FEF & FEI  ; 
assign gee = ~GEE; //complement 
assign gfe =  FEB & fef & fei  |  feb & FEF & fei  |  feb & fef & FEI  |  feb & fef & fei  ; 
assign GFE = ~gfe;  //complement 
assign GEJ =  FDO & fdg & fdk  |  fdo & FDG & fdk  |  fdo & fdg & FDK  |  FDO & FDG & FDK  ; 
assign gej = ~GEJ; //complement 
assign gfj =  FDO & fdg & fdk  |  fdo & FDG & fdk  |  fdo & fdg & FDK  |  fdo & fdg & fdk  ; 
assign GFJ = ~gfj;  //complement 
assign GEF =  FDI & fdb & fdf  |  fdi & FDB & fdf  |  fdi & fdb & FDF  |  FDI & FDB & FDF  ; 
assign gef = ~GEF; //complement 
assign gff =  FDI & fdb & fdf  |  fdi & FDB & fdf  |  fdi & fdb & FDF  |  fdi & fdb & fdf  ; 
assign GFF = ~gff;  //complement 
assign GGD =  FFA & ffe & ffm  |  ffa & FFE & ffm  |  ffa & ffe & FFM  |  FFA & FFE & FFM  ; 
assign ggd = ~GGD; //complement 
assign ghd =  FFA & ffe & ffm  |  ffa & FFE & ffm  |  ffa & ffe & FFM  |  ffa & ffe & ffm  ; 
assign GHD = ~ghd;  //complement 
assign GEI =  FEO & feg & fek  |  feo & FEG & fek  |  feo & feg & FEK  |  FEO & FEG & FEK  ; 
assign gei = ~GEI; //complement 
assign gfi =  FEO & feg & fek  |  feo & FEG & fek  |  feo & feg & FEK  |  feo & feg & fek  ; 
assign GFI = ~gfi;  //complement 
assign GEG =  FEJ & fen & fec  |  fej & FEN & fec  |  fej & fen & FEC  |  FEJ & FEN & FEC  ; 
assign geg = ~GEG; //complement 
assign gfg =  FEJ & fen & fec  |  fej & FEN & fec  |  fej & fen & FEC  |  fej & fen & fec  ; 
assign GFG = ~gfg;  //complement 
assign GEC =  FEE & fem & feh  |  fee & FEM & feh  |  fee & fem & FEH  |  FEE & FEM & FEH  ; 
assign gec = ~GEC; //complement 
assign gfc =  FEE & fem & feh  |  fee & FEM & feh  |  fee & fem & FEH  |  fee & fem & feh  ; 
assign GFC = ~gfc;  //complement 
assign GGJ =  FFO & ffg & ffk  |  ffo & FFG & ffk  |  ffo & ffg & FFK  |  FFO & FFG & FFK  ; 
assign ggj = ~GGJ; //complement 
assign ghj =  FFO & ffg & ffk  |  ffo & FFG & ffk  |  ffo & ffg & FFK  |  ffo & ffg & ffk  ; 
assign GHJ = ~ghj;  //complement 
assign GGF =  FFI & ffb & fff  |  ffi & FFB & fff  |  ffi & ffb & FFF  |  FFI & FFB & FFF  ; 
assign ggf = ~GGF; //complement 
assign ghf =  FFI & ffb & fff  |  ffi & FFB & fff  |  ffi & ffb & FFF  |  ffi & ffb & fff  ; 
assign GHF = ~ghf;  //complement 
assign GGB =  FFD & ffl & ffh  |  ffd & FFL & ffh  |  ffd & ffl & FFH  |  FFD & FFL & FFH  ; 
assign ggb = ~GGB; //complement 
assign ghb =  FFD & ffl & ffh  |  ffd & FFL & ffh  |  ffd & ffl & FFH  |  ffd & ffl & ffh  ; 
assign GHB = ~ghb;  //complement 
assign GGH =  FFC & ffj & ffn  |  ffc & FFJ & ffn  |  ffc & ffj & FFN  |  FFC & FFJ & FFN  ; 
assign ggh = ~GGH; //complement 
assign ghh =  FFC & ffj & ffn  |  ffc & FFJ & ffn  |  ffc & ffj & FFN  |  ffc & ffj & ffn  ; 
assign GHH = ~ghh;  //complement 
assign GGG =  FGJ & fgn & fgc  |  fgj & FGN & fgc  |  fgj & fgn & FGC  |  FGJ & FGN & FGC  ; 
assign ggg = ~GGG; //complement 
assign ghg =  FGJ & fgn & fgc  |  fgj & FGN & fgc  |  fgj & fgn & FGC  |  fgj & fgn & fgc  ; 
assign GHG = ~ghg;  //complement 
assign GGC =  FGE & fgm & fgh  |  fge & FGM & fgh  |  fge & fgm & FGH  |  FGE & FGM & FGH  ; 
assign ggc = ~GGC; //complement 
assign ghc =  FGE & fgm & fgh  |  fge & FGM & fgh  |  fge & fgm & FGH  |  fge & fgm & fgh  ; 
assign GHC = ~ghc;  //complement 
assign GGA =  FGD & fga & fgl  |  fgd & FGA & fgl  |  fgd & fga & FGL  |  FGD & FGA & FGL  ; 
assign gga = ~GGA; //complement 
assign gha =  FGD & fga & fgl  |  fgd & FGA & fgl  |  fgd & fga & FGL  |  fgd & fga & fgl  ; 
assign GHA = ~gha;  //complement 
assign GGE =  FGB & fgf & fgi  |  fgb & FGF & fgi  |  fgb & fgf & FGI  |  FGB & FGF & FGI  ; 
assign gge = ~GGE; //complement 
assign ghe =  FGB & fgf & fgi  |  fgb & FGF & fgi  |  fgb & fgf & FGI  |  fgb & fgf & fgi  ; 
assign GHE = ~ghe;  //complement 
assign BBA = ~bba;  //complement 
assign BBB = ~bbb;  //complement 
assign BBC = ~bbc;  //complement 
assign BBD = ~bbd;  //complement 
assign BBE = ~bbe;  //complement 
assign BBF = ~bbf;  //complement 
assign BBG = ~bbg;  //complement 
assign BBH = ~bbh;  //complement 
assign BBI = ~bbi;  //complement 
assign BBJ = ~bbj;  //complement 
assign BBK = ~bbk;  //complement 
assign BBL = ~bbl;  //complement 
assign BBM = ~bbm;  //complement 
assign BBN = ~bbn;  //complement 
assign BBO = ~bbo;  //complement 
assign BBP = ~bbp;  //complement 
assign bca = ~BCA;  //complement 
assign bcb = ~BCB;  //complement 
assign bcc = ~BCC;  //complement 
assign bcd = ~BCD;  //complement 
assign bce = ~BCE;  //complement 
assign bcf = ~BCF;  //complement 
assign bcg = ~BCG;  //complement 
assign bch = ~BCH;  //complement 
assign bci = ~BCI;  //complement 
assign bcj = ~BCJ;  //complement 
assign bck = ~BCK;  //complement 
assign bcl = ~BCL;  //complement 
assign bcm = ~BCM;  //complement 
assign bcn = ~BCN;  //complement 
assign bco = ~BCO;  //complement 
assign bcp = ~BCP;  //complement 
assign GAB =  FAE & fam & fah  |  fae & FAM & fah  |  fae & fam & FAH  |  FAE & FAM & FAH  ; 
assign gab = ~GAB; //complement 
assign gbb =  FAE & fam & fah  |  fae & FAM & fah  |  fae & fam & FAH  |  fae & fam & fah  ; 
assign GBB = ~gbb;  //complement 
assign GAA =  FAD & faa & fal  |  fad & FAA & fal  |  fad & faa & FAL  |  FAD & FAA & FAL  ; 
assign gaa = ~GAA; //complement 
assign gba =  FAD & faa & fal  |  fad & FAA & fal  |  fad & faa & FAL  |  fad & faa & fal  ; 
assign GBA = ~gba;  //complement 
assign GAC =  FAB & fan & faf  |  fab & FAN & faf  |  fab & fan & FAF  |  FAB & FAN & FAF  ; 
assign gac = ~GAC; //complement 
assign gbc =  FAB & fan & faf  |  fab & FAN & faf  |  fab & fan & FAF  |  fab & fan & faf  ; 
assign GBC = ~gbc;  //complement 
assign HAE =  FAQ & gae & ilh  |  faq & GAE & ilh  |  faq & gae & ILH  |  FAQ & GAE & ILH  ; 
assign hae = ~HAE; //complement 
assign hbe =  FAQ & gae & ilh  |  faq & GAE & ilh  |  faq & gae & ILH  |  faq & gae & ilh  ; 
assign HBE = ~hbe;  //complement 
assign GAE =  FAP & fak & fao  |  fap & FAK & fao  |  fap & fak & FAO  |  FAP & FAK & FAO  ; 
assign gae = ~GAE; //complement 
assign gbe =  FAP & fak & fao  |  fap & FAK & fao  |  fap & fak & FAO  |  fap & fak & fao  ; 
assign GBE = ~gbe;  //complement 
assign GAD =  FAJ & fac & fag  |  faj & FAC & fag  |  faj & fac & FAG  |  FAJ & FAC & FAG  ; 
assign gad = ~GAD; //complement 
assign gbd =  FAJ & fac & fag  |  faj & FAC & fag  |  faj & fac & FAG  |  faj & fac & fag  ; 
assign GBD = ~gbd;  //complement 
assign GCB =  FBD & fbl & fbh  |  fbd & FBL & fbh  |  fbd & fbl & FBH  |  FBD & FBL & FBH  ; 
assign gcb = ~GCB; //complement 
assign gdb =  FBD & fbl & fbh  |  fbd & FBL & fbh  |  fbd & fbl & FBH  |  fbd & fbl & fbh  ; 
assign GDB = ~gdb;  //complement 
assign GCH =  FBC & fbj & fbn  |  fbc & FBJ & fbn  |  fbc & fbj & FBN  |  FBC & FBJ & FBN  ; 
assign gch = ~GCH; //complement 
assign gdh =  FBC & fbj & fbn  |  fbc & FBJ & fbn  |  fbc & fbj & FBN  |  fbc & fbj & fbn  ; 
assign GDH = ~gdh;  //complement 
assign GCD =  FBA & fbe & fbm  |  fba & FBE & fbm  |  fba & fbe & FBM  |  FBA & FBE & FBM  ; 
assign gcd = ~GCD; //complement 
assign gdd =  FBA & fbe & fbm  |  fba & FBE & fbm  |  fba & fbe & FBM  |  fba & fbe & fbm  ; 
assign GDD = ~gdd;  //complement 
assign GCE =  FCB & fcf & fci  |  fcb & FCF & fci  |  fcb & fcf & FCI  |  FCB & FCF & FCI  ; 
assign gce = ~GCE; //complement 
assign gde =  FCB & fcf & fci  |  fcb & FCF & fci  |  fcb & fcf & FCI  |  fcb & fcf & fci  ; 
assign GDE = ~gde;  //complement 
assign GCJ =  FBO & fbg & fbk  |  fbo & FBG & fbk  |  fbo & fbg & FBK  |  FBO & FBG & FBK  ; 
assign gcj = ~GCJ; //complement 
assign gdj =  FBO & fbg & fbk  |  fbo & FBG & fbk  |  fbo & fbg & FBK  |  fbo & fbg & fbk  ; 
assign GDJ = ~gdj;  //complement 
assign GCF =  FBI & fbb & fbf  |  fbi & FBB & fbf  |  fbi & fbb & FBF  |  FBI & FBB & FBF  ; 
assign gcf = ~GCF; //complement 
assign gdf =  FBI & fbb & fbf  |  fbi & FBB & fbf  |  fbi & fbb & FBF  |  fbi & fbb & fbf  ; 
assign GDF = ~gdf;  //complement 
assign GCG =  FCJ & fcn & fcc  |  fcj & FCN & fcc  |  fcj & fcn & FCC  |  FCJ & FCN & FCC  ; 
assign gcg = ~GCG; //complement 
assign gdg =  FCJ & fcn & fcc  |  fcj & FCN & fcc  |  fcj & fcn & FCC  |  fcj & fcn & fcc  ; 
assign GDG = ~gdg;  //complement 
assign qta = ~QTA;  //complement 
assign tta = ~TTA;  //complement 
assign ttb = ~TTB;  //complement 
assign ttc = ~TTC;  //complement 
assign GCC =  FCE & fcm & fch  |  fce & FCM & fch  |  fce & fcm & FCH  |  FCE & FCM & FCH  ; 
assign gcc = ~GCC; //complement 
assign gdc =  FCE & fcm & fch  |  fce & FCM & fch  |  fce & fcm & FCH  |  fce & fcm & fch  ; 
assign GDC = ~gdc;  //complement 
assign GCA =  FCD & fca & fcl  |  fcd & FCA & fcl  |  fcd & fca & FCL  |  FCD & FCA & FCL  ; 
assign gca = ~GCA; //complement 
assign gda =  FCD & fca & fcl  |  fcd & FCA & fcl  |  fcd & fca & FCL  |  fcd & fca & fcl  ; 
assign GDA = ~gda;  //complement 
assign EAK = DAK & CCH ; 
assign eak = ~EAK ; //complement 
assign ECK = DAK & CCI ; 
assign eck = ~ECK ;  //complement 
assign EEK = DAK & CCJ ; 
assign eek = ~EEK ;  //complement 
assign EIK = DAK & CCL; 
assign eik = ~EIK; 
assign ECL = DAL & CCH ; 
assign ecl = ~ECL ; //complement 
assign EEL = DAL & CCI ; 
assign eel = ~EEL ;  //complement 
assign EIL = DAL & CCK ; 
assign eil = ~EIL ;  //complement 
assign EKL = DAL & CCL; 
assign ekl = ~EKL; 
assign opi = ~OPI;  //complement 
assign OQI = ~oqi;  //complement 
assign cbe = ~CBE;  //complement 
assign cee = ~CEE;  //complement 
assign cbf = ~CBF;  //complement 
assign cef = ~CEF;  //complement 
assign EAM = DAM & CCF ; 
assign eam = ~EAM ; //complement 
assign ECM = DAM & CCG ; 
assign ecm = ~ECM ;  //complement 
assign EEM = DAM & CCH ; 
assign eem = ~EEM ;  //complement 
assign EIM = DAM & CCJ; 
assign eim = ~EIM; 
assign EAN = DAN & CCE ; 
assign ean = ~EAN ; //complement 
assign ECN = DAN & CCF ; 
assign ecn = ~ECN ;  //complement 
assign EEN = DAN & CCG ; 
assign een = ~EEN ;  //complement 
assign EIN = DAN & CCI; 
assign ein = ~EIN; 
assign bdm = ~BDM;  //complement 
assign bdn = ~BDN;  //complement 
assign bdo = ~BDO;  //complement 
assign bdp = ~BDP;  //complement 
assign cbg = ~CBG;  //complement 
assign cbh = ~CBH;  //complement 
assign cbi = ~CBI;  //complement 
assign EEO = DAO & CCF ; 
assign eeo = ~EEO ; //complement 
assign EAO = DAO & CCD ; 
assign eao = ~EAO ;  //complement 
assign ECO = DAO & CCE ; 
assign eco = ~ECO ;  //complement 
assign EIO = DAO & CCH; 
assign eio = ~EIO; 
assign EAP = DAP & CCC ; 
assign eap = ~EAP ; //complement 
assign ECP = DAP & CCD ; 
assign ecp = ~ECP ;  //complement 
assign EEP = DAP & CCE ; 
assign eep = ~EEP ;  //complement 
assign EIP = DAP & CCG; 
assign eip = ~EIP; 
assign opo = ~OPO;  //complement 
assign OQO = ~oqo;  //complement 
assign ceg = ~CEG;  //complement 
assign ceh = ~CEH;  //complement 
assign cei = ~CEI;  //complement 
assign EAQ = DBA & CCB ; 
assign eaq = ~EAQ ; //complement 
assign ECQ = DBA & CCC ; 
assign ecq = ~ECQ ;  //complement 
assign EEQ = DBA & CCD ; 
assign eeq = ~EEQ ;  //complement 
assign EIQ = DBA & CCF; 
assign eiq = ~EIQ; 
assign EAR = DBB & CCA ; 
assign ear = ~EAR ; //complement 
assign ECR = DBB & CCB ; 
assign ecr = ~ECR ;  //complement 
assign EER = DBB & CCC ; 
assign eer = ~EER ;  //complement 
assign opq = ~OPQ;  //complement 
assign OQQ = ~oqq;  //complement 
assign opr = ~OPR;  //complement 
assign EKN = DAN & CCJ ; 
assign ekn = ~EKN ; //complement 
assign EAS = DBC & CBP ; 
assign eas = ~EAS ; //complement 
assign ECS = DBC & CCA ; 
assign ecs = ~ECS ;  //complement 
assign EES = DBC & CCB ; 
assign ees = ~EES ;  //complement 
assign EIS = DBC & CCD; 
assign eis = ~EIS; 
assign EAT = DBD & CBO ; 
assign eat = ~EAT ; //complement 
assign ECT = DBD & CBP ; 
assign ect = ~ECT ;  //complement 
assign EET = DBD & CCA ; 
assign eet = ~EET ;  //complement 
assign EIT = DBD & CCC; 
assign eit = ~EIT; 
assign qka = ~QKA;  //complement 
assign tka = ~TKA;  //complement 
assign tkb = ~TKB;  //complement 
assign tkc = ~TKC;  //complement 
assign dca = ~DCA;  //complement 
assign DFA = ~dfa;  //complement 
assign dcb = ~DCB;  //complement 
assign DFB = ~dfb;  //complement 
assign EAU = DBE & CBN ; 
assign eau = ~EAU ; //complement 
assign ECU = DBE & CBO ; 
assign ecu = ~ECU ;  //complement 
assign EEU = DBE & CBP ; 
assign eeu = ~EEU ;  //complement 
assign EAV = DBF & CBM ; 
assign eav = ~EAV ; //complement 
assign ECV = DBF & CBN ; 
assign ecv = ~ECV ;  //complement 
assign EEV = DBF & CBO ; 
assign eev = ~EEV ;  //complement 
assign EIV = DBF & CCA; 
assign eiv = ~EIV; 
assign tkd = ~TKD;  //complement 
assign tke = ~TKE;  //complement 
assign tkf = ~TKF;  //complement 
assign dcc = ~DCC;  //complement 
assign DFC = ~dfc;  //complement 
assign dcd = ~DCD;  //complement 
assign DFD = ~dfd;  //complement 
assign EAW = DBG & CBL ; 
assign eaw = ~EAW ; //complement 
assign ECW = DBG & CBM ; 
assign ecw = ~ECW ;  //complement 
assign EEW = DBG & CBN ; 
assign eew = ~EEW ;  //complement 
assign EIW = DBG & CBP; 
assign eiw = ~EIW; 
assign EAX = DBH & CBK ; 
assign eax = ~EAX ; //complement 
assign ECX = DBH & CBL ; 
assign ecx = ~ECX ;  //complement 
assign EEX = DBH & CBM ; 
assign eex = ~EEX ;  //complement 
assign EIX = DBH & CBO; 
assign eix = ~EIX; 
assign opk = ~OPK;  //complement 
assign OQK = ~oqk;  //complement 
assign dce = ~DCE;  //complement 
assign DFE = ~dfe;  //complement 
assign dcf = ~DCF;  //complement 
assign DFF = ~dff;  //complement 
assign bda = ~BDA;  //complement 
assign bdb = ~BDB;  //complement 
assign bdc = ~BDC;  //complement 
assign bdd = ~BDD;  //complement 
assign bde = ~BDE;  //complement 
assign bdf = ~BDF;  //complement 
assign bdg = ~BDG;  //complement 
assign bdh = ~BDH;  //complement 
assign bdi = ~BDI;  //complement 
assign bdj = ~BDJ;  //complement 
assign bdk = ~BDK;  //complement 
assign bdl = ~BDL;  //complement 
assign dcg = ~DCG;  //complement 
assign DFG = ~dfg;  //complement 
assign dch = ~DCH;  //complement 
assign DFH = ~dfh;  //complement 
assign GMI =  FMI & fmj & fmf  |  fmi & FMJ & fmf  |  fmi & fmj & FMF  |  FMI & FMJ & FMF  ; 
assign gmi = ~GMI; //complement 
assign gni =  FMI & fmj & fmf  |  fmi & FMJ & fmf  |  fmi & fmj & FMF  |  fmi & fmj & fmf  ; 
assign GNI = ~gni;  //complement 
assign GMD =  FMA & fmg & fmd  |  fma & FMG & fmd  |  fma & fmg & FMD  |  FMA & FMG & FMD  ; 
assign gmd = ~GMD; //complement 
assign gnd =  FMA & fmg & fmd  |  fma & FMG & fmd  |  fma & fmg & FMD  |  fma & fmg & fmd  ; 
assign GND = ~gnd;  //complement 
assign GMF =  FLN & flf & fmb  |  fln & FLF & fmb  |  fln & flf & FMB  |  FLN & FLF & FMB  ; 
assign gmf = ~GMF; //complement 
assign gnf =  FLN & flf & fmb  |  fln & FLF & fmb  |  fln & flf & FMB  |  fln & flf & fmb  ; 
assign GNF = ~gnf;  //complement 
assign GMG =  FLJ & flc & fme  |  flj & FLC & fme  |  flj & flc & FME  |  FLJ & FLC & FME  ; 
assign gmg = ~GMG; //complement 
assign gng =  FLJ & flc & fme  |  flj & FLC & fme  |  flj & flc & FME  |  flj & flc & fme  ; 
assign GNG = ~gng;  //complement 
assign GOC =  FND & fnl & fol  |  fnd & FNL & fol  |  fnd & fnl & FOL  |  FND & FNL & FOL  ; 
assign goc = ~GOC; //complement 
assign gpc =  FND & fnl & fol  |  fnd & FNL & fol  |  fnd & fnl & FOL  |  fnd & fnl & fol  ; 
assign GPC = ~gpc;  //complement 
assign GOA =  FNC & fnk & foc  |  fnc & FNK & foc  |  fnc & fnk & FOC  |  FNC & FNK & FOC  ; 
assign goa = ~GOA; //complement 
assign gpa =  FNC & fnk & foc  |  fnc & FNK & foc  |  fnc & fnk & FOC  |  fnc & fnk & foc  ; 
assign GPA = ~gpa;  //complement 
assign GOE =  FNB & fnh & foh  |  fnb & FNH & foh  |  fnb & fnh & FOH  |  FNB & FNH & FOH  ; 
assign goe = ~GOE; //complement 
assign gpe =  FNB & fnh & foh  |  fnb & FNH & foh  |  fnb & fnh & FOH  |  fnb & fnh & foh  ; 
assign GPE = ~gpe;  //complement 
assign GOB =  FNA & fng & fok  |  fna & FNG & fok  |  fna & fng & FOK  |  FNA & FNG & FOK  ; 
assign gob = ~GOB; //complement 
assign gpb =  FNA & fng & fok  |  fna & FNG & fok  |  fna & fng & FOK  |  fna & fng & fok  ; 
assign GPB = ~gpb;  //complement 
assign GOD =  FOG & foa & fod  |  fog & FOA & fod  |  fog & foa & FOD  |  FOG & FOA & FOD  ; 
assign god = ~GOD; //complement 
assign gpd =  FOG & foa & fod  |  fog & FOA & fod  |  fog & foa & FOD  |  fog & foa & fod  ; 
assign GPD = ~gpd;  //complement 
assign GOG =  FNI & foe & fom  |  fni & FOE & fom  |  fni & foe & FOM  |  FNI & FOE & FOM  ; 
assign gog = ~GOG; //complement 
assign gpg =  FNI & foe & fom  |  fni & FOE & fom  |  fni & foe & FOM  |  fni & foe & fom  ; 
assign GPG = ~gpg;  //complement 
assign GOH =  FNF & fnj & fon  |  fnf & FNJ & fon  |  fnf & fnj & FON  |  FNF & FNJ & FON  ; 
assign goh = ~GOH; //complement 
assign gph =  FNF & fnj & fon  |  fnf & FNJ & fon  |  fnf & fnj & FON  |  fnf & fnj & fon  ; 
assign GPH = ~gph;  //complement 
assign GOF =  FNE & fnm & fob  |  fne & FNM & fob  |  fne & fnm & FOB  |  FNE & FNM & FOB  ; 
assign gof = ~GOF; //complement 
assign gpf =  FNE & fnm & fob  |  fne & FNM & fob  |  fne & fnm & FOB  |  fne & fnm & fob  ; 
assign GPF = ~gpf;  //complement 
assign GQA =  FPC & fqc & fpk  |  fpc & FQC & fpk  |  fpc & fqc & FPK  |  FPC & FQC & FPK  ; 
assign gqa = ~GQA; //complement 
assign gra =  FPC & fqc & fpk  |  fpc & FQC & fpk  |  fpc & fqc & FPK  |  fpc & fqc & fpk  ; 
assign GRA = ~gra;  //complement 
assign GQC =  FPD & fpl & fql  |  fpd & FPL & fql  |  fpd & fpl & FQL  |  FPD & FPL & FQL  ; 
assign gqc = ~GQC; //complement 
assign grc =  FPD & fpl & fql  |  fpd & FPL & fql  |  fpd & fpl & FQL  |  fpd & fpl & fql  ; 
assign GRC = ~grc;  //complement 
assign GQB =  FPA & fpg & fqk  |  fpa & FPG & fqk  |  fpa & fpg & FQK  |  FPA & FPG & FQK  ; 
assign gqb = ~GQB; //complement 
assign grb =  FPA & fpg & fqk  |  fpa & FPG & fqk  |  fpa & fpg & FQK  |  fpa & fpg & fqk  ; 
assign GRB = ~grb;  //complement 
assign GOI =  FOJ & foi & fof  |  foj & FOI & fof  |  foj & foi & FOF  |  FOJ & FOI & FOF  ; 
assign goi = ~GOI; //complement 
assign gpi =  FOJ & foi & fof  |  foj & FOI & fof  |  foj & foi & FOF  |  foj & foi & fof  ; 
assign GPI = ~gpi;  //complement 
assign bem = ~BEM;  //complement 
assign ben = ~BEN;  //complement 
assign beo = ~BEO;  //complement 
assign bep = ~BEP;  //complement 
assign GQH =  FPJ & fpf & fqf  |  fpj & FPF & fqf  |  fpj & fpf & FQF  |  FPJ & FPF & FQF  ; 
assign gqh = ~GQH; //complement 
assign grh =  FPJ & fpf & fqf  |  fpj & FPF & fqf  |  fpj & fpf & FQF  |  fpj & fpf & fqf  ; 
assign GRH = ~grh;  //complement 
assign GQG =  FPI & fqi & fqm  |  fpi & FQI & fqm  |  fpi & fqi & FQM  |  FPI & FQI & FQM  ; 
assign gqg = ~GQG; //complement 
assign grg =  FPI & fqi & fqm  |  fpi & FQI & fqm  |  fpi & fqi & FQM  |  fpi & fqi & fqm  ; 
assign GRG = ~grg;  //complement 
assign GQE =  FPH & fpb & fqh  |  fph & FPB & fqh  |  fph & fpb & FQH  |  FPH & FPB & FQH  ; 
assign gqe = ~GQE; //complement 
assign gre =  FPH & fpb & fqh  |  fph & FPB & fqh  |  fph & fpb & FQH  |  fph & fpb & fqh  ; 
assign GRE = ~gre;  //complement 
assign GQF =  FPE & fqb & fpm  |  fpe & FQB & fpm  |  fpe & fqb & FPM  |  FPE & FQB & FPM  ; 
assign gqf = ~GQF; //complement 
assign grf =  FPE & fqb & fpm  |  fpe & FQB & fpm  |  fpe & fqb & FPM  |  fpe & fqb & fpm  ; 
assign GRF = ~grf;  //complement 
assign bea = ~BEA;  //complement 
assign beb = ~BEB;  //complement 
assign bec = ~BEC;  //complement 
assign bed = ~BED;  //complement 
assign bee = ~BEE;  //complement 
assign bef = ~BEF;  //complement 
assign beg = ~BEG;  //complement 
assign beh = ~BEH;  //complement 
assign bei = ~BEI;  //complement 
assign bej = ~BEJ;  //complement 
assign bek = ~BEK;  //complement 
assign bel = ~BEL;  //complement 
assign GQD =  FQA & fqg & fqd  |  fqa & FQG & fqd  |  fqa & fqg & FQD  |  FQA & FQG & FQD  ; 
assign gqd = ~GQD; //complement 
assign grd =  FQA & fqg & fqd  |  fqa & FQG & fqd  |  fqa & fqg & FQD  |  fqa & fqg & fqd  ; 
assign GRD = ~grd;  //complement 
assign cbj = ~CBJ;  //complement 
assign cbk = ~CBK;  //complement 
assign cbl = ~CBL;  //complement 
assign cej = ~CEJ;  //complement 
assign cek = ~CEK;  //complement 
assign cel = ~CEL;  //complement 
assign GIH =  FHC & fhj & fhn  |  fhc & FHJ & fhn  |  fhc & fhj & FHN  |  FHC & FHJ & FHN  ; 
assign gih = ~GIH; //complement 
assign gjh =  FHC & fhj & fhn  |  fhc & FHJ & fhn  |  fhc & fhj & FHN  |  fhc & fhj & fhn  ; 
assign GJH = ~gjh;  //complement 
assign GID =  FHA & fhe & fhm  |  fha & FHE & fhm  |  fha & fhe & FHM  |  FHA & FHE & FHM  ; 
assign gid = ~GID; //complement 
assign gjd =  FHA & fhe & fhm  |  fha & FHE & fhm  |  fha & fhe & FHM  |  fha & fhe & fhm  ; 
assign GJD = ~gjd;  //complement 
assign GGI =  FGP & fgg & fgk  |  fgp & FGG & fgk  |  fgp & fgg & FGK  |  FGP & FGG & FGK  ; 
assign ggi = ~GGI; //complement 
assign ghi =  FGP & fgg & fgk  |  fgp & FGG & fgk  |  fgp & fgg & FGK  |  fgp & fgg & fgk  ; 
assign GHI = ~ghi;  //complement 
assign GIE =  FIB & fif & fii  |  fib & FIF & fii  |  fib & fif & FII  |  FIB & FIF & FII  ; 
assign gie = ~GIE; //complement 
assign gje =  FIB & fif & fii  |  fib & FIF & fii  |  fib & fif & FII  |  fib & fif & fii  ; 
assign GJE = ~gje;  //complement 
assign GIF =  FHI & fhb & fhf  |  fhi & FHB & fhf  |  fhi & fhb & FHF  |  FHI & FHB & FHF  ; 
assign gif = ~GIF; //complement 
assign gjf =  FHI & fhb & fhf  |  fhi & FHB & fhf  |  fhi & fhb & FHF  |  fhi & fhb & fhf  ; 
assign GJF = ~gjf;  //complement 
assign GIB =  FHD & fhl & fhh  |  fhd & FHL & fhh  |  fhd & fhl & FHH  |  FHD & FHL & FHH  ; 
assign gib = ~GIB; //complement 
assign gjb =  FHD & fhl & fhh  |  fhd & FHL & fhh  |  fhd & fhl & FHH  |  fhd & fhl & fhh  ; 
assign GJB = ~gjb;  //complement 
assign GIG =  FIJ & fin & fic  |  fij & FIN & fic  |  fij & fin & FIC  |  FIJ & FIN & FIC  ; 
assign gig = ~GIG; //complement 
assign gjg =  FIJ & fin & fic  |  fij & FIN & fic  |  fij & fin & FIC  |  fij & fin & fic  ; 
assign GJG = ~gjg;  //complement 
assign GIC =  FIE & fim & fih  |  fie & FIM & fih  |  fie & fim & FIH  |  FIE & FIM & FIH  ; 
assign gic = ~GIC; //complement 
assign gjc =  FIE & fim & fih  |  fie & FIM & fih  |  fie & fim & FIH  |  fie & fim & fih  ; 
assign GJC = ~gjc;  //complement 
assign GIA =  FID & fia & fil  |  fid & FIA & fil  |  fid & fia & FIL  |  FID & FIA & FIL  ; 
assign gia = ~GIA; //complement 
assign gja =  FID & fia & fil  |  fid & FIA & fil  |  fid & fia & FIL  |  fid & fia & fil  ; 
assign GJA = ~gja;  //complement 
assign GKH =  FJC & fjj & fjn  |  fjc & FJJ & fjn  |  fjc & fjj & FJN  |  FJC & FJJ & FJN  ; 
assign gkh = ~GKH; //complement 
assign glh =  FJC & fjj & fjn  |  fjc & FJJ & fjn  |  fjc & fjj & FJN  |  fjc & fjj & fjn  ; 
assign GLH = ~glh;  //complement 
assign GKD =  FJA & fje & fjm  |  fja & FJE & fjm  |  fja & fje & FJM  |  FJA & FJE & FJM  ; 
assign gkd = ~GKD; //complement 
assign gld =  FJA & fje & fjm  |  fja & FJE & fjm  |  fja & fje & FJM  |  fja & fje & fjm  ; 
assign GLD = ~gld;  //complement 
assign GII =  FIO & fig & fik  |  fio & FIG & fik  |  fio & fig & FIK  |  FIO & FIG & FIK  ; 
assign gii = ~GII; //complement 
assign gji =  FIO & fig & fik  |  fio & FIG & fik  |  fio & fig & FIK  |  fio & fig & fik  ; 
assign GJI = ~gji;  //complement 
assign GKE =  FKB & fkf & fki  |  fkb & FKF & fki  |  fkb & fkf & FKI  |  FKB & FKF & FKI  ; 
assign gke = ~GKE; //complement 
assign gle =  FKB & fkf & fki  |  fkb & FKF & fki  |  fkb & fkf & FKI  |  fkb & fkf & fki  ; 
assign GLE = ~gle;  //complement 
assign GKF =  FJI & fjb & fjf  |  fji & FJB & fjf  |  fji & fjb & FJF  |  FJI & FJB & FJF  ; 
assign gkf = ~GKF; //complement 
assign glf =  FJI & fjb & fjf  |  fji & FJB & fjf  |  fji & fjb & FJF  |  fji & fjb & fjf  ; 
assign GLF = ~glf;  //complement 
assign GKB =  FJD & fjl & fjh  |  fjd & FJL & fjh  |  fjd & fjl & FJH  |  FJD & FJL & FJH  ; 
assign gkb = ~GKB; //complement 
assign glb =  FJD & fjl & fjh  |  fjd & FJL & fjh  |  fjd & fjl & FJH  |  fjd & fjl & fjh  ; 
assign GLB = ~glb;  //complement 
assign GKG =  FKJ & fkn & fkc  |  fkj & FKN & fkc  |  fkj & fkn & FKC  |  FKJ & FKN & FKC  ; 
assign gkg = ~GKG; //complement 
assign glg =  FKJ & fkn & fkc  |  fkj & FKN & fkc  |  fkj & fkn & FKC  |  fkj & fkn & fkc  ; 
assign GLG = ~glg;  //complement 
assign NQA =  MQA & mqb & mqc  |  mqa & MQB & mqc  |  mqa & mqb & MQC  |  MQA & MQB & MQC  ; 
assign nqa = ~NQA; //complement 
assign nra =  MQA & mqb & mqc  |  mqa & MQB & mqc  |  mqa & mqb & MQC  |  mqa & mqb & mqc  ; 
assign NRA = ~nra;  //complement 
assign GKC =  FKE & fkm & fkh  |  fke & FKM & fkh  |  fke & fkm & FKH  |  FKE & FKM & FKH  ; 
assign gkc = ~GKC; //complement 
assign glc =  FKE & fkm & fkh  |  fke & FKM & fkh  |  fke & fkm & FKH  |  fke & fkm & fkh  ; 
assign GLC = ~glc;  //complement 
assign GKA =  FKD & fka & fkl  |  fkd & FKA & fkl  |  fkd & fka & FKL  |  FKD & FKA & FKL  ; 
assign gka = ~GKA; //complement 
assign gla =  FKD & fka & fkl  |  fkd & FKA & fkl  |  fkd & fka & FKL  |  fkd & fka & fkl  ; 
assign GLA = ~gla;  //complement 
assign GME =  FLB & fli & fmh  |  flb & FLI & fmh  |  flb & fli & FMH  |  FLB & FLI & FMH  ; 
assign gme = ~GME; //complement 
assign gne =  FLB & fli & fmh  |  flb & FLI & fmh  |  flb & fli & FMH  |  flb & fli & fmh  ; 
assign GNE = ~gne;  //complement 
assign GMB =  FLA & flh & fmk  |  fla & FLH & fmk  |  fla & flh & FMK  |  FLA & FLH & FMK  ; 
assign gmb = ~GMB; //complement 
assign gnb =  FLA & flh & fmk  |  fla & FLH & fmk  |  fla & flh & FMK  |  fla & flh & fmk  ; 
assign GNB = ~gnb;  //complement 
assign GKI =  FKK & fkg & fjk  |  fkk & FKG & fjk  |  fkk & fkg & FJK  |  FKK & FKG & FJK  ; 
assign gki = ~GKI; //complement 
assign gli =  FKK & fkg & fjk  |  fkk & FKG & fjk  |  fkk & fkg & FJK  |  fkk & fkg & fjk  ; 
assign GLI = ~gli;  //complement 
assign GMH =  FLG & flk & fmn  |  flg & FLK & fmn  |  flg & flk & FMN  |  FLG & FLK & FMN  ; 
assign gmh = ~GMH; //complement 
assign gnh =  FLG & flk & fmn  |  flg & FLK & fmn  |  flg & flk & FMN  |  flg & flk & fmn  ; 
assign GNH = ~gnh;  //complement 
assign GMC =  FLE & flm & fml  |  fle & FLM & fml  |  fle & flm & FML  |  FLE & FLM & FML  ; 
assign gmc = ~GMC; //complement 
assign gnc =  FLE & flm & fml  |  fle & FLM & fml  |  fle & flm & FML  |  fle & flm & fml  ; 
assign GNC = ~gnc;  //complement 
assign GMA =  FLD & fmc & fll  |  fld & FMC & fll  |  fld & fmc & FLL  |  FLD & FMC & FLL  ; 
assign gma = ~GMA; //complement 
assign gna =  FLD & fmc & fll  |  fld & FMC & fll  |  fld & fmc & FLL  |  fld & fmc & fll  ; 
assign GNA = ~gna;  //complement 
assign ope = ~OPE;  //complement 
assign OQE = ~oqe;  //complement 
assign opf = ~OPF;  //complement 
assign EBB = DBJ & CBI ; 
assign ebb = ~EBB ; //complement 
assign EDB = DBJ & CBJ ; 
assign edb = ~EDB ;  //complement 
assign EFB = DBJ & CBK ; 
assign efb = ~EFB ;  //complement 
assign EJB = DBJ & CBM; 
assign ejb = ~EJB; 
assign opg = ~OPG;  //complement 
assign oph = ~OPH;  //complement 
assign cbm = ~CBM;  //complement 
assign cbn = ~CBN;  //complement 
assign cbo = ~CBO;  //complement 
assign EBC = DBK & CBH ; 
assign ebc = ~EBC ; //complement 
assign EDC = DBK & CBI ; 
assign edc = ~EDC ;  //complement 
assign EFC = DBK & CBJ ; 
assign efc = ~EFC ;  //complement 
assign EJC = DBK & CBL; 
assign ejc = ~EJC; 
assign EBD = DBL & CBG ; 
assign ebd = ~EBD ; //complement 
assign EDD = DBL & CBH ; 
assign edd = ~EDD ;  //complement 
assign EFD = DBL & CBI ; 
assign efd = ~EFD ;  //complement 
assign EJD = DBL & CBK; 
assign ejd = ~EJD; 
assign opm = ~OPM;  //complement 
assign OQM = ~oqm;  //complement 
assign cem = ~CEM;  //complement 
assign cen = ~CEN;  //complement 
assign ceo = ~CEO;  //complement 
assign opa = ~OPA;  //complement 
assign OQA = ~oqa;  //complement 
assign opb = ~OPB;  //complement 
assign EBF = DBN & CBE ; 
assign ebf = ~EBF ; //complement 
assign EDF = DBN & CBF ; 
assign edf = ~EDF ;  //complement 
assign EFF = DBN & CBG ; 
assign eff = ~EFF ;  //complement 
assign EJF = DBN & CBI; 
assign ejf = ~EJF; 
assign cbp = ~CBP;  //complement 
assign cep = ~CEP;  //complement 
assign EBG = DBO & CBD ; 
assign ebg = ~EBG ; //complement 
assign EDG = DBO & CBE ; 
assign edg = ~EDG ;  //complement 
assign EFG = DBO & CBF ; 
assign efg = ~EFG ;  //complement 
assign EJG = DBO & CBH; 
assign ejg = ~EJG; 
assign EBH = DBP & CBC ; 
assign ebh = ~EBH ; //complement 
assign EDH = DBP & CBD ; 
assign edh = ~EDH ;  //complement 
assign EFH = DBP & CBE ; 
assign efh = ~EFH ;  //complement 
assign EJH = DBP & CBG; 
assign ejh = ~EJH; 
assign opc = ~OPC;  //complement 
assign OQC = ~oqc;  //complement 
assign opd = ~OPD;  //complement 
assign qga = ~QGA;  //complement 
assign tga = ~TGA;  //complement 
assign tgb = ~TGB;  //complement 
assign tgc = ~TGC;  //complement 
assign EBI = DCA & CBB ; 
assign ebi = ~EBI ; //complement 
assign EDI = DCA & CBC ; 
assign edi = ~EDI ;  //complement 
assign EFI = DCA & CBD ; 
assign efi = ~EFI ;  //complement 
assign EJI = DCA & CBF; 
assign eji = ~EJI; 
assign EBK = DCC & CAP ; 
assign ebk = ~EBK ; //complement 
assign EDK = DCC & CBA ; 
assign edk = ~EDK ;  //complement 
assign EFK = DCC & CBB ; 
assign efk = ~EFK ;  //complement 
assign EJK = DCC & CBD; 
assign ejk = ~EJK; 
assign dci = ~DCI;  //complement 
assign DFI = ~dfi;  //complement 
assign dcj = ~DCJ;  //complement 
assign DFJ = ~dfj;  //complement 
assign EBL = DCD & CAO ; 
assign ebl = ~EBL ; //complement 
assign EDL = DCD & CAP ; 
assign edl = ~EDL ;  //complement 
assign EFL = DCD & CBA ; 
assign efl = ~EFL ;  //complement 
assign EJL = DCD & CBC; 
assign ejl = ~EJL; 
assign EBM = DCE & CAN ; 
assign ebm = ~EBM ; //complement 
assign EDM = DCE & CAO ; 
assign edm = ~EDM ;  //complement 
assign EFM = DCE & CAP ; 
assign efm = ~EFM ;  //complement 
assign EJM = DCE & CBB; 
assign ejm = ~EJM; 
assign dck = ~DCK;  //complement 
assign DFK = ~dfk;  //complement 
assign dcl = ~DCL;  //complement 
assign DFL = ~dfl;  //complement 
assign EBN = DCF & CAM ; 
assign ebn = ~EBN ; //complement 
assign EDN = DCF & CAN ; 
assign edn = ~EDN ;  //complement 
assign EFN = DCF & CAO ; 
assign efn = ~EFN ;  //complement 
assign EJN = DCF & CBA; 
assign ejn = ~EJN; 
assign EBO = DCG & CAL ; 
assign ebo = ~EBO ; //complement 
assign EDO = DCG & CAM ; 
assign edo = ~EDO ;  //complement 
assign EFO = DCG & CAN ; 
assign efo = ~EFO ;  //complement 
assign EJO = DCG & CAP; 
assign ejo = ~EJO; 
assign EBE = DBM & CBF ; 
assign ebe = ~EBE ; //complement 
assign EDE = DBM & CBG ; 
assign ede = ~EDE ;  //complement 
assign EFE = DBM & CBH ; 
assign efe = ~EFE ;  //complement 
assign EJE = DBM & CBJ; 
assign eje = ~EJE; 
assign dcm = ~DCM;  //complement 
assign DFM = ~dfm;  //complement 
assign dcn = ~DCN;  //complement 
assign DFN = ~dfn;  //complement 
assign EBP = DCH & CAK ; 
assign ebp = ~EBP ; //complement 
assign EDP = DCH & CAL ; 
assign edp = ~EDP ;  //complement 
assign EFP = DCH & CAM ; 
assign efp = ~EFP ;  //complement 
assign EJP = DCH & CAO; 
assign ejp = ~EJP; 
assign EBQ = DCI & CAJ ; 
assign ebq = ~EBQ ; //complement 
assign EDQ = DCI & CAK ; 
assign edq = ~EDQ ;  //complement 
assign EFQ = DCI & CAL ; 
assign efq = ~EFQ ;  //complement 
assign EJQ = DCI & CAN; 
assign ejq = ~EJQ; 
assign EBA = DBI & CBJ ; 
assign eba = ~EBA ; //complement 
assign EDA = DBI & CBK ; 
assign eda = ~EDA ;  //complement 
assign EFA = DBI & CBL ; 
assign efa = ~EFA ;  //complement 
assign EJA = DBI & CBN; 
assign eja = ~EJA; 
assign dco = ~DCO;  //complement 
assign DFO = ~dfo;  //complement 
assign dcp = ~DCP;  //complement 
assign DFP = ~dfp;  //complement 
assign hib = ~HIB;  //complement 
assign HJB = ~hjb;  //complement 
assign hgg = ~HGG;  //complement 
assign HHG = ~hhg;  //complement 
assign hgd = ~HGD;  //complement 
assign HHD = ~hhd;  //complement 
assign hqf = ~HQF;  //complement 
assign OHF = ~ohf;  //complement 
assign hqg = ~HQG;  //complement 
assign hie = ~HIE;  //complement 
assign HJE = ~hje;  //complement 
assign hif = ~HIF;  //complement 
assign HJF = ~hjf;  //complement 
assign hic = ~HIC;  //complement 
assign HJC = ~hjc;  //complement 
assign hia = ~HIA;  //complement 
assign HJA = ~hja;  //complement 
assign hka = ~HKA;  //complement 
assign HLA = ~hla;  //complement 
assign hkb = ~HKB;  //complement 
assign HLB = ~hlb;  //complement 
assign hig = ~HIG;  //complement 
assign HJG = ~hjg;  //complement 
assign hid = ~HID;  //complement 
assign HJD = ~hjd;  //complement 
assign hke = ~HKE;  //complement 
assign HLE = ~hle;  //complement 
assign hkc = ~HKC;  //complement 
assign HLC = ~hlc;  //complement 
assign hkf = ~HKF;  //complement 
assign HLF = ~hlf;  //complement 
assign hkg = ~HKG;  //complement 
assign hkd = ~HKD;  //complement 
assign HLD = ~hld;  //complement 
assign hmc = ~HMC;  //complement 
assign HNC = ~hnc;  //complement 
assign hmd = ~HMD;  //complement 
assign HND = ~hnd;  //complement 
assign hma = ~HMA;  //complement 
assign HNA = ~hna;  //complement 
assign hmb = ~HMB;  //complement 
assign HNB = ~hnb;  //complement 
assign hod = ~HOD;  //complement 
assign HPD = ~hpd;  //complement 
assign hob = ~HOB;  //complement 
assign HPB = ~hpb;  //complement 
assign hme = ~HME;  //complement 
assign HNE = ~hne;  //complement 
assign hmh = ~HMH;  //complement 
assign hmf = ~HMF;  //complement 
assign HNF = ~hnf;  //complement 
assign hmg = ~HMG;  //complement 
assign hoe = ~HOE;  //complement 
assign HPE = ~hpe;  //complement 
assign hoc = ~HOC;  //complement 
assign HPC = ~hpc;  //complement 
assign hoa = ~HOA;  //complement 
assign HPA = ~hpa;  //complement 
assign hof = ~HOF;  //complement 
assign HPF = ~hpf;  //complement 
assign hac = ~HAC;  //complement 
assign HBC = ~hbc;  //complement 
assign hab = ~HAB;  //complement 
assign HBB = ~hbb;  //complement 
assign haa = ~HAA;  //complement 
assign HBA = ~hba;  //complement 
assign hce = ~HCE;  //complement 
assign HDE = ~hde;  //complement 
assign hcf = ~HCF;  //complement 
assign hcb = ~HCB;  //complement 
assign HDB = ~hdb;  //complement 
assign had = ~HAD;  //complement 
assign HBD = ~hbd;  //complement 
assign hcc = ~HCC;  //complement 
assign HDC = ~hdc;  //complement 
assign hcd = ~HCD;  //complement 
assign HDD = ~hdd;  //complement 
assign hca = ~HCA;  //complement 
assign HDA = ~hda;  //complement 
assign hec = ~HEC;  //complement 
assign HFC = ~hfc;  //complement 
assign hea = ~HEA;  //complement 
assign HFA = ~hfa;  //complement 
assign heb = ~HEB;  //complement 
assign HFB = ~hfb;  //complement 
assign hee = ~HEE;  //complement 
assign HFE = ~hfe;  //complement 
assign hed = ~HED;  //complement 
assign HFD = ~hfd;  //complement 
assign heh = ~HEH;  //complement 
assign hef = ~HEF;  //complement 
assign HFF = ~hff;  //complement 
assign heg = ~HEG;  //complement 
assign hqc = ~HQC;  //complement 
assign OHC = ~ohc;  //complement 
assign hga = ~HGA;  //complement 
assign HHA = ~hha;  //complement 
assign hgb = ~HGB;  //complement 
assign HHB = ~hhb;  //complement 
assign hge = ~HGE;  //complement 
assign HHE = ~hhe;  //complement 
assign hgf = ~HGF;  //complement 
assign HHF = ~hhf;  //complement 
assign hgc = ~HGC;  //complement 
assign HHC = ~hhc;  //complement 
assign EBR = DCJ & CAI ; 
assign ebr = ~EBR ; //complement 
assign EDR = DCJ & CAJ ; 
assign edr = ~EDR ;  //complement 
assign EFR = DCJ & CAK ; 
assign efr = ~EFR ;  //complement 
assign EJR = DCJ & CAM; 
assign ejr = ~EJR; 
assign EBS = DCK & CAH ; 
assign ebs = ~EBS ; //complement 
assign EDS = DCK & CAI ; 
assign eds = ~EDS ;  //complement 
assign EFS = DCK & CAJ ; 
assign efs = ~EFS ;  //complement 
assign EJS = DCK & CAL; 
assign ejs = ~EJS; 
assign NCA =  MCA & mba & mcb  |  mca & MBA & mcb  |  mca & mba & MCB  |  MCA & MBA & MCB  ; 
assign nca = ~NCA; //complement 
assign nda =  MCA & mba & mcb  |  mca & MBA & mcb  |  mca & mba & MCB  |  mca & mba & mcb  ; 
assign NDA = ~nda;  //complement 
assign cca = ~CCA;  //complement 
assign cfa = ~CFA;  //complement 
assign ccb = ~CCB;  //complement 
assign cfb = ~CFB;  //complement 
assign EBT = DCL & CAG ; 
assign ebt = ~EBT ; //complement 
assign EDT = DCL & CAH ; 
assign edt = ~EDT ;  //complement 
assign EFT = DCL & CAI ; 
assign eft = ~EFT ;  //complement 
assign EJT = DCL & CAK; 
assign ejt = ~EJT; 
assign EBU = DCM & CAF ; 
assign ebu = ~EBU ; //complement 
assign EDU = DCM & CAG ; 
assign edu = ~EDU ;  //complement 
assign EFU = DCM & CAH ; 
assign efu = ~EFU ;  //complement 
assign EJU = DCM & CAJ; 
assign eju = ~EJU; 
assign ccc = ~CCC;  //complement 
assign cfc = ~CFC;  //complement 
assign ccd = ~CCD;  //complement 
assign cfd = ~CFD;  //complement 
assign EBV = DCN & CAE ; 
assign ebv = ~EBV ; //complement 
assign EDV = DCN & CAF ; 
assign edv = ~EDV ;  //complement 
assign EFV = DCN & CAG ; 
assign efv = ~EFV ;  //complement 
assign EJV = DCN & CAI; 
assign ejv = ~EJV; 
assign ENW = DCO & CAJ ; 
assign enw = ~ENW ; //complement 
assign ELW = DCO & CAI ; 
assign elw = ~ELW ;  //complement 
assign EJW = DCO & CAH ; 
assign ejw = ~EJW ;  //complement 
assign EFW = DCO & CAF; 
assign efw = ~EFW; 
assign NEA =  MDB & meb & mec  |  mdb & MEB & mec  |  mdb & meb & MEC  |  MDB & MEB & MEC  ; 
assign nea = ~NEA; //complement 
assign nfa =  MDB & meb & mec  |  mdb & MEB & mec  |  mdb & meb & MEC  |  mdb & meb & mec  ; 
assign NFA = ~nfa;  //complement 
assign EFX = DCP & CAE ; 
assign efx = ~EFX ; //complement 
assign EJX = DCP & CAG ; 
assign ejx = ~EJX ;  //complement 
assign ELX = DCP & CAH ; 
assign elx = ~ELX ;  //complement 
assign ENX = DCP & CAI; 
assign enx = ~ENX; 
assign EDJ = DCB & CBB ; 
assign edj = ~EDJ ; //complement 
assign EFJ = DCB & CBC ; 
assign efj = ~EFJ ;  //complement 
assign EJJ = DCB & CBE ; 
assign ejj = ~EJJ ;  //complement 
assign ELJ = DCB & CBF; 
assign elj = ~ELJ; 
assign NGA =  MFA & mga & mgb  |  mfa & MGA & mgb  |  mfa & mga & MGB  |  MFA & MGA & MGB  ; 
assign nga = ~NGA; //complement 
assign nha =  MFA & mga & mgb  |  mfa & MGA & mgb  |  mfa & mga & MGB  |  mfa & mga & mgb  ; 
assign NHA = ~nha;  //complement 
assign EHI =  CBE & DFA  ; 
assign ehi = ~EHI;  //complement 
assign EHK = DFC & CBC ; 
assign ehk = ~EHK ; //complement 
assign EPK = DFC & CBG ; 
assign epk = ~EPK ;  //complement 
assign ERK = DFC & CBH ; 
assign erk = ~ERK ;  //complement 
assign NIA =  MIA & mib & mha  |  mia & MIB & mha  |  mia & mib & MHA  |  MIA & MIB & MHA  ; 
assign nia = ~NIA; //complement 
assign nja =  MIA & mib & mha  |  mia & MIB & mha  |  mia & mib & MHA  |  mia & mib & mha  ; 
assign NJA = ~nja;  //complement 
assign EHL = DFD & CBB ; 
assign ehl = ~EHL ; //complement 
assign EPL = DFD & CBF ; 
assign epl = ~EPL ;  //complement 
assign ERL = DFD & CBG ; 
assign erl = ~ERL ;  //complement 
assign EHM = DFE & CBA ; 
assign ehm = ~EHM ; //complement 
assign EPM = DFE & CBE ; 
assign epm = ~EPM ;  //complement 
assign ERM = DFE & CBF ; 
assign erm = ~ERM ;  //complement 
assign NKA =  MKA & mkb & mkc  |  mka & MKB & mkc  |  mka & mkb & MKC  |  MKA & MKB & MKC  ; 
assign nka = ~NKA; //complement 
assign nla =  MKA & mkb & mkc  |  mka & MKB & mkc  |  mka & mkb & MKC  |  mka & mkb & mkc  ; 
assign NLA = ~nla;  //complement 
assign EHN = DFF & CAP ; 
assign ehn = ~EHN ; //complement 
assign EPN = DFF & CBD ; 
assign epn = ~EPN ;  //complement 
assign ERN = DFF & CBE ; 
assign ern = ~ERN ;  //complement 
assign EHO = DFG & CAO ; 
assign eho = ~EHO ; //complement 
assign EPO = DFG & CBC ; 
assign epo = ~EPO ;  //complement 
assign ERO = DFG & CBD ; 
assign ero = ~ERO ;  //complement 
assign NMA =  MMA & mmb & mla  |  mma & MMB & mla  |  mma & mmb & MLA  |  MMA & MMB & MLA  ; 
assign nma = ~NMA; //complement 
assign nna =  MMA & mmb & mla  |  mma & MMB & mla  |  mma & mmb & MLA  |  mma & mmb & mla  ; 
assign NNA = ~nna;  //complement 
assign NOA =  MOA & mob & moc  |  moa & MOB & moc  |  moa & mob & MOC  |  MOA & MOB & MOC  ; 
assign noa = ~NOA; //complement 
assign npa =  MOA & mob & moc  |  moa & MOB & moc  |  moa & mob & MOC  |  moa & mob & moc  ; 
assign NPA = ~npa;  //complement 
assign EHP = DFH & CAN ; 
assign ehp = ~EHP ; //complement 
assign EPP = DFH & CBB ; 
assign epp = ~EPP ;  //complement 
assign ERP = DFH & CBC ; 
assign erp = ~ERP ;  //complement 
assign EHQ = DFI & CAM ; 
assign ehq = ~EHQ ; //complement 
assign EPQ = DFI & CBA ; 
assign epq = ~EPQ ;  //complement 
assign ERQ = DFI & CBB ; 
assign erq = ~ERQ ;  //complement 
assign NAA =  MAA & mac & mad  |  maa & MAC & mad  |  maa & mac & MAD  |  MAA & MAC & MAD  ; 
assign naa = ~NAA; //complement 
assign nba =  MAA & mac & mad  |  maa & MAC & mad  |  maa & mac & MAD  |  maa & mac & mad  ; 
assign NBA = ~nba;  //complement 
assign JOA =  HNB & hoa & hna  |  hnb & HOA & hna  |  hnb & hoa & HNA  |  HNB & HOA & HNA  ; 
assign joa = ~JOA; //complement 
assign jpa =  HNB & hoa & hna  |  hnb & HOA & hna  |  hnb & hoa & HNA  |  hnb & hoa & hna  ; 
assign JPA = ~jpa;  //complement 
assign JMB =  HMC & hld & hmd  |  hmc & HLD & hmd  |  hmc & hld & HMD  |  HMC & HLD & HMD  ; 
assign jmb = ~JMB; //complement 
assign jnb =  HMC & hld & hmd  |  hmc & HLD & hmd  |  hmc & hld & HMD  |  hmc & hld & hmd  ; 
assign JNB = ~jnb;  //complement 
assign JMA =  HMB & hlb & hma  |  hmb & HLB & hma  |  hmb & hlb & HMA  |  HMB & HLB & HMA  ; 
assign jma = ~JMA; //complement 
assign jna =  HMB & hlb & hma  |  hmb & HLB & hma  |  hmb & hlb & HMA  |  hmb & hlb & hma  ; 
assign JNA = ~jna;  //complement 
assign JMD =  HLF & hmg & hmh  |  hlf & HMG & hmh  |  hlf & hmg & HMH  |  HLF & HMG & HMH  ; 
assign jmd = ~JMD; //complement 
assign jnd =  HLF & hmg & hmh  |  hlf & HMG & hmh  |  hlf & hmg & HMH  |  hlf & hmg & hmh  ; 
assign JND = ~jnd;  //complement 
assign JQD =  HPF & hqg & hqf  |  hpf & HQG & hqf  |  hpf & hqg & HQF  |  HPF & HQG & HQF  ; 
assign jqd = ~JQD; //complement 
assign jrd =  HPF & hqg & hqf  |  hpf & HQG & hqf  |  hpf & hqg & HQF  |  hpf & hqg & hqf  ; 
assign JRD = ~jrd;  //complement 
assign JOD =  HOF & hnf & hne  |  hof & HNF & hne  |  hof & hnf & HNE  |  HOF & HNF & HNE  ; 
assign jod = ~JOD; //complement 
assign jpd =  HOF & hnf & hne  |  hof & HNF & hne  |  hof & hnf & HNE  |  hof & hnf & hne  ; 
assign JPD = ~jpd;  //complement 
assign JOC =  HOE & hnc & hod  |  hoe & HNC & hod  |  hoe & hnc & HOD  |  HOE & HNC & HOD  ; 
assign joc = ~JOC; //complement 
assign jpc =  HOE & hnc & hod  |  hoe & HNC & hod  |  hoe & hnc & HOD  |  hoe & hnc & hod  ; 
assign JPC = ~jpc;  //complement 
assign JOB =  HND & hob & hoc  |  hnd & HOB & hoc  |  hnd & hob & HOC  |  HND & HOB & HOC  ; 
assign job = ~JOB; //complement 
assign jpb =  HND & hob & hoc  |  hnd & HOB & hoc  |  hnd & hob & HOC  |  hnd & hob & hoc  ; 
assign JPB = ~jpb;  //complement 
assign JQC =  HQE & hpe & hpd  |  hqe & HPE & hpd  |  hqe & hpe & HPD  |  HQE & HPE & HPD  ; 
assign jqc = ~JQC; //complement 
assign jrc =  HQE & hpe & hpd  |  hqe & HPE & hpd  |  hqe & hpe & HPD  |  hqe & hpe & hpd  ; 
assign JRC = ~jrc;  //complement 
assign JQB =  HQD & hpc & hqc  |  hqd & HPC & hqc  |  hqd & hpc & HQC  |  HQD & HPC & HQC  ; 
assign jqb = ~JQB; //complement 
assign jrb =  HQD & hpc & hqc  |  hqd & HPC & hqc  |  hqd & hpc & HQC  |  hqd & hpc & hqc  ; 
assign JRB = ~jrb;  //complement 
assign JQA =  HQB & hqa & hpa  |  hqb & HQA & hpa  |  hqb & hqa & HPA  |  HQB & HQA & HPA  ; 
assign jqa = ~JQA; //complement 
assign jra =  HQB & hqa & hpa  |  hqb & HQA & hpa  |  hqb & hqa & HPA  |  hqb & hqa & hpa  ; 
assign JRA = ~jra;  //complement 
assign hqb = ~HQB;  //complement 
assign OHB = ~ohb;  //complement 
assign ohg = ~OHG;  //complement 
assign OIG = ~oig;  //complement 
assign hqe = ~HQE;  //complement 
assign OHE = ~ohe;  //complement 
assign hqd = ~HQD;  //complement 
assign OHD = ~ohd;  //complement 
assign hqa = ~HQA;  //complement 
assign OHA = ~oha;  //complement 
assign ohj = ~OHJ;  //complement 
assign ohh = ~OHH;  //complement 
assign OIH = ~oih;  //complement 
assign ohi = ~OHI;  //complement 
assign JAC =  HAF & hag & hae  |  haf & HAG & hae  |  haf & hag & HAE  |  HAF & HAG & HAE  ; 
assign jac = ~JAC; //complement 
assign jbc =  HAF & hag & hae  |  haf & HAG & hae  |  haf & hag & HAE  |  haf & hag & hae  ; 
assign JBC = ~jbc;  //complement 
assign JAB =  HAD & hai & hac  |  had & HAI & hac  |  had & hai & HAC  |  HAD & HAI & HAC  ; 
assign jab = ~JAB; //complement 
assign jbb =  HAD & hai & hac  |  had & HAI & hac  |  had & hai & HAC  |  had & hai & hac  ; 
assign JBB = ~jbb;  //complement 
assign JAA =  HAA & hah & hab  |  haa & HAH & hab  |  haa & hah & HAB  |  HAA & HAH & HAB  ; 
assign jaa = ~JAA; //complement 
assign jba =  HAA & hah & hab  |  haa & HAH & hab  |  haa & hah & HAB  |  haa & hah & hab  ; 
assign JBA = ~jba;  //complement 
assign JCA =  HCB & hba & hca  |  hcb & HBA & hca  |  hcb & hba & HCA  |  HCB & HBA & HCA  ; 
assign jca = ~JCA; //complement 
assign jda =  HCB & hba & hca  |  hcb & HBA & hca  |  hcb & hba & HCA  |  hcb & hba & hca  ; 
assign JDA = ~jda;  //complement 
assign JCC =  HBG & hbf & hcf  |  hbg & HBF & hcf  |  hbg & hbf & HCF  |  HBG & HBF & HCF  ; 
assign jcc = ~JCC; //complement 
assign jdc =  HBG & hbf & hcf  |  hbg & HBF & hcf  |  hbg & hbf & HCF  |  hbg & hbf & hcf  ; 
assign JDC = ~jdc;  //complement 
assign JCD =  HBD & hce & hbe  |  hbd & HCE & hbe  |  hbd & hce & HBE  |  HBD & HCE & HBE  ; 
assign jcd = ~JCD; //complement 
assign jdd =  HBD & hce & hbe  |  hbd & HCE & hbe  |  hbd & hce & HBE  |  hbd & hce & hbe  ; 
assign JDD = ~jdd;  //complement 
assign JCB =  HBC & hcd & hcc  |  hbc & HCD & hcc  |  hbc & hcd & HCC  |  HBC & HCD & HCC  ; 
assign jcb = ~JCB; //complement 
assign jdb =  HBC & hcd & hcc  |  hbc & HCD & hcc  |  hbc & hcd & HCC  |  hbc & hcd & hcc  ; 
assign JDB = ~jdb;  //complement 
assign JEC =  HEF & heh & hdc  |  hef & HEH & hdc  |  hef & heh & HDC  |  HEF & HEH & HDC  ; 
assign jec = ~JEC; //complement 
assign jfc =  HEF & heh & hdc  |  hef & HEH & hdc  |  hef & heh & HDC  |  hef & heh & hdc  ; 
assign JFC = ~jfc;  //complement 
assign JED =  HEE & heg & hde  |  hee & HEG & hde  |  hee & heg & HDE  |  HEE & HEG & HDE  ; 
assign jed = ~JED; //complement 
assign jfd =  HEE & heg & hde  |  hee & HEG & hde  |  hee & heg & HDE  |  hee & heg & hde  ; 
assign JFD = ~jfd;  //complement 
assign JEB =  HED & hdd & hec  |  hed & HDD & hec  |  hed & hdd & HEC  |  HED & HDD & HEC  ; 
assign jeb = ~JEB; //complement 
assign jfb =  HED & hdd & hec  |  hed & HDD & hec  |  hed & hdd & HEC  |  hed & hdd & hec  ; 
assign JFB = ~jfb;  //complement 
assign JEA =  HEB & hdb & hea  |  heb & HDB & hea  |  heb & hdb & HEA  |  HEB & HDB & HEA  ; 
assign jea = ~JEA; //complement 
assign jfa =  HEB & hdb & hea  |  heb & HDB & hea  |  heb & hdb & HEA  |  heb & hdb & hea  ; 
assign JFA = ~jfa;  //complement 
assign JGC =  HGG & hgf & hff  |  hgg & HGF & hff  |  hgg & hgf & HFF  |  HGG & HGF & HFF  ; 
assign jgc = ~JGC; //complement 
assign jhc =  HGG & hgf & hff  |  hgg & HGF & hff  |  hgg & hgf & HFF  |  hgg & hgf & hff  ; 
assign JHC = ~jhc;  //complement 
assign JGD =  HGE & hfe & hfc  |  hge & HFE & hfc  |  hge & hfe & HFC  |  HGE & HFE & HFC  ; 
assign jgd = ~JGD; //complement 
assign jhd =  HGE & hfe & hfc  |  hge & HFE & hfc  |  hge & hfe & HFC  |  hge & hfe & hfc  ; 
assign JHD = ~jhd;  //complement 
assign JGB =  HGD & hfd & hgc  |  hgd & HFD & hgc  |  hgd & hfd & HGC  |  HGD & HFD & HGC  ; 
assign jgb = ~JGB; //complement 
assign jhb =  HGD & hfd & hgc  |  hgd & HFD & hgc  |  hgd & hfd & HGC  |  hgd & hfd & hgc  ; 
assign JHB = ~jhb;  //complement 
assign JGA =  HFB & hgb & hga  |  hfb & HGB & hga  |  hfb & hgb & HGA  |  HFB & HGB & HGA  ; 
assign jga = ~JGA; //complement 
assign jha =  HFB & hgb & hga  |  hfb & HGB & hga  |  hfb & hgb & HGA  |  hfb & hgb & hga  ; 
assign JHA = ~jha;  //complement 
assign JID =  HIE & hhe & hif  |  hie & HHE & hif  |  hie & hhe & HIF  |  HIE & HHE & HIF  ; 
assign jid = ~JID; //complement 
assign jjd =  HIE & hhe & hif  |  hie & HHE & hif  |  hie & hhe & HIF  |  hie & hhe & hif  ; 
assign JJD = ~jjd;  //complement 
assign JIA =  HIB & hhb & hia  |  hib & HHB & hia  |  hib & hhb & HIA  |  HIB & HHB & HIA  ; 
assign jia = ~JIA; //complement 
assign jja =  HIB & hhb & hia  |  hib & HHB & hia  |  hib & hhb & HIA  |  hib & hhb & hia  ; 
assign JJA = ~jja;  //complement 
assign JIB =  HHC & hic & hid  |  hhc & HIC & hid  |  hhc & hic & HID  |  HHC & HIC & HID  ; 
assign jib = ~JIB; //complement 
assign jjb =  HHC & hic & hid  |  hhc & HIC & hid  |  hhc & hic & HID  |  hhc & hic & hid  ; 
assign JJB = ~jjb;  //complement 
assign JKB =  HKC & hkd & hja  |  hkc & HKD & hja  |  hkc & hkd & HJA  |  HKC & HKD & HJA  ; 
assign jkb = ~JKB; //complement 
assign jlb =  HKC & hkd & hja  |  hkc & HKD & hja  |  hkc & hkd & HJA  |  hkc & hkd & hja  ; 
assign JLB = ~jlb;  //complement 
assign JKA =  HKA & hkb & hjb  |  hka & HKB & hjb  |  hka & hkb & HJB  |  HKA & HKB & HJB  ; 
assign jka = ~JKA; //complement 
assign jla =  HKA & hkb & hjb  |  hka & HKB & hjb  |  hka & hkb & HJB  |  hka & hkb & hjb  ; 
assign JLA = ~jla;  //complement 
assign JIC =  HIG & hhg & hhf  |  hig & HHG & hhf  |  hig & hhg & HHF  |  HIG & HHG & HHF  ; 
assign jic = ~JIC; //complement 
assign jjc =  HIG & hhg & hhf  |  hig & HHG & hhf  |  hig & hhg & HHF  |  hig & hhg & hhf  ; 
assign JJC = ~jjc;  //complement 
assign JMC =  HLC & hle & hmf  |  hlc & HLE & hmf  |  hlc & hle & HMF  |  HLC & HLE & HMF  ; 
assign jmc = ~JMC; //complement 
assign jnc =  HLC & hle & hmf  |  hlc & HLE & hmf  |  hlc & hle & HMF  |  hlc & hle & hmf  ; 
assign JNC = ~jnc;  //complement 
assign JKD =  HKF & hkg & hjg  |  hkf & HKG & hjg  |  hkf & hkg & HJG  |  HKF & HKG & HJG  ; 
assign jkd = ~JKD; //complement 
assign jld =  HKF & hkg & hjg  |  hkf & HKG & hjg  |  hkf & hkg & HJG  |  hkf & hkg & hjg  ; 
assign JLD = ~jld;  //complement 
assign JKC =  HKE & hjd & hjc  |  hke & HJD & hjc  |  hke & hjd & HJC  |  HKE & HJD & HJC  ; 
assign jkc = ~JKC; //complement 
assign jlc =  HKE & hjd & hjc  |  hke & HJD & hjc  |  hke & hjd & HJC  |  hke & hjd & hjc  ; 
assign JLC = ~jlc;  //complement 
assign ERR = DFJ & CBA ; 
assign err = ~ERR ; //complement 
assign EPR = DFJ & CAP ; 
assign epr = ~EPR ;  //complement 
assign EHR = DFJ & CAL ; 
assign ehr = ~EHR ;  //complement 
assign EHS = DFK & CAK ; 
assign ehs = ~EHS ; //complement 
assign EPS = DFK & CAO ; 
assign eps = ~EPS ;  //complement 
assign ERS = DFK & CAP ; 
assign ers = ~ERS ;  //complement 
assign cce = ~CCE;  //complement 
assign cfe = ~CFE;  //complement 
assign ccf = ~CCF;  //complement 
assign cff = ~CFF;  //complement 
assign EHT = DFL & CAJ ; 
assign eht = ~EHT ; //complement 
assign EPT = DFL & CAN ; 
assign ept = ~EPT ;  //complement 
assign ERT = DFL & CAO ; 
assign ert = ~ERT ;  //complement 
assign EHU = DFM & CAI ; 
assign ehu = ~EHU ; //complement 
assign EPU = DFM & CAM ; 
assign epu = ~EPU ;  //complement 
assign ERU = DFM & CAN ; 
assign eru = ~ERU ;  //complement 
assign ccg = ~CCG;  //complement 
assign cfg = ~CFG;  //complement 
assign cch = ~CCH;  //complement 
assign cfh = ~CFH;  //complement 
assign EHV =  CAH & DFN  ; 
assign ehv = ~EHV;  //complement 
assign EPV =  CAL & DFN  ; 
assign epv = ~EPV;  //complement 
assign ERV =  CAM & DFN  ; 
assign erv = ~ERV;  //complement 
assign EHW =  CAG & DFO  ; 
assign ehw = ~EHW;  //complement 
assign EPW =  CAK & DFO  ; 
assign epw = ~EPW;  //complement 
assign ERW =  CAL & DFO  ; 
assign erw = ~ERW;  //complement 
assign cci = ~CCI;  //complement 
assign cfi = ~CFI;  //complement 
assign ccj = ~CCJ;  //complement 
assign cfj = ~CFJ;  //complement 
assign EHX = DFP & CAF ; 
assign ehx = ~EHX ; //complement 
assign EPX = DFP & CAJ ; 
assign epx = ~EPX ;  //complement 
assign ERX = DFP & CAK ; 
assign erx = ~ERX ;  //complement 
assign EMK = DGK & CCN ; 
assign emk = ~EMK ; //complement 
assign EOK = DGK & CCO ; 
assign eok = ~EOK ;  //complement 
assign EQK = DGK & CCP ; 
assign eqk = ~EQK ;  //complement 
assign EML = DGL & CCM ; 
assign eml = ~EML ; //complement 
assign EOL = DGL & CCN ; 
assign eol = ~EOL ;  //complement 
assign EQL = DGL & CCO ; 
assign eql = ~EQL ;  //complement 
assign EMM = DGM & CCL ; 
assign emm = ~EMM ; //complement 
assign EOM = DGM & CCM ; 
assign eom = ~EOM ;  //complement 
assign EQM = DGM & CCN ; 
assign eqm = ~EQM ;  //complement 
assign EMN = DGN & CCK ; 
assign emn = ~EMN ; //complement 
assign EON = DGN & CCL ; 
assign eon = ~EON ;  //complement 
assign EQN = DGN & CCM ; 
assign eqn = ~EQN ;  //complement 
assign EMO = DGO & CCJ ; 
assign emo = ~EMO ; //complement 
assign EOO = DGO & CCK ; 
assign eoo = ~EOO ;  //complement 
assign EQO = DGO & CCL ; 
assign eqo = ~EQO ;  //complement 
assign mia = ~MIA;  //complement 
assign MJA = ~mja;  //complement 
assign mib = ~MIB;  //complement 
assign EMP = DGP & CCI ; 
assign emp = ~EMP ; //complement 
assign EOP = DGP & CCJ ; 
assign eop = ~EOP ;  //complement 
assign EQP = DGP & CCK ; 
assign eqp = ~EQP ;  //complement 
assign EMQ = DHA & CCH ; 
assign emq = ~EMQ ; //complement 
assign EOQ = DHA & CCI ; 
assign eoq = ~EOQ ;  //complement 
assign EQQ = DHA & CCJ ; 
assign eqq = ~EQQ ;  //complement 
assign mka = ~MKA;  //complement 
assign MLA = ~mla;  //complement 
assign mkb = ~MKB;  //complement 
assign EMR = DHB & CCG ; 
assign emr = ~EMR ; //complement 
assign EOR = DHB & CCH ; 
assign eor = ~EOR ;  //complement 
assign EQR = DHB & CCI ; 
assign eqr = ~EQR ;  //complement 
assign mma = ~MMA;  //complement 
assign MNA = ~mna;  //complement 
assign mmb = ~MMB;  //complement 
assign EMS = DHC & CCF ; 
assign ems = ~EMS ; //complement 
assign EOS = DHC & CCG ; 
assign eos = ~EOS ;  //complement 
assign EQS = DHC & CCH ; 
assign eqs = ~EQS ;  //complement 
assign kqa = ~KQA;  //complement 
assign OKA = ~oka;  //complement 
assign kqb = ~KQB;  //complement 
assign OKB = ~okb;  //complement 
assign koa = ~KOA;  //complement 
assign KPA = ~kpa;  //complement 
assign kod = ~KOD;  //complement 
assign kob = ~KOB;  //complement 
assign KPB = ~kpb;  //complement 
assign koc = ~KOC;  //complement 
assign LAB =  KAB & kaf & kad  |  kab & KAF & kad  |  kab & kaf & KAD  |  KAB & KAF & KAD  ; 
assign lab = ~LAB; //complement 
assign lbb =  KAB & kaf & kad  |  kab & KAF & kad  |  kab & kaf & KAD  |  kab & kaf & kad  ; 
assign LBB = ~lbb;  //complement 
assign LAA =  KAA & kae & kac  |  kaa & KAE & kac  |  kaa & kae & KAC  |  KAA & KAE & KAC  ; 
assign laa = ~LAA; //complement 
assign lba =  KAA & kae & kac  |  kaa & KAE & kac  |  kaa & kae & KAC  |  kaa & kae & kac  ; 
assign LBA = ~lba;  //complement 
assign okd = ~OKD;  //complement 
assign OLD = ~old;  //complement 
assign oke = ~OKE;  //complement 
assign kqc = ~KQC;  //complement 
assign OKC = ~okc;  //complement 
assign LEA =  KEA & kda & kec  |  kea & KDA & kec  |  kea & kda & KEC  |  KEA & KDA & KEC  ; 
assign lea = ~LEA; //complement 
assign lfa =  KEA & kda & kec  |  kea & KDA & kec  |  kea & kda & KEC  |  kea & kda & kec  ; 
assign LFA = ~lfa;  //complement 
assign LCB =  KCB & kcd & kbb  |  kcb & KCD & kbb  |  kcb & kcd & KBB  |  KCB & KCD & KBB  ; 
assign lcb = ~LCB; //complement 
assign ldb =  KCB & kcd & kbb  |  kcb & KCD & kbb  |  kcb & kcd & KBB  |  kcb & kcd & kbb  ; 
assign LDB = ~ldb;  //complement 
assign LCA =  KCA & kce & kba  |  kca & KCE & kba  |  kca & kce & KBA  |  KCA & KCE & KBA  ; 
assign lca = ~LCA; //complement 
assign lda =  KCA & kce & kba  |  kca & KCE & kba  |  kca & kce & KBA  |  kca & kce & kba  ; 
assign LDA = ~lda;  //complement 
assign LCC =  KBC & kcc & kbd  |  kbc & KCC & kbd  |  kbc & kcc & KBD  |  KBC & KCC & KBD  ; 
assign lcc = ~LCC; //complement 
assign ldc =  KBC & kcc & kbd  |  kbc & KCC & kbd  |  kbc & kcc & KBD  |  kbc & kcc & kbd  ; 
assign LDC = ~ldc;  //complement 
assign LIB =  KHB & kib & kid  |  khb & KIB & kid  |  khb & kib & KID  |  KHB & KIB & KID  ; 
assign lib = ~LIB; //complement 
assign ljb =  KHB & kib & kid  |  khb & KIB & kid  |  khb & kib & KID  |  khb & kib & kid  ; 
assign LJB = ~ljb;  //complement 
assign LGB =  KGB & kfb & kfc  |  kgb & KFB & kfc  |  kgb & kfb & KFC  |  KGB & KFB & KFC  ; 
assign lgb = ~LGB; //complement 
assign lhb =  KGB & kfb & kfc  |  kgb & KFB & kfc  |  kgb & kfb & KFC  |  kgb & kfb & kfc  ; 
assign LHB = ~lhb;  //complement 
assign LGA =  KGA & kfa & kgc  |  kga & KFA & kgc  |  kga & kfa & KGC  |  KGA & KFA & KGC  ; 
assign lga = ~LGA; //complement 
assign lha =  KGA & kfa & kgc  |  kga & KFA & kgc  |  kga & kfa & KGC  |  kga & kfa & kgc  ; 
assign LHA = ~lha;  //complement 
assign LEB =  KEB & kdb & kdc  |  keb & KDB & kdc  |  keb & kdb & KDC  |  KEB & KDB & KDC  ; 
assign leb = ~LEB; //complement 
assign lfb =  KEB & kdb & kdc  |  keb & KDB & kdc  |  keb & kdb & KDC  |  keb & kdb & kdc  ; 
assign LFB = ~lfb;  //complement 
assign LMA =  KMA & kla & kmc  |  kma & KLA & kmc  |  kma & kla & KMC  |  KMA & KLA & KMC  ; 
assign lma = ~LMA; //complement 
assign lna =  KMA & kla & kmc  |  kma & KLA & kmc  |  kma & kla & KMC  |  kma & kla & kmc  ; 
assign LNA = ~lna;  //complement 
assign LKB =  KKB & kkd & kjb  |  kkb & KKD & kjb  |  kkb & kkd & KJB  |  KKB & KKD & KJB  ; 
assign lkb = ~LKB; //complement 
assign llb =  KKB & kkd & kjb  |  kkb & KKD & kjb  |  kkb & kkd & KJB  |  kkb & kkd & kjb  ; 
assign LLB = ~llb;  //complement 
assign LKA =  KKA & kja & kkc  |  kka & KJA & kkc  |  kka & kja & KKC  |  KKA & KJA & KKC  ; 
assign lka = ~LKA; //complement 
assign lla =  KKA & kja & kkc  |  kka & KJA & kkc  |  kka & kja & KKC  |  kka & kja & kkc  ; 
assign LLA = ~lla;  //complement 
assign LIA =  KIA & kha & kic  |  kia & KHA & kic  |  kia & kha & KIC  |  KIA & KHA & KIC  ; 
assign lia = ~LIA; //complement 
assign lja =  KIA & kha & kic  |  kia & KHA & kic  |  kia & kha & KIC  |  kia & kha & kic  ; 
assign LJA = ~lja;  //complement 
assign oab = ~OAB;  //complement 
assign obb = ~OBB;  //complement 
assign oac = ~OAC;  //complement 
assign obc = ~OBC;  //complement 
assign oad = ~OAD;  //complement 
assign obd = ~OBD;  //complement 
assign oaf = ~OAF;  //complement 
assign obf = ~OBF;  //complement 
assign LQA =  KQC & kpa & kpb  |  kqc & KPA & kpb  |  kqc & kpa & KPB  |  KQC & KPA & KPB  ; 
assign lqa = ~LQA; //complement 
assign lra =  KQC & kpa & kpb  |  kqc & KPA & kpb  |  kqc & kpa & KPB  |  kqc & kpa & kpb  ; 
assign LRA = ~lra;  //complement 
assign LOA =  KOC & kod & kna  |  koc & KOD & kna  |  koc & kod & KNA  |  KOC & KOD & KNA  ; 
assign loa = ~LOA; //complement 
assign lpa =  KOC & kod & kna  |  koc & KOD & kna  |  koc & kod & KNA  |  koc & kod & kna  ; 
assign LPA = ~lpa;  //complement 
assign LOB =  KOB & knb & koa  |  kob & KNB & koa  |  kob & knb & KOA  |  KOB & KNB & KOA  ; 
assign lob = ~LOB; //complement 
assign lpb =  KOB & knb & koa  |  kob & KNB & koa  |  kob & knb & KOA  |  kob & knb & koa  ; 
assign LPB = ~lpb;  //complement 
assign LMB =  KMB & klb & kmd  |  kmb & KLB & kmd  |  kmb & klb & KMD  |  KMB & KLB & KMD  ; 
assign lmb = ~LMB; //complement 
assign lnb =  KMB & klb & kmd  |  kmb & KLB & kmd  |  kmb & klb & KMD  |  kmb & klb & kmd  ; 
assign LNB = ~lnb;  //complement 
assign oaa = ~OAA;  //complement 
assign oba = ~OBA;  //complement 
assign oae = ~OAE;  //complement 
assign obe = ~OBE;  //complement 
assign oai = ~OAI;  //complement 
assign obi = ~OBI;  //complement 
assign oam = ~OAM;  //complement 
assign obm = ~OBM;  //complement 
assign kad = ~KAD;  //complement 
assign KBD = ~kbd;  //complement 
assign kae = ~KAE;  //complement 
assign hag = ~HAG;  //complement 
assign HBG = ~hbg;  //complement 
assign hah = ~HAH;  //complement 
assign haf = ~HAF;  //complement 
assign HBF = ~hbf;  //complement 
assign hai = ~HAI;  //complement 
assign kab = ~KAB;  //complement 
assign KBB = ~kbb;  //complement 
assign kac = ~KAC;  //complement 
assign KBC = ~kbc;  //complement 
assign kaf = ~KAF;  //complement 
assign kaa = ~KAA;  //complement 
assign KBA = ~kba;  //complement 
assign kcb = ~KCB;  //complement 
assign KDB = ~kdb;  //complement 
assign kce = ~KCE;  //complement 
assign kca = ~KCA;  //complement 
assign KDA = ~kda;  //complement 
assign kcc = ~KCC;  //complement 
assign KDC = ~kdc;  //complement 
assign kcd = ~KCD;  //complement 
assign kec = ~KEC;  //complement 
assign KFC = ~kfc;  //complement 
assign kea = ~KEA;  //complement 
assign KFA = ~kfa;  //complement 
assign keb = ~KEB;  //complement 
assign KFB = ~kfb;  //complement 
assign kgc = ~KGC;  //complement 
assign KHC = ~khc;  //complement 
assign kga = ~KGA;  //complement 
assign KHA = ~kha;  //complement 
assign kgb = ~KGB;  //complement 
assign KHB = ~khb;  //complement 
assign kib = ~KIB;  //complement 
assign KJB = ~kjb;  //complement 
assign kia = ~KIA;  //complement 
assign KJA = ~kja;  //complement 
assign kic = ~KIC;  //complement 
assign KJC = ~kjc;  //complement 
assign kid = ~KID;  //complement 
assign kka = ~KKA;  //complement 
assign KLA = ~kla;  //complement 
assign kkb = ~KKB;  //complement 
assign KLB = ~klb;  //complement 
assign kkc = ~KKC;  //complement 
assign KLC = ~klc;  //complement 
assign kkd = ~KKD;  //complement 
assign kmb = ~KMB;  //complement 
assign KNB = ~knb;  //complement 
assign kmc = ~KMC;  //complement 
assign KNC = ~knc;  //complement 
assign kmd = ~KMD;  //complement 
assign kma = ~KMA;  //complement 
assign KNA = ~kna;  //complement 
assign mqa = ~MQA;  //complement 
assign OMA = ~oma;  //complement 
assign mqb = ~MQB;  //complement 
assign EMU = DHE & CCD ; 
assign emu = ~EMU ; //complement 
assign EOU = DHE & CCE ; 
assign eou = ~EOU ;  //complement 
assign EQU = DHE & CCF ; 
assign equ = ~EQU ;  //complement 
assign oak = ~OAK;  //complement 
assign obk = ~OBK;  //complement 
assign cck = ~CCK;  //complement 
assign cfk = ~CFK;  //complement 
assign ccl = ~CCL;  //complement 
assign cfl = ~CFL;  //complement 
assign EMV = DHF & CCC ; 
assign emv = ~EMV ; //complement 
assign EOV = DHF & CCD ; 
assign eov = ~EOV ;  //complement 
assign EQV = DHF & CCE ; 
assign eqv = ~EQV ;  //complement 
assign EMW = DHG & CCB ; 
assign emw = ~EMW ; //complement 
assign EOW = DHG & CCC ; 
assign eow = ~EOW ;  //complement 
assign EQW = DHG & CCD ; 
assign eqw = ~EQW ;  //complement 
assign moa = ~MOA;  //complement 
assign MPA = ~mpa;  //complement 
assign mob = ~MOB;  //complement 
assign ccm = ~CCM;  //complement 
assign cfm = ~CFM;  //complement 
assign ccn = ~CCN;  //complement 
assign cfn = ~CFN;  //complement 
assign EMX = DHH & CCA ; 
assign emx = ~EMX ; //complement 
assign EOX = DHH & CCB ; 
assign eox = ~EOX ;  //complement 
assign EQX = DHH & CCC ; 
assign eqx = ~EQX ;  //complement 
assign ENA = DHI & CBP ; 
assign ena = ~ENA ; //complement 
assign EPA = DHI & CCA ; 
assign epa = ~EPA ;  //complement 
assign ERA = DHI & CCB ; 
assign era = ~ERA ;  //complement 
assign maa = ~MAA;  //complement 
assign MBA = ~mba;  //complement 
assign mac = ~MAC;  //complement 
assign cco = ~CCO;  //complement 
assign cfo = ~CFO;  //complement 
assign ccp = ~CCP;  //complement 
assign cfp = ~CFP;  //complement 
assign ENB = DHJ & CBO ; 
assign enb = ~ENB ; //complement 
assign EPB = DHJ & CBP ; 
assign epb = ~EPB ;  //complement 
assign ERB = DHJ & CCA ; 
assign erb = ~ERB ;  //complement 
assign ENC = DHK & CBN ; 
assign enc = ~ENC ; //complement 
assign EPC = DHK & CBO ; 
assign epc = ~EPC ;  //complement 
assign ERC = DHK & CBP ; 
assign erc = ~ERC ;  //complement 
assign mab = ~MAB;  //complement 
assign MBB = ~mbb;  //complement 
assign mad = ~MAD;  //complement 
assign ENDD  = DHL & CBM ; 
assign endd = ~ENDD  ; //complement 
assign EPD = DHL & CBN ; 
assign epd = ~EPD ;  //complement 
assign ERD = DHL & CBO ; 
assign erd = ~ERD ;  //complement 
assign mca = ~MCA;  //complement 
assign MDA = ~mda;  //complement 
assign ENE = DHM & CBL ; 
assign ene = ~ENE ; //complement 
assign EPE = DHM & CBM ; 
assign epe = ~EPE ;  //complement 
assign ERE = DHM & CBN ; 
assign ere = ~ERE ;  //complement 
assign oao = ~OAO;  //complement 
assign obo = ~OBO;  //complement 
assign oap = ~OAP;  //complement 
assign obp = ~OBP;  //complement 
assign mcb = ~MCB;  //complement 
assign MDB = ~mdb;  //complement 
assign ENG = DHO & CBJ ; 
assign eng = ~ENG ; //complement 
assign EPG = DHO & CBK ; 
assign epg = ~EPG ;  //complement 
assign ERG = DHO & CBL ; 
assign erg = ~ERG ;  //complement 
assign oal = ~OAL;  //complement 
assign obl = ~OBL;  //complement 
assign oan = ~OAN;  //complement 
assign obn = ~OBN;  //complement 
assign ENH = DHP & CBI ; 
assign enh = ~ENH ; //complement 
assign EPH = DHP & CBJ ; 
assign eph = ~EPH ;  //complement 
assign ERH = DHP & CBK ; 
assign erh = ~ERH ;  //complement 
assign oag = ~OAG;  //complement 
assign obg = ~OBG;  //complement 
assign ENF = DHN & CBK ; 
assign enf = ~ENF ; //complement 
assign EPF = DHN & CBL ; 
assign epf = ~EPF ;  //complement 
assign ERF = DHN & CBM ; 
assign erf = ~ERF ;  //complement 
assign mea = ~MEA;  //complement 
assign MFA = ~mfa;  //complement 
assign mga = ~MGA;  //complement 
assign MHA = ~mha;  //complement 
assign mgb = ~MGB;  //complement 
assign oah = ~OAH;  //complement 
assign obh = ~OBH;  //complement 
assign EMT = DHD & CCE ; 
assign emt = ~EMT ; //complement 
assign EOT = DHD & CCF ; 
assign eot = ~EOT ;  //complement 
assign EQT = DHD & CCG ; 
assign eqt = ~EQT ;  //complement 
assign oaj = ~OAJ;  //complement 
assign obj = ~OBJ;  //complement 
assign iba = ~IBA; //complement 
assign ibb = ~IBB; //complement 
assign ibc = ~IBC; //complement 
assign ibd = ~IBD; //complement 
assign ibe = ~IBE; //complement 
assign ibf = ~IBF; //complement 
assign ibg = ~IBG; //complement 
assign ibh = ~IBH; //complement 
assign ibi = ~IBI; //complement 
assign ibj = ~IBJ; //complement 
assign ibk = ~IBK; //complement 
assign ibl = ~IBL; //complement 
assign ibm = ~IBM; //complement 
assign ibn = ~IBN; //complement 
assign ibo = ~IBO; //complement 
assign ibp = ~IBP; //complement 
assign ica = ~ICA; //complement 
assign icb = ~ICB; //complement 
assign icc = ~ICC; //complement 
assign icd = ~ICD; //complement 
assign ice = ~ICE; //complement 
assign icf = ~ICF; //complement 
assign icg = ~ICG; //complement 
assign ich = ~ICH; //complement 
assign ici = ~ICI; //complement 
assign icj = ~ICJ; //complement 
assign ick = ~ICK; //complement 
assign icl = ~ICL; //complement 
assign icm = ~ICM; //complement 
assign icn = ~ICN; //complement 
assign ico = ~ICO; //complement 
assign icp = ~ICP; //complement 
assign ida = ~IDA; //complement 
assign idb = ~IDB; //complement 
assign idc = ~IDC; //complement 
assign idd = ~IDD; //complement 
assign ide = ~IDE; //complement 
assign idf = ~IDF; //complement 
assign idg = ~IDG; //complement 
assign idh = ~IDH; //complement 
assign idi = ~IDI; //complement 
assign idj = ~IDJ; //complement 
assign idk = ~IDK; //complement 
assign idl = ~IDL; //complement 
assign idm = ~IDM; //complement 
assign idn = ~IDN; //complement 
assign ido = ~IDO; //complement 
assign idp = ~IDP; //complement 
assign iea = ~IEA; //complement 
assign ieb = ~IEB; //complement 
assign iec = ~IEC; //complement 
assign ied = ~IED; //complement 
assign iee = ~IEE; //complement 
assign ief = ~IEF; //complement 
assign ieg = ~IEG; //complement 
assign ieh = ~IEH; //complement 
assign iei = ~IEI; //complement 
assign iej = ~IEJ; //complement 
assign iek = ~IEK; //complement 
assign iel = ~IEL; //complement 
assign iem = ~IEM; //complement 
assign ien = ~IEN; //complement 
assign ieo = ~IEO; //complement 
assign iep = ~IEP; //complement 
assign ieq = ~IEQ; //complement 
assign ier = ~IER; //complement 
assign ies = ~IES; //complement 
assign iet = ~IET; //complement 
assign ieu = ~IEU; //complement 
assign iev = ~IEV; //complement 
assign iew = ~IEW; //complement 
assign iex = ~IEX; //complement 
assign iey = ~IEY; //complement 
assign iez = ~IEZ; //complement 
assign ifa = ~IFA; //complement 
assign ifb = ~IFB; //complement 
assign ifc = ~IFC; //complement 
assign ifd = ~IFD; //complement 
assign ife = ~IFE; //complement 
assign ifff  = ~IFFF ; //complement 
assign ifg = ~IFG; //complement 
assign ifh = ~IFH; //complement 
assign ifi = ~IFI; //complement 
assign ifj = ~IFJ; //complement 
assign ifk = ~IFK; //complement 
assign ifl = ~IFL; //complement 
assign ifm = ~IFM; //complement 
assign ifn = ~IFN; //complement 
assign ifo = ~IFO; //complement 
assign ifp = ~IFP; //complement 
assign iga = ~IGA; //complement 
assign igb = ~IGB; //complement 
assign igc = ~IGC; //complement 
assign igd = ~IGD; //complement 
assign ige = ~IGE; //complement 
assign igf = ~IGF; //complement 
assign igg = ~IGG; //complement 
assign igh = ~IGH; //complement 
assign igi = ~IGI; //complement 
assign igj = ~IGJ; //complement 
assign igk = ~IGK; //complement 
assign igl = ~IGL; //complement 
assign igm = ~IGM; //complement 
assign ign = ~IGN; //complement 
assign igo = ~IGO; //complement 
assign igp = ~IGP; //complement 
assign iha = ~IHA; //complement 
assign iia = ~IIA; //complement 
assign ika = ~IKA; //complement 
assign ila = ~ILA; //complement 
assign ilb = ~ILB; //complement 
assign ilc = ~ILC; //complement 
assign ild = ~ILD; //complement 
assign ile = ~ILE; //complement 
assign ilf = ~ILF; //complement 
assign ilg = ~ILG; //complement 
assign ilh = ~ILH; //complement 
assign ili = ~ILI; //complement 
assign ilj = ~ILJ; //complement 
assign ilk = ~ILK; //complement 
assign ill = ~ILL; //complement 
assign ilm = ~ILM; //complement 
assign iln = ~ILN; //complement 
assign ilo = ~ILO; //complement 
assign ilp = ~ILP; //complement 
assign ima = ~IMA; //complement 
assign imb = ~IMB; //complement 
assign imc = ~IMC; //complement 
assign imd = ~IMD; //complement 
assign ime = ~IME; //complement 
assign imf = ~IMF; //complement 
assign img = ~IMG; //complement 
assign imh = ~IMH; //complement 
assign imi = ~IMI; //complement 
assign imj = ~IMJ; //complement 
assign imk = ~IMK; //complement 
assign iml = ~IML; //complement 
assign imm = ~IMM; //complement 
assign imn = ~IMN; //complement 
assign ina = ~INA; //complement 
assign inb = ~INB; //complement 
assign inc = ~INC; //complement 
assign ind = ~IND; //complement 
assign ine = ~INE; //complement 
assign inf = ~INF; //complement 
assign ing = ~ING; //complement 
assign ioa = ~IOA; //complement 
assign iob = ~IOB; //complement 
assign ioc = ~IOC; //complement 
assign ira = ~IRA; //complement 
assign isa = ~ISA; //complement 
assign ita = ~ITA; //complement 
assign itb = ~ITB; //complement 
always@(posedge IZZ )
   begin 
 FAE <=  EBJ & ebk & ebl  |  ebj & EBK & ebl  |  ebj & ebk & EBL  |  EBJ & EBK & EBL  ;
 fbe <=  EBJ & ebk & ebl  |  ebj & EBK & ebl  |  ebj & ebk & EBL  |  ebj & ebk & ebl  ;
 FAF <=  EBG & ebh & ebi  |  ebg & EBH & ebi  |  ebg & ebh & EBI  |  EBG & EBH & EBI  ;
 fbf <=  EBG & ebh & ebi  |  ebg & EBH & ebi  |  ebg & ebh & EBI  |  ebg & ebh & ebi  ;
 FAG <=  EBD & ebe & ebf  |  ebd & EBE & ebf  |  ebd & ebe & EBF  |  EBD & EBE & EBF  ;
 fbg <=  EBD & ebe & ebf  |  ebd & EBE & ebf  |  ebd & ebe & EBF  |  ebd & ebe & ebf  ;
 FAH <=  EBA & ebb & ebc  |  eba & EBB & ebc  |  eba & ebb & EBC  |  EBA & EBB & EBC  ;
 fbh <=  EBA & ebb & ebc  |  eba & EBB & ebc  |  eba & ebb & EBC  |  eba & ebb & ebc  ;
 AAB <=  ICB & TSA  |  BAB & TKA  |  AAB & THA  ; 
 FAB <=  EBS & ebt & ebu  |  ebs & EBT & ebu  |  ebs & ebt & EBU  |  EBS & EBT & EBU  ;
 fbb <=  EBS & ebt & ebu  |  ebs & EBT & ebu  |  ebs & ebt & EBU  |  ebs & ebt & ebu  ;
 FAC <=  EBP & ebq & ebr  |  ebp & EBQ & ebr  |  ebp & ebq & EBR  |  EBP & EBQ & EBR  ;
 fbc <=  EBP & ebq & ebr  |  ebp & EBQ & ebr  |  ebp & ebq & EBR  |  ebp & ebq & ebr  ;
 FAD <=  EBM & ebn & ebo  |  ebm & EBN & ebo  |  ebm & ebn & EBO  |  EBM & EBN & EBO  ;
 fbd <=  EBM & ebn & ebo  |  ebm & EBN & ebo  |  ebm & ebn & EBO  |  ebm & ebn & ebo  ;
 FCD <=  EDM & edn & edo  |  edm & EDN & edo  |  edm & edn & EDO  |  EDM & EDN & EDO  ;
 fdd <=  EDM & edn & edo  |  edm & EDN & edo  |  edm & edn & EDO  |  edm & edn & edo  ;
 FCE <=  EDJ & edk & edl  |  edj & EDK & edl  |  edj & edk & EDL  |  EDJ & EDK & EDL  ;
 fde <=  EDJ & edk & edl  |  edj & EDK & edl  |  edj & edk & EDL  |  edj & edk & edl  ;
 FCF <=  EDG & edh & edi  |  edg & EDH & edi  |  edg & edh & EDI  |  EDG & EDH & EDI  ;
 fdf <=  EDG & edh & edi  |  edg & EDH & edi  |  edg & edh & EDI  |  edg & edh & edi  ;
 FCG <=  EDD & ede & edf  |  edd & EDE & edf  |  edd & ede & EDF  |  EDD & EDE & EDF  ;
 fdg <=  EDD & ede & edf  |  edd & EDE & edf  |  edd & ede & EDF  |  edd & ede & edf  ;
 AAC <=  ICC & TSB  |  BAC & TKB  |  AAC & THB  ; 
 FCA <=  EDX & edw & edv  |  edx & EDW & edv  |  edx & edw & EDV  |  EDX & EDW & EDV  ;
 fda <=  EDX & edw & edv  |  edx & EDW & edv  |  edx & edw & EDV  |  edx & edw & edv  ;
 FCB <=  EDS & edt & edu  |  eds & EDT & edu  |  eds & edt & EDU  |  EDS & EDT & EDU  ;
 fdb <=  EDS & edt & edu  |  eds & EDT & edu  |  eds & edt & EDU  |  eds & edt & edu  ;
 FCC <=  EDP & edq & edr  |  edp & EDQ & edr  |  edp & edq & EDR  |  EDP & EDQ & EDR  ;
 fdc <=  EDP & edq & edr  |  edp & EDQ & edr  |  edp & edq & EDR  |  edp & edq & edr  ;
 AAD <=  ICD & TSB  |  BAD & TKB  |  AAD & THB  ; 
 AAE <=  ICE & TSA  |  BAE & TKA  |  AAE & THA  ; 
 AAF <=  ICF & TSA  |  BAF & TKA  |  AAF & THA  ; 
 AAG <=  ICG & TSB  |  BAG & TKB  |  AAG & THB  ; 
 FEC <=  EFP & efq & efr  |  efp & EFQ & efr  |  efp & efq & EFR  |  EFP & EFQ & EFR  ;
 ffc <=  EFP & efq & efr  |  efp & EFQ & efr  |  efp & efq & EFR  |  efp & efq & efr  ;
 FED <=  EFM & efn & efo  |  efm & EFN & efo  |  efm & efn & EFO  |  EFM & EFN & EFO  ;
 ffd <=  EFM & efn & efo  |  efm & EFN & efo  |  efm & efn & EFO  |  efm & efn & efo  ;
 FEE <=  EFJ & efk & efl  |  efj & EFK & efl  |  efj & efk & EFL  |  EFJ & EFK & EFL  ;
 ffe <=  EFJ & efk & efl  |  efj & EFK & efl  |  efj & efk & EFL  |  efj & efk & efl  ;
 FEF <=  EFG & efh & efi  |  efg & EFH & efi  |  efg & efh & EFI  |  EFG & EFH & EFI  ;
 fff <=  EFG & efh & efi  |  efg & EFH & efi  |  efg & efh & EFI  |  efg & efh & efi  ;
 oda <= ida ; 
 odb <= idb ; 
 odc <= idc ; 
 odd <= idd ; 
 ode <= ide ; 
 odf <= idf ; 
 odg <= idg ; 
 odh <= idh ; 
 FEA <=  EFX & efw & efv  |  efx & EFW & efv  |  efx & efw & EFV  |  EFX & EFW & EFV  ;
 ffa <=  EFX & efw & efv  |  efx & EFW & efv  |  efx & efw & EFV  |  efx & efw & efv  ;
 FEB <=  EFS & eft & efu  |  efs & EFT & efu  |  efs & eft & EFU  |  EFS & EFT & EFU  ;
 ffb <=  EFS & eft & efu  |  efs & EFT & efu  |  efs & eft & EFU  |  efs & eft & efu  ;
 odi <= idi ; 
 odj <= idj ; 
 odk <= idk ; 
 odl <= idl ; 
 odm <= idm ; 
 odn <= idn ; 
 odo <= ido ; 
 odp <= idp ; 
 AAA <=  ICA & TSA  |  BAA & TKA  |  AAA & THA  ; 
 FAM <=  EAL & eak & eaj  |  eal & EAK & eaj  |  eal & eak & EAJ  |  EAL & EAK & EAJ  ;
 fbm <=  EAL & eak & eaj  |  eal & EAK & eaj  |  eal & eak & EAJ  |  eal & eak & eaj  ;
 QHA <= IHA ; 
 THA <= QHA ; 
 THB <= QHA ; 
 THC <= QHA ; 
 FAN <=  EAI & eah & eag  |  eai & EAH & eag  |  eai & eah & EAG  |  EAI & EAH & EAG  ;
 fbn <=  EAI & eah & eag  |  eai & EAH & eag  |  eai & eah & EAG  |  eai & eah & eag  ;
 FAQ <= QIC ; 
 FAO <=  EAF & eae & ead  |  eaf & EAE & ead  |  eaf & eae & EAD  |  EAF & EAE & EAD  ;
 fbo <=  EAF & eae & ead  |  eaf & EAE & ead  |  eaf & eae & EAD  |  eaf & eae & ead  ;
 FAP <= EAC ; 
 FAJ <=  EAS & eat & eau  |  eas & EAT & eau  |  eas & eat & EAU  |  EAS & EAT & EAU  ;
 fbj <=  EAS & eat & eau  |  eas & EAT & eau  |  eas & eat & EAU  |  eas & eat & eau  ;
 THD <= QHA ; 
 THE <= QHA ; 
 THF <= QHA ; 
 FAK <=  EAP & eaq & ear  |  eap & EAQ & ear  |  eap & eaq & EAR  |  EAP & EAQ & EAR  ;
 fbk <=  EAP & eaq & ear  |  eap & EAQ & ear  |  eap & eaq & EAR  |  eap & eaq & ear  ;
 FAL <=  EAM & ean & eao  |  eam & EAN & eao  |  eam & ean & EAO  |  EAM & EAN & EAO  ;
 fbl <=  EAM & ean & eao  |  eam & EAN & eao  |  eam & ean & EAO  |  eam & ean & eao  ;
 FCN <=  ECI & ech & ecg  |  eci & ECH & ecg  |  eci & ech & ECG  |  ECI & ECH & ECG  ;
 fdn <=  ECI & ech & ecg  |  eci & ECH & ecg  |  eci & ech & ECG  |  eci & ech & ecg  ;
 FCO <=  ECF & ece & qic  |  ecf & ECE & qic  |  ecf & ece & QIC  |  ECF & ECE & QIC  ;
 fdo <=  ECF & ece & qic  |  ecf & ECE & qic  |  ecf & ece & QIC  |  ecf & ece & qic  ;
 FCP <= ECD ; 
 FAA <=  EBX & ebw & ebv  |  ebx & EBW & ebv  |  ebx & ebw & EBV  |  EBX & EBW & EBV  ;
 fba <=  EBX & ebw & ebv  |  ebx & EBW & ebv  |  ebx & ebw & EBV  |  ebx & ebw & ebv  ;
 FAI <=  EAX & eaw & eav  |  eax & EAW & eav  |  eax & eaw & EAV  |  EAX & EAW & EAV  ;
 fbi <=  EAX & eaw & eav  |  eax & EAW & eav  |  eax & eaw & EAV  |  eax & eaw & eav  ;
 FCK <=  ECP & ecq & ecr  |  ecp & ECQ & ecr  |  ecp & ecq & ECR  |  ECP & ECQ & ECR  ;
 fdk <=  ECP & ecq & ecr  |  ecp & ECQ & ecr  |  ecp & ecq & ECR  |  ecp & ecq & ecr  ;
 FCL <=  ECM & ecn & eco  |  ecm & ECN & eco  |  ecm & ecn & ECO  |  ECM & ECN & ECO  ;
 fdl <=  ECM & ecn & eco  |  ecm & ECN & eco  |  ecm & ecn & ECO  |  ecm & ecn & eco  ;
 FCM <=  ECL & eck & ecj  |  ecl & ECK & ecj  |  ecl & eck & ECJ  |  ECL & ECK & ECJ  ;
 fdm <=  ECL & eck & ecj  |  ecl & ECK & ecj  |  ecl & eck & ECJ  |  ecl & eck & ecj  ;
 FCH <=  EDA & edb & edc  |  eda & EDB & edc  |  eda & edb & EDC  |  EDA & EDB & EDC  ;
 fdh <=  EDA & edb & edc  |  eda & EDB & edc  |  eda & edb & EDC  |  eda & edb & edc  ;
 FCI <=  ECX & ecw & ecv  |  ecx & ECW & ecv  |  ecx & ecw & ECV  |  ECX & ECW & ECV  ;
 fdi <=  ECX & ecw & ecv  |  ecx & ECW & ecv  |  ecx & ecw & ECV  |  ecx & ecw & ecv  ;
 FCJ <=  ECS & ect & ecu  |  ecs & ECT & ecu  |  ecs & ect & ECU  |  ECS & ECT & ECU  ;
 fdj <=  ECS & ect & ecu  |  ecs & ECT & ecu  |  ecs & ect & ECU  |  ecs & ect & ecu  ;
 FEM <=  EEL & eek & eej  |  eel & EEK & eej  |  eel & eek & EEJ  |  EEL & EEK & EEJ  ;
 ffm <=  EEL & eek & eej  |  eel & EEK & eej  |  eel & eek & EEJ  |  eel & eek & eej  ;
 TSA <= QAA ; 
 TSB <= QAA ; 
 TSC <= QAA ; 
 TSD <= QAA ; 
 FEN <=  EEI & eeh & eeg  |  eei & EEH & eeg  |  eei & eeh & EEG  |  EEI & EEH & EEG  ;
 ffn <=  EEI & eeh & eeg  |  eei & EEH & eeg  |  eei & eeh & EEG  |  eei & eeh & eeg  ;
 FEO <=  EEF & eee & qic  |  eef & EEE & qic  |  eef & eee & QIC  |  EEF & EEE & QIC  ;
 ffo <=  EEF & eee & qic  |  eef & EEE & qic  |  eef & eee & QIC  |  eef & eee & qic  ;
 FEJ <=  EES & eet & eeu  |  ees & EET & eeu  |  ees & eet & EEU  |  EES & EET & EEU  ;
 ffj <=  EES & eet & eeu  |  ees & EET & eeu  |  ees & eet & EEU  |  ees & eet & eeu  ;
 TRA <= QTB ; 
 TRB <= QTB ; 
 QTB <= IRA ; 
 FEK <=  EEP & eeq & eer  |  eep & EEQ & eer  |  eep & eeq & EER  |  EEP & EEQ & EER  ;
 ffk <=  EEP & eeq & eer  |  eep & EEQ & eer  |  eep & eeq & EER  |  eep & eeq & eer  ;
 FEL <=  EEM & een & eeo  |  eem & EEN & eeo  |  eem & een & EEO  |  EEM & EEN & EEO  ;
 ffl <=  EEM & een & eeo  |  eem & EEN & eeo  |  eem & een & EEO  |  eem & een & eeo  ;
 FEG <=  EFD & efe & eff  |  efd & EFE & eff  |  efd & efe & EFF  |  EFD & EFE & EFF  ;
 ffg <=  EFD & efe & eff  |  efd & EFE & eff  |  efd & efe & EFF  |  efd & efe & eff  ;
 MQC <= LPB ; 
 MOC <= LNA ; 
 MMC <= LLB ; 
 OMB <= LRA ; 
 FEH <=  EFA & efb & efc  |  efa & EFB & efc  |  efa & efb & EFC  |  EFA & EFB & EFC  ;
 ffh <=  EFA & efb & efc  |  efa & EFB & efc  |  efa & efb & EFC  |  efa & efb & efc  ;
 FEI <=  EEX & eew & eev  |  eex & EEW & eev  |  eex & eew & EEV  |  EEX & EEW & EEV  ;
 ffi <=  EEX & eew & eev  |  eex & EEW & eev  |  eex & eew & EEV  |  eex & eew & eev  ;
 DHA <= IFA ; 
 DHB <= IFB ; 
 DHC <= IFC ; 
 DHD <= IFD ; 
 CAC <= AAC ; 
 CDC <= AAC ; 
 CAD <= AAD ; 
 CDD <= AAD ; 
 DHE <= IFE ; 
 DHF <= IFFF  ; 
 DHG <= IFG ; 
 DHH <= IFH ; 
 CAE <= AAE ; 
 CDE <= AAE ; 
 CAH <= AAH ; 
 QAA <= ISA ; 
 DHI <= IFI ; 
 DHJ <= IFJ ; 
 DHK <= IFK ; 
 DHL <= IFL ; 
 CAG <= AAG ; 
 CDG <= AAG ; 
 TSE <= QAA ; 
 DGA <= BAA ; 
 DGB <= BAB ; 
 DGC <= BAC ; 
 DGD <= BAD ; 
 DAC <= BAC ; 
 DAD <= BAD ; 
 DAE <= BAE ; 
 DAF <= BAF ; 
 DHM <= IFM ; 
 DHN <= IFN ; 
 DHO <= IFO ; 
 DHP <= IFP ; 
 DAH <= BAH ; 
 ddh <= bah ; 
 DAG <= BAG ; 
 ddg <= bag ; 
 ddf <= baf ; 
 CDH <= AAH ; 
 TSF <= QAA ; 
 DAI <= BAI ; 
 ddi <= bai ; 
 DAJ <= BAJ ; 
 ddj <= baj ; 
 MKC <= LJB ; 
 MIC <= LHB ; 
 MEB <= LDB ; 
 MEC <= LEB ; 
 DAK <= BAK ; 
 ddk <= bak ; 
 DAL <= BAL ; 
 ddl <= bal ; 
 DAO <= BAO ; 
 ddo <= bao ; 
 DAP <= BAP ; 
 ddp <= bap ; 
 DAM <= BAM ; 
 ddm <= bam ; 
 DAN <= BAN ; 
 ddn <= ban ; 
 FGB <=  EHS & eht & ehu  |  ehs & EHT & ehu  |  ehs & eht & EHU  |  EHS & EHT & EHU  ;
 fhb <=  EHS & eht & ehu  |  ehs & EHT & ehu  |  ehs & eht & EHU  |  ehs & eht & ehu  ;
 FGC <=  EHP & ehq & ehr  |  ehp & EHQ & ehr  |  ehp & ehq & EHR  |  EHP & EHQ & EHR  ;
 fhc <=  EHP & ehq & ehr  |  ehp & EHQ & ehr  |  ehp & ehq & EHR  |  ehp & ehq & ehr  ;
 FGD <=  EHM & ehn & eho  |  ehm & EHN & eho  |  ehm & ehn & EHO  |  EHM & EHN & EHO  ;
 fhd <=  EHM & ehn & eho  |  ehm & EHN & eho  |  ehm & ehn & EHO  |  ehm & ehn & eho  ;
 FGE <=  EHJ & ehk & ehl  |  ehj & EHK & ehl  |  ehj & ehk & EHL  |  EHJ & EHK & EHL  ;
 fhe <=  EHJ & ehk & ehl  |  ehj & EHK & ehl  |  ehj & ehk & EHL  |  ehj & ehk & ehl  ;
 FIC <=  EJP & ejq & ejr  |  ejp & EJQ & ejr  |  ejp & ejq & EJR  |  EJP & EJQ & EJR  ;
 fjc <=  EJP & ejq & ejr  |  ejp & EJQ & ejr  |  ejp & ejq & EJR  |  ejp & ejq & ejr  ;
 FID <=  EJM & ejn & ejo  |  ejm & EJN & ejo  |  ejm & ejn & EJO  |  EJM & EJN & EJO  ;
 fjd <=  EJM & ejn & ejo  |  ejm & EJN & ejo  |  ejm & ejn & EJO  |  ejm & ejn & ejo  ;
 FIE <=  EJJ & ejk & ejl  |  ejj & EJK & ejl  |  ejj & ejk & EJL  |  EJJ & EJK & EJL  ;
 fje <=  EJJ & ejk & ejl  |  ejj & EJK & ejl  |  ejj & ejk & EJL  |  ejj & ejk & ejl  ;
 FGA <=  EHX & ehw & ehv  |  ehx & EHW & ehv  |  ehx & ehw & EHV  |  EHX & EHW & EHV  ;
 fha <=  EHX & ehw & ehv  |  ehx & EHW & ehv  |  ehx & ehw & EHV  |  ehx & ehw & ehv  ;
 FIB <=  EJS & ejt & eju  |  ejs & EJT & eju  |  ejs & ejt & EJU  |  EJS & EJT & EJU  ;
 fjb <=  EJS & ejt & eju  |  ejs & EJT & eju  |  ejs & ejt & EJU  |  ejs & ejt & eju  ;
 FKH <=  ELA & elb & elc  |  ela & ELB & elc  |  ela & elb & ELC  |  ELA & ELB & ELC  ;
 flh <=  ELA & elb & elc  |  ela & ELB & elc  |  ela & elb & ELC  |  ela & elb & elc  ;
 FIA <=  EJX & ejw & ejv  |  ejx & EJW & ejv  |  ejx & ejw & EJV  |  EJX & EJW & EJV  ;
 fja <=  EJX & ejw & ejv  |  ejx & EJW & ejv  |  ejx & ejw & EJV  |  ejx & ejw & ejv  ;
 FKG <=  ELD & ele & elf  |  eld & ELE & elf  |  eld & ele & ELF  |  ELD & ELE & ELF  ;
 flg <=  ELD & ele & elf  |  eld & ELE & elf  |  eld & ele & ELF  |  eld & ele & elf  ;
 AAL <=  ICL & TSB  |  BAL & TKB  |  AAL & THB  ; 
 FKC <=  ELP & elq & elr  |  elp & ELQ & elr  |  elp & elq & ELR  |  ELP & ELQ & ELR  ;
 flc <=  ELP & elq & elr  |  elp & ELQ & elr  |  elp & elq & ELR  |  elp & elq & elr  ;
 FKD <=  ELM & eln & elo  |  elm & ELN & elo  |  elm & eln & ELO  |  ELM & ELN & ELO  ;
 fld <=  ELM & eln & elo  |  elm & ELN & elo  |  elm & eln & ELO  |  elm & eln & elo  ;
 FKE <=  ELJ & elk & ell  |  elj & ELK & ell  |  elj & elk & ELL  |  ELJ & ELK & ELL  ;
 fle <=  ELJ & elk & ell  |  elj & ELK & ell  |  elj & elk & ELL  |  elj & elk & ell  ;
 FKF <=  ELG & elh & eli  |  elg & ELH & eli  |  elg & elh & ELI  |  ELG & ELH & ELI  ;
 flf <=  ELG & elh & eli  |  elg & ELH & eli  |  elg & elh & ELI  |  elg & elh & eli  ;
 AAM <=  ICM & TSA  |  BAM & TKA  |  AAM & THA  ; 
 AAN <=  ICN & TSA  |  BAN & TKA  |  AAN & THA  ; 
 FKA <=  ELX & elw & elv  |  elx & ELW & elv  |  elx & elw & ELV  |  ELX & ELW & ELV  ;
 fla <=  ELX & elw & elv  |  elx & ELW & elv  |  elx & elw & ELV  |  elx & elw & elv  ;
 FKB <=  ELS & elt & elu  |  els & ELT & elu  |  els & elt & ELU  |  ELS & ELT & ELU  ;
 flb <=  ELS & elt & elu  |  els & ELT & elu  |  els & elt & ELU  |  els & elt & elu  ;
 oca <= ida ; 
 ocb <= idb ; 
 occ <= idc ; 
 ocd <= idd ; 
 oce <= ide ; 
 ocf <= idf ; 
 ocg <= idg ; 
 och <= idh ; 
 oci <= idi ; 
 ocj <= idj ; 
 ock <= idk ; 
 ocl <= idl ; 
 ocm <= idm ; 
 ocn <= idn ; 
 oco <= ido ; 
 ocp <= idp ; 
 AAH <=  ICH & TSB  |  BAH & TKB  |  AAH & THB  ; 
 AAI <=  ICI & TSA  |  BAI & TKA  |  AAI & THA  ; 
 AAJ <=  ICJ & TSA  |  BAJ & TKA  |  AAJ & THA  ; 
 AAK <=  ICK & TSB  |  BAK & TKB  |  AAK & THB  ; 
 FGL <=  EGM & egn & ego  |  egm & EGN & ego  |  egm & egn & EGO  |  EGM & EGN & EGO  ;
 fhl <=  EGM & egn & ego  |  egm & EGN & ego  |  egm & egn & EGO  |  egm & egn & ego  ;
 FGP <= EGF ; 
 FGM <=  EGL & egk & egj  |  egl & EGK & egj  |  egl & egk & EGJ  |  EGL & EGK & EGJ  ;
 fhm <=  EGL & egk & egj  |  egl & EGK & egj  |  egl & egk & EGJ  |  egl & egk & egj  ;
 FGO <= QIC ; 
 FGN <=  EGI & egh & egg  |  egi & EGH & egg  |  egi & egh & EGG  |  EGI & EGH & EGG  ;
 fhn <=  EGI & egh & egg  |  egi & EGH & egg  |  egi & egh & EGG  |  egi & egh & egg  ;
 FGI <=  EGX & egw & egv  |  egx & EGW & egv  |  egx & egw & EGV  |  EGX & EGW & EGV  ;
 fhi <=  EGX & egw & egv  |  egx & EGW & egv  |  egx & egw & EGV  |  egx & egw & egv  ;
 FGJ <=  EGS & egt & egu  |  egs & EGT & egu  |  egs & egt & EGU  |  EGS & EGT & EGU  ;
 fhj <=  EGS & egt & egu  |  egs & EGT & egu  |  egs & egt & EGU  |  egs & egt & egu  ;
 FGK <=  EGP & egq & egr  |  egp & EGQ & egr  |  egp & egq & EGR  |  EGP & EGQ & EGR  ;
 fhk <=  EGP & egq & egr  |  egp & EGQ & egr  |  egp & egq & EGR  |  egp & egq & egr  ;
 FGF <=  EHG & ehh & ehi  |  ehg & EHH & ehi  |  ehg & ehh & EHI  |  EHG & EHH & EHI  ;
 fhf <=  EHG & ehh & ehi  |  ehg & EHH & ehi  |  ehg & ehh & EHI  |  ehg & ehh & ehi  ;
 FGG <=  EHD & ehe & ehf  |  ehd & EHE & ehf  |  ehd & ehe & EHF  |  EHD & EHE & EHF  ;
 fhg <=  EHD & ehe & ehf  |  ehd & EHE & ehf  |  ehd & ehe & EHF  |  ehd & ehe & ehf  ;
 FGH <=  EHA & ehb & ehc  |  eha & EHB & ehc  |  eha & ehb & EHC  |  EHA & EHB & EHC  ;
 fhh <=  EHA & ehb & ehc  |  eha & EHB & ehc  |  eha & ehb & EHC  |  eha & ehb & ehc  ;
 FIL <=  EIM & ein & eio  |  eim & EIN & eio  |  eim & ein & EIO  |  EIM & EIN & EIO  ;
 fjl <=  EIM & ein & eio  |  eim & EIN & eio  |  eim & ein & EIO  |  eim & ein & eio  ;
 FIM <=  EIL & eik & eij  |  eil & EIK & eij  |  eil & eik & EIJ  |  EIL & EIK & EIJ  ;
 fjm <=  EIL & eik & eij  |  eil & EIK & eij  |  eil & eik & EIJ  |  eil & eik & eij  ;
 FIN <=  EII & eih & qid  |  eii & EIH & qid  |  eii & eih & QID  |  EII & EIH & QID  ;
 fjn <=  EII & eih & qid  |  eii & EIH & qid  |  eii & eih & QID  |  eii & eih & qid  ;
 FIO <= EIG ; 
 FII <=  EIX & eiw & eiv  |  eix & EIW & eiv  |  eix & eiw & EIV  |  EIX & EIW & EIV  ;
 fji <=  EIX & eiw & eiv  |  eix & EIW & eiv  |  eix & eiw & EIV  |  eix & eiw & eiv  ;
 FIJ <=  EIS & eit & eiu  |  eis & EIT & eiu  |  eis & eit & EIU  |  EIS & EIT & EIU  ;
 fjj <=  EIS & eit & eiu  |  eis & EIT & eiu  |  eis & eit & EIU  |  eis & eit & eiu  ;
 FIK <=  EIP & eiq & eir  |  eip & EIQ & eir  |  eip & eiq & EIR  |  EIP & EIQ & EIR  ;
 fjk <=  EIP & eiq & eir  |  eip & EIQ & eir  |  eip & eiq & EIR  |  eip & eiq & eir  ;
 FIF <=  EJG & ejh & eji  |  ejg & EJH & eji  |  ejg & ejh & EJI  |  EJG & EJH & EJI  ;
 fjf <=  EJG & ejh & eji  |  ejg & EJH & eji  |  ejg & ejh & EJI  |  ejg & ejh & eji  ;
 FIG <=  EJD & eje & ejf  |  ejd & EJE & ejf  |  ejd & eje & EJF  |  EJD & EJE & EJF  ;
 fjg <=  EJD & eje & ejf  |  ejd & EJE & ejf  |  ejd & eje & EJF  |  ejd & eje & ejf  ;
 FIH <=  EJA & ejb & ejc  |  eja & EJB & ejc  |  eja & ejb & EJC  |  EJA & EJB & EJC  ;
 fjh <=  EJA & ejb & ejc  |  eja & EJB & ejc  |  eja & ejb & EJC  |  eja & ejb & ejc  ;
 FKL <=  EKM & ekn & eko  |  ekm & EKN & eko  |  ekm & ekn & EKO  |  EKM & EKN & EKO  ;
 fll <=  EKM & ekn & eko  |  ekm & EKN & eko  |  ekm & ekn & EKO  |  ekm & ekn & eko  ;
 QIE <= QIA ; 
 FKM <=  EKL & ekk & ekj  |  ekl & EKK & ekj  |  ekl & ekk & EKJ  |  EKL & EKK & EKJ  ;
 flm <=  EKL & ekk & ekj  |  ekl & EKK & ekj  |  ekl & ekk & EKJ  |  ekl & ekk & ekj  ;
 FKN <=  EKI & ekh & qid  |  eki & EKH & qid  |  eki & ekh & QID  |  EKI & EKH & QID  ;
 fln <=  EKI & ekh & qid  |  eki & EKH & qid  |  eki & ekh & QID  |  eki & ekh & qid  ;
 FKI <=  EKX & ekw & ekv  |  ekx & EKW & ekv  |  ekx & ekw & EKV  |  EKX & EKW & EKV  ;
 fli <=  EKX & ekw & ekv  |  ekx & EKW & ekv  |  ekx & ekw & EKV  |  ekx & ekw & ekv  ;
 QIA <= ITB ; 
 QIB <= QIA ; 
 QIC <= QIA ; 
 QID <= QIA ; 
 FKJ <=  EKS & ekt & eku  |  eks & EKT & eku  |  eks & ekt & EKU  |  EKS & EKT & EKU  ;
 flj <=  EKS & ekt & eku  |  eks & EKT & eku  |  eks & ekt & EKU  |  eks & ekt & eku  ;
 FKK <=  EKP & ekq & ekr  |  ekp & EKQ & ekr  |  ekp & ekq & EKR  |  EKP & EKQ & EKR  ;
 flk <=  EKP & ekq & ekr  |  ekp & EKQ & ekr  |  ekp & ekq & EKR  |  ekp & ekq & ekr  ;
 CAI <= AAI ; 
 CDI <= AAI ; 
 CAJ <= AAJ ; 
 CDJ <= AAJ ; 
 CAK <= AAK ; 
 CDK <= AAK ; 
 CAL <= AAL ; 
 CDL <= AAL ; 
 CAM <= AAM ; 
 CDM <= AAM ; 
 CAN <= AAN ; 
 CDN <= AAN ; 
 DBA <= IFA ; 
 dea <= ifa ; 
 DBB <= IFB ; 
 deb <= ifb ; 
 DBC <= IFC ; 
 dec <= ifc ; 
 DBD <= IFD ; 
 ded <= ifd ; 
 DGI <= BAI ; 
 DGJ <= BAJ ; 
 DGK <= BAK ; 
 DGL <= BAL ; 
 DBE <= IFE ; 
 dee <= ife ; 
 DBF <= IFFF  ; 
 def <= ifff  ; 
 DGE <= BAE ; 
 DGF <= BAF ; 
 DGG <= BAG ; 
 DGH <= BAH ; 
 DBG <= IFG ; 
 deg <= ifg ; 
 DBH <= IFH ; 
 deh <= ifh ; 
 FQL <=  EQM & eqn & eqo  |  eqm & EQN & eqo  |  eqm & eqn & EQO  |  EQM & EQN & EQO  ;
 ogl <=  EQM & eqn & eqo  |  eqm & EQN & eqo  |  eqm & eqn & EQO  |  eqm & eqn & eqo  ;
 FQM <=  EQL & eqk & qie  |  eql & EQK & qie  |  eql & eqk & QIE  |  EQL & EQK & QIE  ;
 ogm <=  EQL & eqk & qie  |  eql & EQK & qie  |  eql & eqk & QIE  |  eql & eqk & qie  ;
 FOA <=  EPX & epw & epv  |  epx & EPW & epv  |  epx & epw & EPV  |  EPX & EPW & EPV  ;
 fpa <=  EPX & epw & epv  |  epx & EPW & epv  |  epx & epw & EPV  |  epx & epw & epv  ;
 FOB <=  EPS & ept & epu  |  eps & EPT & epu  |  eps & ept & EPU  |  EPS & EPT & EPU  ;
 fpb <=  EPS & ept & epu  |  eps & EPT & epu  |  eps & ept & EPU  |  eps & ept & epu  ;
 FQH <=  ERA & erb & erc  |  era & ERB & erc  |  era & erb & ERC  |  ERA & ERB & ERC  ;
 ogh <=  ERA & erb & erc  |  era & ERB & erc  |  era & erb & ERC  |  era & erb & erc  ;
 FQI <=  EQX & eqw & eqv  |  eqx & EQW & eqv  |  eqx & eqw & EQV  |  EQX & EQW & EQV  ;
 ogi <=  EQX & eqw & eqv  |  eqx & EQW & eqv  |  eqx & eqw & EQV  |  eqx & eqw & eqv  ;
 FQJ <=  EQS & eqt & equ  |  eqs & EQT & equ  |  eqs & eqt & EQU  |  EQS & EQT & EQU  ;
 ogj <=  EQS & eqt & equ  |  eqs & EQT & equ  |  eqs & eqt & EQU  |  eqs & eqt & equ  ;
 FQK <=  EQP & eqq & eqr  |  eqp & EQQ & eqr  |  eqp & eqq & EQR  |  EQP & EQQ & EQR  ;
 ogk <=  EQP & eqq & eqr  |  eqp & EQQ & eqr  |  eqp & eqq & EQR  |  eqp & eqq & eqr  ;
 FQD <=  ERM & ern & ero  |  erm & ERN & ero  |  erm & ern & ERO  |  ERM & ERN & ERO  ;
 ogd <=  ERM & ern & ero  |  erm & ERN & ero  |  erm & ern & ERO  |  erm & ern & ero  ;
 FQE <=  ERJ & erk & erl  |  erj & ERK & erl  |  erj & erk & ERL  |  ERJ & ERK & ERL  ;
 oge <=  ERJ & erk & erl  |  erj & ERK & erl  |  erj & erk & ERL  |  erj & erk & erl  ;
 FQF <=  ERG & erh & eri  |  erg & ERH & eri  |  erg & erh & ERI  |  ERG & ERH & ERI  ;
 ogf <=  ERG & erh & eri  |  erg & ERH & eri  |  erg & erh & ERI  |  erg & erh & eri  ;
 FQG <=  ERD & ere & erf  |  erd & ERE & erf  |  erd & ere & ERF  |  ERD & ERE & ERF  ;
 ogg <=  ERD & ere & erf  |  erd & ERE & erf  |  erd & ere & ERF  |  erd & ere & erf  ;
 FQA <=  ERX & erw & erv  |  erx & ERW & erv  |  erx & erw & ERV  |  ERX & ERW & ERV  ;
 oga <=  ERX & erw & erv  |  erx & ERW & erv  |  erx & erw & ERV  |  erx & erw & erv  ;
 BAC <=  IDC & TTB  |  BEC & TGB  ; 
 FQB <=  ERS & ert & eru  |  ers & ERT & eru  |  ers & ert & ERU  |  ERS & ERT & ERU  ;
 ogb <=  ERS & ert & eru  |  ers & ERT & eru  |  ers & ert & ERU  |  ers & ert & eru  ;
 FQC <=  ERP & erq & err  |  erp & ERQ & err  |  erp & erq & ERR  |  ERP & ERQ & ERR  ;
 ogc <=  ERP & erq & err  |  erp & ERQ & err  |  erp & erq & ERR  |  erp & erq & err  ;
 BAD <=  IDD & TTB  |  BED & TGB  ; 
 BAE <=  IDE & TTA  |  BEE & TGA  ; 
 BAF <=  IDF & TTA  |  BEF & TGA  ; 
 BAG <=  IDG & TTB  |  BEG & TGB  ; 
 BAH <=  IDH & TTB  |  BEH & TGB  ; 
 BAI <=  IDI & TTA  |  BEI & TGA  ; 
 BAJ <=  IDJ & TTA  |  BEJ & TGA  ; 
 BAK <=  IDK & TTB  |  BEK & TGB  ; 
 AAO <=  ICO & TSB  |  BAO & TKB  |  AAO & THB  ; 
 AAP <=  ICP & TSB  |  BAP & TKB  |  AAP & THB  ; 
 BAA <=  IDA & TTA  |  BEA & TGA  ; 
 BAB <=  IDB & TTA  |  BEB & TGA  ; 
 FMK <=  EMP & emq & emr  |  emp & EMQ & emr  |  emp & emq & EMR  |  EMP & EMQ & EMR  ;
 fnk <=  EMP & emq & emr  |  emp & EMQ & emr  |  emp & emq & EMR  |  emp & emq & emr  ;
 FML <=  EMM & emn & emo  |  emm & EMN & emo  |  emm & emn & EMO  |  EMM & EMN & EMO  ;
 fnl <=  EMM & emn & emo  |  emm & EMN & emo  |  emm & emn & EMO  |  emm & emn & emo  ;
 FMO <= QIE ; 
 FMM <=  EML & emk & emj  |  eml & EMK & emj  |  eml & emk & EMJ  |  EML & EMK & EMJ  ;
 fnm <=  EML & emk & emj  |  eml & EMK & emj  |  eml & emk & EMJ  |  eml & emk & emj  ;
 FMN <= EMI ; 
 FMH <=  ENA & enb & enc  |  ena & ENB & enc  |  ena & enb & ENC  |  ENA & ENB & ENC  ;
 fnh <=  ENA & enb & enc  |  ena & ENB & enc  |  ena & enb & ENC  |  ena & enb & enc  ;
 FMI <=  EMX & emw & emv  |  emx & EMW & emv  |  emx & emw & EMV  |  EMX & EMW & EMV  ;
 fni <=  EMX & emw & emv  |  emx & EMW & emv  |  emx & emw & EMV  |  emx & emw & emv  ;
 FMJ <=  EMS & emt & emu  |  ems & EMT & emu  |  ems & emt & EMU  |  EMS & EMT & EMU  ;
 fnj <=  EMS & emt & emu  |  ems & EMT & emu  |  ems & emt & EMU  |  ems & emt & emu  ;
 FME <=  ENJ & enk & enl  |  enj & ENK & enl  |  enj & enk & ENL  |  ENJ & ENK & ENL  ;
 fne <=  ENJ & enk & enl  |  enj & ENK & enl  |  enj & enk & ENL  |  enj & enk & enl  ;
 FMF <=  ENG & enh & eni  |  eng & ENH & eni  |  eng & enh & ENI  |  ENG & ENH & ENI  ;
 fnf <=  ENG & enh & eni  |  eng & ENH & eni  |  eng & enh & ENI  |  eng & enh & eni  ;
 FMG <=  ENDD  & ene & enf  |  endd & ENE & enf  |  endd & ene & ENF  |  ENDD  & ENE & ENF  ;
 fng <=  ENDD  & ene & enf  |  endd & ENE & enf  |  endd & ene & ENF  |  endd & ene & enf  ;
 FMB <=  ENS & ent & enu  |  ens & ENT & enu  |  ens & ent & ENU  |  ENS & ENT & ENU  ;
 fnb <=  ENS & ent & enu  |  ens & ENT & enu  |  ens & ent & ENU  |  ens & ent & enu  ;
 FMC <=  ENP & enq & enr  |  enp & ENQ & enr  |  enp & enq & ENR  |  ENP & ENQ & ENR  ;
 fnc <=  ENP & enq & enr  |  enp & ENQ & enr  |  enp & enq & ENR  |  enp & enq & enr  ;
 FMD <=  ENM & enn & eno  |  enm & ENN & eno  |  enm & enn & ENO  |  ENM & ENN & ENO  ;
 fnd <=  ENM & enn & eno  |  enm & ENN & eno  |  enm & enn & ENO  |  enm & enn & eno  ;
 FOL <=  EOM & eon & eoo  |  eom & EON & eoo  |  eom & eon & EOO  |  EOM & EON & EOO  ;
 fpl <=  EOM & eon & eoo  |  eom & EON & eoo  |  eom & eon & EOO  |  eom & eon & eoo  ;
 FOM <=  QIE & eok & eol  |  qie & EOK & eol  |  qie & eok & EOL  |  QIE & EOK & EOL  ;
 fpm <=  QIE & eok & eol  |  qie & EOK & eol  |  qie & eok & EOL  |  qie & eok & eol  ;
 FON <= EOJ ; 
 FMA <=  ENX & enw & env  |  enx & ENW & env  |  enx & enw & ENV  |  ENX & ENW & ENV  ;
 fna <=  ENX & enw & env  |  enx & ENW & env  |  enx & enw & ENV  |  enx & enw & env  ;
 FOI <=  EOX & eow & eov  |  eox & EOW & eov  |  eox & eow & EOV  |  EOX & EOW & EOV  ;
 fpi <=  EOX & eow & eov  |  eox & EOW & eov  |  eox & eow & EOV  |  eox & eow & eov  ;
 FOJ <=  EOS & eot & eou  |  eos & EOT & eou  |  eos & eot & EOU  |  EOS & EOT & EOU  ;
 fpj <=  EOS & eot & eou  |  eos & EOT & eou  |  eos & eot & EOU  |  eos & eot & eou  ;
 FOK <=  EOP & eoq & eor  |  eop & EOQ & eor  |  eop & eoq & EOR  |  EOP & EOQ & EOR  ;
 fpk <=  EOP & eoq & eor  |  eop & EOQ & eor  |  eop & eoq & EOR  |  eop & eoq & eor  ;
 FOF <=  EPG & eph & epi  |  epg & EPH & epi  |  epg & eph & EPI  |  EPG & EPH & EPI  ;
 fpf <=  EPG & eph & epi  |  epg & EPH & epi  |  epg & eph & EPI  |  epg & eph & epi  ;
 FOG <=  EPD & epe & epf  |  epd & EPE & epf  |  epd & epe & EPF  |  EPD & EPE & EPF  ;
 fpg <=  EPD & epe & epf  |  epd & EPE & epf  |  epd & epe & EPF  |  epd & epe & epf  ;
 FOH <=  EPA & epb & epc  |  epa & EPB & epc  |  epa & epb & EPC  |  EPA & EPB & EPC  ;
 fph <=  EPA & epb & epc  |  epa & EPB & epc  |  epa & epb & EPC  |  epa & epb & epc  ;
 FOC <=  EPP & epq & epr  |  epp & EPQ & epr  |  epp & epq & EPR  |  EPP & EPQ & EPR  ;
 fpc <=  EPP & epq & epr  |  epp & EPQ & epr  |  epp & epq & EPR  |  epp & epq & epr  ;
 FOD <=  EPM & epn & epo  |  epm & EPN & epo  |  epm & epn & EPO  |  EPM & EPN & EPO  ;
 fpd <=  EPM & epn & epo  |  epm & EPN & epo  |  epm & epn & EPO  |  epm & epn & epo  ;
 FOE <=  EPJ & epk & epl  |  epj & EPK & epl  |  epj & epk & EPL  |  EPJ & EPK & EPL  ;
 fpe <=  EPJ & epk & epl  |  epj & EPK & epl  |  epj & epk & EPL  |  epj & epk & epl  ;
 BAP <=  IDP & TTB  |  BEP & TGB  ; 
 CAO <= AAO ; 
 CDO <= AAO ; 
 CAF <= AAF ; 
 CDF <= AAF ; 
 CAP <= AAP ; 
 CDP <= AAP ; 
 CBA <= IBA ; 
 CEA <= IBA ; 
 CBB <= IBB ; 
 CEB <= IBB ; 
 CBC <= IBC ; 
 CEC <= IBC ; 
 CBD <= IBD ; 
 CED <= IBD ; 
 DBI <= IFI ; 
 dei <= ifi ; 
 DBJ <= IFJ ; 
 dej <= ifj ; 
 DGM <= BAM ; 
 DGN <= BAN ; 
 DGO <= BAO ; 
 DGP <= BAP ; 
 DBK <= IFK ; 
 dek <= ifk ; 
 DBL <= IFL ; 
 del <= ifl ; 
 BAL <=  IDL & TTB  |  BEL & TGB  ; 
 DBM <= IFM ; 
 dem <= ifm ; 
 DBN <= IFN ; 
 den <= ifn ; 
 BAM <=  IDM & TTA  |  BEM & TGA  ; 
 BAN <=  IDN & TTA  |  BEN & TGA  ; 
 BAO <=  IDO & TTB  |  BEO & TGB  ; 
 DBO <= IFO ; 
 deo <= ifo ; 
 DBP <= IFP ; 
 dep <= ifp ; 
 bba <= ida ; 
 bbb <= idb ; 
 bbc <= idc ; 
 bbd <= idd ; 
 bbe <= ide ; 
 bbf <= idf ; 
 bbg <= idg ; 
 bbh <= idh ; 
 bbi <= idi ; 
 bbj <= idj ; 
 bbk <= idk ; 
 bbl <= idl ; 
 bbm <= idm ; 
 bbn <= idn ; 
 bbo <= ido ; 
 bbp <= idp ; 
 BCA <= BBA ; 
 BCB <= BBB ; 
 BCC <= BBC ; 
 BCD <= BBD ; 
 BCE <= BBE ; 
 BCF <= BBF ; 
 BCG <= BBG ; 
 BCH <= BBH ; 
 BCI <= BBI ; 
 BCJ <= BBJ ; 
 BCK <= BBK ; 
 BCL <= BBL ; 
 BCM <= BBM ; 
 BCN <= BBN ; 
 BCO <= BBO ; 
 BCP <= BBP ; 
 QTA <= ITA ; 
 TTA <= QTA ; 
 TTB <= QTA ; 
 TTC <= QTA ; 
 OPI <=  NIA & nha & mic  |  nia & NHA & mic  |  nia & nha & MIC  |  NIA & NHA & MIC  ;
 oqi <=  NIA & nha & mic  |  nia & NHA & mic  |  nia & nha & MIC  |  nia & nha & mic  ;
 CBE <= IBE ; 
 CEE <= IBE ; 
 CBF <= IBF ; 
 CEF <= IBF ; 
 BDM <= BCM ; 
 BDN <= BCN ; 
 BDO <= BCO ; 
 BDP <= BCP ; 
 CBG <= IEA & TRB |  IBG & trb ; 
 CBH <= IEB & TRB |  IBH & trb ; 
 CBI <= IEC & TRB |  IBI & trb ; 
 OPO <=  NNA & mna & noa  |  nna & MNA & noa  |  nna & mna & NOA  |  NNA & MNA & NOA  ;
 oqo <=  NNA & mna & noa  |  nna & MNA & noa  |  nna & mna & NOA  |  nna & mna & noa  ;
 CEG <= IEA & TRA |  IBG & tra ; 
 CEH <= IEB & TRA |  IBH & tra ; 
 CEI <= IEC & TRA |  IBI & tra ; 
 OPQ <=  NQA & npa & mpa  |  nqa & NPA & mpa  |  nqa & npa & MPA  |  NQA & NPA & MPA  ;
 oqq <=  NQA & npa & mpa  |  nqa & NPA & mpa  |  nqa & npa & MPA  |  nqa & npa & mpa  ;
 OPR <= NRA ; 
 QKA <= IKA ; 
 TKA <= QKA ; 
 TKB <= QKA ; 
 TKC <= QKA ; 
 DCA <= IGA ; 
 dfa <= iga ; 
 DCB <= IGB ; 
 dfb <= igb ; 
 TKD <= QKA ; 
 TKE <= QKA ; 
 TKF <= QKA ; 
 DCC <= IGC ; 
 dfc <= igc ; 
 DCD <= IGD ; 
 dfd <= igd ; 
 OPK <=  NJA & nka & mja  |  nja & NKA & mja  |  nja & nka & MJA  |  NJA & NKA & MJA  ;
 oqk <=  NJA & nka & mja  |  nja & NKA & mja  |  nja & nka & MJA  |  nja & nka & mja  ;
 DCE <= IGE ; 
 dfe <= ige ; 
 DCF <= IGF ; 
 dff <= igf ; 
 BDA <= BCA ; 
 BDB <= BCB ; 
 BDC <= BCC ; 
 BDD <= BCD ; 
 BDE <= BCE ; 
 BDF <= BCF ; 
 BDG <= BCG ; 
 BDH <= BCH ; 
 BDI <= BCI ; 
 BDJ <= BCJ ; 
 BDK <= BCK ; 
 BDL <= BCL ; 
 DCG <= IGG ; 
 dfg <= igg ; 
 DCH <= IGH ; 
 dfh <= igh ; 
 BEM <= BDM ; 
 BEN <= BDN ; 
 BEO <= BDO ; 
 BEP <= BDP ; 
 BEA <= BDA ; 
 BEB <= BDB ; 
 BEC <= BDC ; 
 BED <= BDD ; 
 BEE <= BDE ; 
 BEF <= BDF ; 
 BEG <= BDG ; 
 BEH <= BDH ; 
 BEI <= BDI ; 
 BEJ <= BDJ ; 
 BEK <= BDK ; 
 BEL <= BDL ; 
 CBJ <= IED & TRB |  IBJ & trb ; 
 CBK <= IEE & TRB |  IBK & trb ; 
 CBL <= IEF & TRB |  IBL & trb ; 
 CEJ <= IED & TRA |  IBJ & tra ; 
 CEK <= IEE & TRA |  IBK & tra ; 
 CEL <= IEF & TRA |  IBL & tra ; 
 OPE <=  MEA & mda & nda  |  mea & MDA & nda  |  mea & mda & NDA  |  MEA & MDA & NDA  ;
 oqe <=  MEA & mda & nda  |  mea & MDA & nda  |  mea & mda & NDA  |  mea & mda & nda  ;
 OPF <= NEA ; 
 OPG <= NFA ; 
 OPH <= NGA ; 
 CBM <= IEG & TRB |  IBM & trb ; 
 CBN <= IEH & TRB |  IBN & trb ; 
 CBO <= IEI & TRB |  IBO & trb ; 
 OPM <=  MMC & nla & nma  |  mmc & NLA & nma  |  mmc & nla & NMA  |  MMC & NLA & NMA  ;
 oqm <=  MMC & nla & nma  |  mmc & NLA & nma  |  mmc & nla & NMA  |  mmc & nla & nma  ;
 CEM <= IEG & TRA |  IBM & tra ; 
 CEN <= IEH & TRA |  IBN & tra ; 
 CEO <= IEI & TRA |  IBO & tra ; 
 OPA <=  NAA & mab & ioa  |  naa & MAB & ioa  |  naa & mab & IOA  |  NAA & MAB & IOA  ;
 oqa <=  NAA & mab & ioa  |  naa & MAB & ioa  |  naa & mab & IOA  |  naa & mab & ioa  ;
 OPB <= IOB ; 
 CBP <= IEJ & TRB |  IBP & trb ; 
 CEP <= IEJ & TRB |  IBP & trb ; 
 OPC <=  NCA & nba & mbb  |  nca & NBA & mbb  |  nca & nba & MBB  |  NCA & NBA & MBB  ;
 oqc <=  NCA & nba & mbb  |  nca & NBA & mbb  |  nca & nba & MBB  |  nca & nba & mbb  ;
 OPD <= IOC ; 
 QGA <= IIA ; 
 TGA <= QGA ; 
 TGB <= QGA ; 
 TGC <= QGA ; 
 DCI <= IGI ; 
 dfi <= igi ; 
 DCJ <= IGJ ; 
 dfj <= igj ; 
 DCK <= IGK ; 
 dfk <= igk ; 
 DCL <= IGL ; 
 dfl <= igl ; 
 DCM <= IGM ; 
 dfm <= igm ; 
 DCN <= IGN ; 
 dfn <= ign ; 
 DCO <= IGO ; 
 dfo <= igo ; 
 DCP <= IGP ; 
 dfp <= igp ; 
 HIB <=  GHA & gia & ghd  |  gha & GIA & ghd  |  gha & gia & GHD  |  GHA & GIA & GHD  ;
 hjb <=  GHA & gia & ghd  |  gha & GIA & ghd  |  gha & gia & GHD  |  gha & gia & ghd  ;
 HGG <=  GGI & gfi & fgo  |  ggi & GFI & fgo  |  ggi & gfi & FGO  |  GGI & GFI & FGO  ;
 hhg <=  GGI & gfi & fgo  |  ggi & GFI & fgo  |  ggi & gfi & FGO  |  ggi & gfi & fgo  ;
 HGD <=  GGE & gfe & ggd  |  gge & GFE & ggd  |  gge & gfe & GGD  |  GGE & GFE & GGD  ;
 hhd <=  GGE & gfe & ggd  |  gge & GFE & ggd  |  gge & gfe & GGD  |  gge & gfe & ggd  ;
 HQF <=  GPH & gqh & gpi  |  gph & GQH & gpi  |  gph & gqh & GPI  |  GPH & GQH & GPI  ;
 ohf <=  GPH & gqh & gpi  |  gph & GQH & gpi  |  gph & gqh & GPI  |  gph & gqh & gpi  ;
 HQG <= FQJ ; 
 HIE <=  GHH & gih & gig  |  ghh & GIH & gig  |  ghh & gih & GIG  |  GHH & GIH & GIG  ;
 hje <=  GHH & gih & gig  |  ghh & GIH & gig  |  ghh & gih & GIG  |  ghh & gih & gig  ;
 HIF <=  GHG & fhg & ghj  |  ghg & FHG & ghj  |  ghg & fhg & GHJ  |  GHG & FHG & GHJ  ;
 hjf <=  GHG & fhg & ghj  |  ghg & FHG & ghj  |  ghg & fhg & GHJ  |  ghg & fhg & ghj  ;
 HIC <=  GHF & gif & gic  |  ghf & GIF & gic  |  ghf & gif & GIC  |  GHF & GIF & GIC  ;
 hjc <=  GHF & gif & gic  |  ghf & GIF & gic  |  ghf & gif & GIC  |  ghf & gif & gic  ;
 HIA <=  GHB & gib & ghc  |  ghb & GIB & ghc  |  ghb & gib & GHC  |  GHB & GIB & GHC  ;
 hja <=  GHB & gib & ghc  |  ghb & GIB & ghc  |  ghb & gib & GHC  |  ghb & gib & ghc  ;
 HKA <=  GJB & gkb & gjc  |  gjb & GKB & gjc  |  gjb & gkb & GJC  |  GJB & GKB & GJC  ;
 hla <=  GJB & gkb & gjc  |  gjb & GKB & gjc  |  gjb & gkb & GJC  |  gjb & gkb & gjc  ;
 HKB <=  GJA & gka & gjd  |  gja & GKA & gjd  |  gja & gka & GJD  |  GJA & GKA & GJD  ;
 hlb <=  GJA & gka & gjd  |  gja & GKA & gjd  |  gja & gka & GJD  |  gja & gka & gjd  ;
 HIG <=  GII & ghi & fhk  |  gii & GHI & fhk  |  gii & ghi & FHK  |  GII & GHI & FHK  ;
 hjg <=  GII & ghi & fhk  |  gii & GHI & fhk  |  gii & ghi & FHK  |  gii & ghi & fhk  ;
 HID <=  GID & ghe & gie  |  gid & GHE & gie  |  gid & ghe & GIE  |  GID & GHE & GIE  ;
 hjd <=  GID & ghe & gie  |  gid & GHE & gie  |  gid & ghe & GIE  |  gid & ghe & gie  ;
 HKE <=  GJH & gkh & gjg  |  gjh & GKH & gjg  |  gjh & gkh & GJG  |  GJH & GKH & GJG  ;
 hle <=  GJH & gkh & gjg  |  gjh & GKH & gjg  |  gjh & gkh & GJG  |  gjh & gkh & gjg  ;
 HKC <=  GJF & gkf & gkc  |  gjf & GKF & gkc  |  gjf & gkf & GKC  |  GJF & GKF & GKC  ;
 hlc <=  GJF & gkf & gkc  |  gjf & GKF & gkc  |  gjf & gkf & GKC  |  gjf & gkf & gkc  ;
 HKF <=  GKI & gji & gkg  |  gki & GJI & gkg  |  gki & gji & GKG  |  GKI & GJI & GKG  ;
 hlf <=  GKI & gji & gkg  |  gki & GJI & gkg  |  gki & gji & GKG  |  gki & gji & gkg  ;
 HKG <= FJG ; 
 HKD <=  GKD & gje & gke  |  gkd & GJE & gke  |  gkd & gje & GKE  |  GKD & GJE & GKE  ;
 hld <=  GKD & gje & gke  |  gkd & GJE & gke  |  gkd & gje & GKE  |  gkd & gje & gke  ;
 HMC <=  GLF & gme & fmo  |  glf & GME & fmo  |  glf & gme & FMO  |  GLF & GME & FMO  ;
 hnc <=  GLF & gme & fmo  |  glf & GME & fmo  |  glf & gme & FMO  |  glf & gme & fmo  ;
 HMD <=  GLD & gmc & gle  |  gld & GMC & gle  |  gld & gmc & GLE  |  GLD & GMC & GLE  ;
 hnd <=  GLD & gmc & gle  |  gld & GMC & gle  |  gld & gmc & GLE  |  gld & gmc & gle  ;
 HMA <=  GLC & glb & gmb  |  glc & GLB & gmb  |  glc & glb & GMB  |  GLC & GLB & GMB  ;
 hna <=  GLC & glb & gmb  |  glc & GLB & gmb  |  glc & glb & GMB  |  glc & glb & gmb  ;
 HMB <=  GLA & gma & gmd  |  gla & GMA & gmd  |  gla & gma & GMD  |  GLA & GMA & GMD  ;
 hnb <=  GLA & gma & gmd  |  gla & GMA & gmd  |  gla & gma & GMD  |  gla & gma & gmd  ;
 HOD <=  GNF & gnh & gng  |  gnf & GNH & gng  |  gnf & gnh & GNG  |  GNF & GNH & GNG  ;
 hpd <=  GNF & gnh & gng  |  gnf & GNH & gng  |  gnf & gnh & GNG  |  gnf & gnh & gng  ;
 HOB <=  GNC & gne & gnb  |  gnc & GNE & gnb  |  gnc & gne & GNB  |  GNC & GNE & GNB  ;
 hpb <=  GNC & gne & gnb  |  gnc & GNE & gnb  |  gnc & gne & GNB  |  gnc & gne & gnb  ;
 HME <=  GMH & gli & glh  |  gmh & GLI & glh  |  gmh & gli & GLH  |  GMH & GLI & GLH  ;
 hne <=  GMH & gli & glh  |  gmh & GLI & glh  |  gmh & gli & GLH  |  gmh & gli & glh  ;
 HMH <= GMF ; 
 HMF <=  GLG & gmg & gmi  |  glg & GMG & gmi  |  glg & gmg & GMI  |  GLG & GMG & GMI  ;
 hnf <=  GLG & gmg & gmi  |  glg & GMG & gmi  |  glg & gmg & GMI  |  glg & gmg & gmi  ;
 HMG <= FMM ; 
 HOE <=  GOF & goe & gog  |  gof & GOE & gog  |  gof & goe & GOG  |  GOF & GOE & GOG  ;
 hpe <=  GOF & goe & gog  |  gof & GOE & gog  |  gof & goe & GOG  |  gof & goe & gog  ;
 HOC <=  GOC & gnd & god  |  goc & GND & god  |  goc & gnd & GOD  |  GOC & GND & GOD  ;
 hpc <=  GOC & gnd & god  |  goc & GND & god  |  goc & gnd & GOD  |  goc & gnd & god  ;
 HOA <=  GOA & gob & gna  |  goa & GOB & gna  |  goa & gob & GNA  |  GOA & GOB & GNA  ;
 hpa <=  GOA & gob & gna  |  goa & GOB & gna  |  goa & gob & GNA  |  goa & gob & gna  ;
 HOF <=  GNI & goi & goh  |  gni & GOI & goh  |  gni & goi & GOH  |  GNI & GOI & GOH  ;
 hpf <=  GNI & goi & goh  |  gni & GOI & goh  |  gni & goi & GOH  |  gni & goi & goh  ;
 HAC <=  GAC & ile & fai  |  gac & ILE & fai  |  gac & ile & FAI  |  GAC & ILE & FAI  ;
 hbc <=  GAC & ile & fai  |  gac & ILE & fai  |  gac & ile & FAI  |  gac & ile & fai  ;
 HAB <=  GAB & ilc & ild  |  gab & ILC & ild  |  gab & ilc & ILD  |  GAB & ILC & ILD  ;
 hbb <=  GAB & ilc & ild  |  gab & ILC & ild  |  gab & ilc & ILD  |  gab & ilc & ild  ;
 HAA <=  GAA & ila & ilb  |  gaa & ILA & ilb  |  gaa & ila & ILB  |  GAA & ILA & ILB  ;
 hba <=  GAA & ila & ilb  |  gaa & ILA & ilb  |  gaa & ila & ILB  |  gaa & ila & ilb  ;
 HCE <=  GBE & gci & fcp  |  gbe & GCI & fcp  |  gbe & gci & FCP  |  GBE & GCI & FCP  ;
 hde <=  GBE & gci & fcp  |  gbe & GCI & fcp  |  gbe & gci & FCP  |  gbe & gci & fcp  ;
 HCF <= GCJ ; 
 HCB <=  GBA & gca & gcd  |  gba & GCA & gcd  |  gba & gca & GCD  |  GBA & GCA & GCD  ;
 hdb <=  GBA & gca & gcd  |  gba & GCA & gcd  |  gba & gca & GCD  |  gba & gca & gcd  ;
 HAD <=  GAD & ilf & ilg  |  gad & ILF & ilg  |  gad & ilf & ILG  |  GAD & ILF & ILG  ;
 hbd <=  GAD & ilf & ilg  |  gad & ILF & ilg  |  gad & ilf & ILG  |  gad & ilf & ilg  ;
 HCC <=  GCF & gbd & gcg  |  gcf & GBD & gcg  |  gcf & gbd & GCG  |  GCF & GBD & GCG  ;
 hdc <=  GCF & gbd & gcg  |  gcf & GBD & gcg  |  gcf & gbd & GCG  |  gcf & gbd & gcg  ;
 HCD <=  GCE & gbc & gch  |  gce & GBC & gch  |  gce & gbc & GCH  |  GCE & GBC & GCH  ;
 hdd <=  GCE & gbc & gch  |  gce & GBC & gch  |  gce & gbc & GCH  |  gce & gbc & gch  ;
 HCA <=  GCB & gbb & gcc  |  gcb & GBB & gcc  |  gcb & gbb & GCC  |  GCB & GBB & GCC  ;
 hda <=  GCB & gbb & gcc  |  gcb & GBB & gcc  |  gcb & gbb & GCC  |  gcb & gbb & gcc  ;
 HEC <=  GDF & gef & gec  |  gdf & GEF & gec  |  gdf & gef & GEC  |  GDF & GEF & GEC  ;
 hfc <=  GDF & gef & gec  |  gdf & GEF & gec  |  gdf & gef & GEC  |  gdf & gef & gec  ;
 HEA <=  GDB & geb & gdc  |  gdb & GEB & gdc  |  gdb & geb & GDC  |  GDB & GEB & GDC  ;
 hfa <=  GDB & geb & gdc  |  gdb & GEB & gdc  |  gdb & geb & GDC  |  gdb & geb & gdc  ;
 HEB <=  GDA & gea & gdd  |  gda & GEA & gdd  |  gda & gea & GDD  |  GDA & GEA & GDD  ;
 hfb <=  GDA & gea & gdd  |  gda & GEA & gdd  |  gda & gea & GDD  |  gda & gea & gdd  ;
 HEE <=  GEH & gdi & gei  |  geh & GDI & gei  |  geh & gdi & GEI  |  GEH & GDI & GEI  ;
 hfe <=  GEH & gdi & gei  |  geh & GDI & gei  |  geh & gdi & GEI  |  geh & gdi & gei  ;
 HED <=  GEE & gde & ged  |  gee & GDE & ged  |  gee & gde & GED  |  GEE & GDE & GED  ;
 hfd <=  GEE & gde & ged  |  gee & GDE & ged  |  gee & gde & GED  |  gee & gde & ged  ;
 HEH <= GDJ ; 
 HEF <=  GDG & geg & gej  |  gdg & GEG & gej  |  gdg & geg & GEJ  |  GDG & GEG & GEJ  ;
 hff <=  GDG & geg & gej  |  gdg & GEG & gej  |  gdg & geg & GEJ  |  gdg & geg & gej  ;
 HEG <= GDH ; 
 HQC <=  GPC & gpe & gqe  |  gpc & GPE & gqe  |  gpc & gpe & GQE  |  GPC & GPE & GQE  ;
 ohc <=  GPC & gpe & gqe  |  gpc & GPE & gqe  |  gpc & gpe & GQE  |  gpc & gpe & gqe  ;
 HGA <=  GFB & ggb & gfc  |  gfb & GGB & gfc  |  gfb & ggb & GFC  |  GFB & GGB & GFC  ;
 hha <=  GFB & ggb & gfc  |  gfb & GGB & gfc  |  gfb & ggb & GFC  |  gfb & ggb & gfc  ;
 HGB <=  GFA & gga & gfd  |  gfa & GGA & gfd  |  gfa & gga & GFD  |  GFA & GGA & GFD  ;
 hhb <=  GFA & gga & gfd  |  gfa & GGA & gfd  |  gfa & gga & GFD  |  gfa & gga & gfd  ;
 HGE <=  GFH & ggh & ggg  |  gfh & GGH & ggg  |  gfh & ggh & GGG  |  GFH & GGH & GGG  ;
 hhe <=  GFH & ggh & ggg  |  gfh & GGH & ggg  |  gfh & ggh & GGG  |  gfh & ggh & ggg  ;
 HGF <=  GFG & gfj & ggj  |  gfg & GFJ & ggj  |  gfg & gfj & GGJ  |  GFG & GFJ & GGJ  ;
 hhf <=  GFG & gfj & ggj  |  gfg & GFJ & ggj  |  gfg & gfj & GGJ  |  gfg & gfj & ggj  ;
 HGC <=  GFF & ggf & ggc  |  gff & GGF & ggc  |  gff & ggf & GGC  |  GFF & GGF & GGC  ;
 hhc <=  GFF & ggf & ggc  |  gff & GGF & ggc  |  gff & ggf & GGC  |  gff & ggf & ggc  ;
 CCA <= IEK ; 
 CFA <= IEK ; 
 CCB <= IEL ; 
 CFB <= IEL ; 
 CCC <= IEM ; 
 CFC <= IEM ; 
 CCD <= IEN ; 
 CFD <= IEN ; 
 HQB <=  GQA & gpd & gqd  |  gqa & GPD & gqd  |  gqa & gpd & GQD  |  GQA & GPD & GQD  ;
 ohb <=  GQA & gpd & gqd  |  gqa & GPD & gqd  |  gqa & gpd & GQD  |  gqa & gpd & gqd  ;
 OHG <=  GRB & grd & gra  |  grb & GRD & gra  |  grb & grd & GRA  |  GRB & GRD & GRA  ;
 oig <=  GRB & grd & gra  |  grb & GRD & gra  |  grb & grd & GRA  |  grb & grd & gra  ;
 HQE <=  GQF & gpg & gqg  |  gqf & GPG & gqg  |  gqf & gpg & GQG  |  GQF & GPG & GQG  ;
 ohe <=  GQF & gpg & gqg  |  gqf & GPG & gqg  |  gqf & gpg & GQG  |  gqf & gpg & gqg  ;
 HQD <=  GQC & gpf & fqe  |  gqc & GPF & fqe  |  gqc & gpf & FQE  |  GQC & GPF & FQE  ;
 ohd <=  GQC & gpf & fqe  |  gqc & GPF & fqe  |  gqc & gpf & FQE  |  gqc & gpf & fqe  ;
 HQA <=  GPA & gpb & gqb  |  gpa & GPB & gqb  |  gpa & gpb & GQB  |  GPA & GPB & GQB  ;
 oha <=  GPA & gpb & gqb  |  gpa & GPB & gqb  |  gpa & gpb & GQB  |  gpa & gpb & gqb  ;
 OHJ <= GRC ; 
 OHH <=  GRF & grh & grg  |  grf & GRH & grg  |  grf & grh & GRG  |  GRF & GRH & GRG  ;
 oih <=  GRF & grh & grg  |  grf & GRH & grg  |  grf & grh & GRG  |  grf & grh & grg  ;
 OHI <= GRE ; 
 CCE <= IEO ; 
 CFE <= IEO ; 
 CCF <= IEP ; 
 CFF <= IEP ; 
 CCG <= IEQ ; 
 CFG <= IEQ ; 
 CCH <= IER ; 
 CFH <= IER ; 
 CCI <= IES ; 
 CFI <= IES ; 
 CCJ <= IET ; 
 CFJ <= IET ; 
 MIA <=  LHA & lia & khc  |  lha & LIA & khc  |  lha & lia & KHC  |  LHA & LIA & KHC  ;
 mja <=  LHA & lia & khc  |  lha & LIA & khc  |  lha & lia & KHC  |  lha & lia & khc  ;
 MIB <= LIB ; 
 MKA <=  LJA & lka & kjc  |  lja & LKA & kjc  |  lja & lka & KJC  |  LJA & LKA & KJC  ;
 mla <=  LJA & lka & kjc  |  lja & LKA & kjc  |  lja & lka & KJC  |  lja & lka & kjc  ;
 MKB <= LKB ; 
 MMA <=  LLA & lma & klc  |  lla & LMA & klc  |  lla & lma & KLC  |  LLA & LMA & KLC  ;
 mna <=  LLA & lma & klc  |  lla & LMA & klc  |  lla & lma & KLC  |  lla & lma & klc  ;
 MMB <= LMB ; 
 KQA <=  JQA & jpa & hpb  |  jqa & JPA & hpb  |  jqa & jpa & HPB  |  JQA & JPA & HPB  ;
 oka <=  JQA & jpa & hpb  |  jqa & JPA & hpb  |  jqa & jpa & HPB  |  jqa & jpa & hpb  ;
 KQB <=  JPB & jqb & jpc  |  jpb & JQB & jpc  |  jpb & jqb & JPC  |  JPB & JQB & JPC  ;
 okb <=  JPB & jqb & jpc  |  jpb & JQB & jpc  |  jpb & jqb & JPC  |  jpb & jqb & jpc  ;
 KOA <=  JOD & jnd & jnc  |  jod & JND & jnc  |  jod & jnd & JNC  |  JOD & JND & JNC  ;
 kpa <=  JOD & jnd & jnc  |  jod & JND & jnc  |  jod & jnd & JNC  |  jod & jnd & jnc  ;
 KOD <= JNA ; 
 KOB <=  JOB & jnb & joc  |  job & JNB & joc  |  job & jnb & JOC  |  JOB & JNB & JOC  ;
 kpb <=  JOB & jnb & joc  |  job & JNB & joc  |  job & jnb & JOC  |  job & jnb & joc  ;
 KOC <= JOA ; 
 OKD <=  JRA & jrb & jrc  |  jra & JRB & jrc  |  jra & jrb & JRC  |  JRA & JRB & JRC  ;
 old <=  JRA & jrb & jrc  |  jra & JRB & jrc  |  jra & jrb & JRC  |  jra & jrb & jrc  ;
 OKE <= JRD ; 
 KQC <=  JQD & jpd & jqc  |  jqd & JPD & jqc  |  jqd & jpd & JQC  |  JQD & JPD & JQC  ;
 okc <=  JQD & jpd & jqc  |  jqd & JPD & jqc  |  jqd & jpd & JQC  |  jqd & jpd & jqc  ;
 OAB <=  ICB & TSD  |  BAA & TKD  |  AAB & THD  ; 
 OBB <=  ICA & TSD  |  BAA & TKD  |  AAB & THD  ; 
 OAC <=  ICC & TSE  |  BAC & TKE  |  AAC & THE  ; 
 OBC <=  ICC & TSE  |  BAC & TKE  |  AAC & THE  ; 
 OAD <=  ICD & TSF  |  BAD & TKF  |  AAD & THF  ; 
 OBD <=  ICD & TSF  |  BAD & TKF  |  AAD & THF  ; 
 OAF <=  ICF & TSD  |  BAF & TKD  |  AAF & THD  ; 
 OBF <=  ICF & TSD  |  BAF & TKD  |  AAF & THD  ; 
 OAA <=  ICA & TSC  |  BAA & TKC  |  AAA & THC  ; 
 OBA <=  ICA & TSC  |  BAA & TKC  |  AAA & THC  ; 
 OAE <=  ICE & TSC  |  BAE & TKC  |  AAE & THC  ; 
 OBE <=  ICE & TSC  |  BAE & TKC  |  AAE & THC  ; 
 OAI <=  ICI & TSC  |  BAI & TKC  |  AAI & THC  ; 
 OBI <=  ICI & TSC  |  BAI & TKC  |  AAI & THC  ; 
 OAM <=  ICM & TSC  |  BAM & TKC  |  AAM & THC  ; 
 OBM <=  ICM & TSC  |  BAM & TKC  |  AAM & THC  ; 
 KAD <=  IMG & imh & imi  |  img & IMH & imi  |  img & imh & IMI  |  IMG & IMH & IMI  ;
 kbd <=  IMG & imh & imi  |  img & IMH & imi  |  img & imh & IMI  |  img & imh & imi  ;
 KAE <= IMJ ; 
 HAG <=  ILL & ilm & iln  |  ill & ILM & iln  |  ill & ilm & ILN  |  ILL & ILM & ILN  ;
 hbg <=  ILL & ilm & iln  |  ill & ILM & iln  |  ill & ilm & ILN  |  ill & ilm & iln  ;
 HAH <= ILO ; 
 HAF <=  ILI & ilj & ilk  |  ili & ILJ & ilk  |  ili & ilj & ILK  |  ILI & ILJ & ILK  ;
 hbf <=  ILI & ilj & ilk  |  ili & ILJ & ilk  |  ili & ilj & ILK  |  ili & ilj & ilk  ;
 HAI <= ILP ; 
 KAB <=  JAC & imc & imd  |  jac & IMC & imd  |  jac & imc & IMD  |  JAC & IMC & IMD  ;
 kbb <=  JAC & imc & imd  |  jac & IMC & imd  |  jac & imc & IMD  |  jac & imc & imd  ;
 KAC <=  JAB & ime & imf  |  jab & IME & imf  |  jab & ime & IMF  |  JAB & IME & IMF  ;
 kbc <=  JAB & ime & imf  |  jab & IME & imf  |  jab & ime & IMF  |  jab & ime & imf  ;
 KAF <= IMK ; 
 KAA <=  JAA & ima & imb  |  jaa & IMA & imb  |  jaa & ima & IMB  |  JAA & IMA & IMB  ;
 kba <=  JAA & ima & imb  |  jaa & IMA & imb  |  jaa & ima & IMB  |  jaa & ima & imb  ;
 KCB <=  JCC & jbc & jcd  |  jcc & JBC & jcd  |  jcc & jbc & JCD  |  JCC & JBC & JCD  ;
 kdb <=  JCC & jbc & jcd  |  jcc & JBC & jcd  |  jcc & jbc & JCD  |  jcc & jbc & jcd  ;
 KCE <= HBB ; 
 KCA <=  JCA & jba & iml  |  jca & JBA & iml  |  jca & jba & IML  |  JCA & JBA & IML  ;
 kda <=  JCA & jba & iml  |  jca & JBA & iml  |  jca & jba & IML  |  jca & jba & iml  ;
 KCC <=  JBB & jcb & imm  |  jbb & JCB & imm  |  jbb & jcb & IMM  |  JBB & JCB & IMM  ;
 kdc <=  JBB & jcb & imm  |  jbb & JCB & imm  |  jbb & jcb & IMM  |  jbb & jcb & imm  ;
 KCD <= IMN ; 
 KEC <=  JEB & jdb & jed  |  jeb & JDB & jed  |  jeb & jdb & JED  |  JEB & JDB & JED  ;
 kfc <=  JEB & jdb & jed  |  jeb & JDB & jed  |  jeb & jdb & JED  |  jeb & jdb & jed  ;
 KEA <=  JEA & jda & hda  |  jea & JDA & hda  |  jea & jda & HDA  |  JEA & JDA & HDA  ;
 kfa <=  JEA & jda & hda  |  jea & JDA & hda  |  jea & jda & HDA  |  jea & jda & hda  ;
 KEB <=  JDC & jec & jdd  |  jdc & JEC & jdd  |  jdc & jec & JDD  |  JDC & JEC & JDD  ;
 kfb <=  JDC & jec & jdd  |  jdc & JEC & jdd  |  jdc & jec & JDD  |  jdc & jec & jdd  ;
 KGC <=  JGB & jfb & jgd  |  jgb & JFB & jgd  |  jgb & jfb & JGD  |  JGB & JFB & JGD  ;
 khc <=  JGB & jfb & jgd  |  jgb & JFB & jgd  |  jgb & jfb & JGD  |  jgb & jfb & jgd  ;
 KGA <=  JGA & jfa & hfa  |  jga & JFA & hfa  |  jga & jfa & HFA  |  JGA & JFA & HFA  ;
 kha <=  JGA & jfa & hfa  |  jga & JFA & hfa  |  jga & jfa & HFA  |  jga & jfa & hfa  ;
 KGB <=  JFC & jgc & jfd  |  jfc & JGC & jfd  |  jfc & jgc & JFD  |  JFC & JGC & JFD  ;
 khb <=  JFC & jgc & jfd  |  jfc & JGC & jfd  |  jfc & jgc & JFD  |  jfc & jgc & jfd  ;
 KIB <=  JIC & jid & jhd  |  jic & JID & jhd  |  jic & jid & JHD  |  JIC & JID & JHD  ;
 kjb <=  JIC & jid & jhd  |  jic & JID & jhd  |  jic & jid & JHD  |  jic & jid & jhd  ;
 KIA <=  JIA & jha & hha  |  jia & JHA & hha  |  jia & jha & HHA  |  JIA & JHA & HHA  ;
 kja <=  JIA & jha & hha  |  jia & JHA & hha  |  jia & jha & HHA  |  jia & jha & hha  ;
 KIC <=  JIB & jhb & hhd  |  jib & JHB & hhd  |  jib & jhb & HHD  |  JIB & JHB & HHD  ;
 kjc <=  JIB & jhb & hhd  |  jib & JHB & hhd  |  jib & jhb & HHD  |  jib & jhb & hhd  ;
 KID <= JHC ; 
 KKA <=  JKA & jja & jkb  |  jka & JJA & jkb  |  jka & jja & JKB  |  JKA & JJA & JKB  ;
 kla <=  JKA & jja & jkb  |  jka & JJA & jkb  |  jka & jja & JKB  |  jka & jja & jkb  ;
 KKB <=  JJC & jkd & jjd  |  jjc & JKD & jjd  |  jjc & jkd & JJD  |  JJC & JKD & JJD  ;
 klb <=  JJC & jkd & jjd  |  jjc & JKD & jjd  |  jjc & jkd & JJD  |  jjc & jkd & jjd  ;
 KKC <=  JJB & jkc & hje  |  jjb & JKC & hje  |  jjb & jkc & HJE  |  JJB & JKC & HJE  ;
 klc <=  JJB & jkc & hje  |  jjb & JKC & hje  |  jjb & jkc & HJE  |  jjb & jkc & hje  ;
 KKD <= HJF ; 
 KMB <=  JMD & jld & hme  |  jmd & JLD & hme  |  jmd & jld & HME  |  JMD & JLD & HME  ;
 knb <=  JMD & jld & hme  |  jmd & JLD & hme  |  jmd & jld & HME  |  jmd & jld & hme  ;
 KMC <=  JMB & jlb & jmc  |  jmb & JLB & jmc  |  jmb & jlb & JMC  |  JMB & JLB & JMC  ;
 knc <=  JMB & jlb & jmc  |  jmb & JLB & jmc  |  jmb & jlb & JMC  |  jmb & jlb & jmc  ;
 KMD <= JLC ; 
 KMA <=  JLA & jma & hla  |  jla & JMA & hla  |  jla & jma & HLA  |  JLA & JMA & HLA  ;
 kna <=  JLA & jma & hla  |  jla & JMA & hla  |  jla & jma & HLA  |  jla & jma & hla  ;
 MQA <=  KQA & lpa & kqb  |  kqa & LPA & kqb  |  kqa & lpa & KQB  |  KQA & LPA & KQB  ;
 oma <=  KQA & lpa & kqb  |  kqa & LPA & kqb  |  kqa & lpa & KQB  |  kqa & lpa & kqb  ;
 MQB <= LQA ; 
 OAK <=  ICK & TSE  |  BAK & TKE  |  AAK & THE  ; 
 OBK <=  ICK & TSE  |  BAK & TKE  |  AAK & THE  ; 
 CCK <= IEU ; 
 CFK <= IEU ; 
 CCL <= IEV ; 
 CFL <= IEV ; 
 MOA <=  KNC & lob & lnb  |  knc & LOB & lnb  |  knc & lob & LNB  |  KNC & LOB & LNB  ;
 mpa <=  KNC & lob & lnb  |  knc & LOB & lnb  |  knc & lob & LNB  |  knc & lob & lnb  ;
 MOB <= LOA ; 
 CCM <= IEW ; 
 CFM <= IEW ; 
 CCN <= IEX ; 
 CFN <= IEX ; 
 MAA <=  LAA & ina & inb  |  laa & INA & inb  |  laa & ina & INB  |  LAA & INA & INB  ;
 mba <=  LAA & ina & inb  |  laa & INA & inb  |  laa & ina & INB  |  laa & ina & inb  ;
 MAC <= INE ; 
 CCO <= IEY ; 
 CFO <= IEY ; 
 CCP <= IEZ ; 
 CFP <= IEZ ; 
 MAB <=  LAB & inc & ind  |  lab & INC & ind  |  lab & inc & IND  |  LAB & INC & IND  ;
 mbb <=  LAB & inc & ind  |  lab & INC & ind  |  lab & inc & IND  |  lab & inc & ind  ;
 MAD <= INF ; 
 MCA <=  LCA & lba & lcc  |  lca & LBA & lcc  |  lca & lba & LCC  |  LCA & LBA & LCC  ;
 mda <=  LCA & lba & lcc  |  lca & LBA & lcc  |  lca & lba & LCC  |  lca & lba & lcc  ;
 OAO <=  ICO & TSE  |  BAO & TKE  |  AAO & THE  ; 
 OBO <=  ICO & TSE  |  BAO & TKE  |  AAO & THE  ; 
 OAP <=  ICP & TSF  |  BAP & TKF  |  AAP & THF  ; 
 OBP <=  ICP & TSF  |  BAP & TKF  |  AAP & THF  ; 
 MCB <=  LCB & lbb & ing  |  lcb & LBB & ing  |  lcb & lbb & ING  |  LCB & LBB & ING  ;
 mdb <=  LCB & lbb & ing  |  lcb & LBB & ing  |  lcb & lbb & ING  |  lcb & lbb & ing  ;
 OAL <=  ICL & TSF  |  BAL & TKF  |  AAL & THF  ; 
 OBL <=  ICL & TSF  |  BAL & TKF  |  AAL & THF  ; 
 OAN <=  ICN & TSD  |  BAN & TKD  |  AAN & THD  ; 
 OBN <=  ICN & TSD  |  BAM & TKD  |  AAN & THD  ; 
 OAG <=  ICG & TSE  |  BAG & TKE  |  AAG & THE  ; 
 OBG <=  ICG & TSE  |  BAG & TKE  |  AAG & THE  ; 
 MEA <=  LEA & lda & ldc  |  lea & LDA & ldc  |  lea & lda & LDC  |  LEA & LDA & LDC  ;
 mfa <=  LEA & lda & ldc  |  lea & LDA & ldc  |  lea & lda & LDC  |  lea & lda & ldc  ;
 MGA <=  LGA & lfa & lgb  |  lga & LFA & lgb  |  lga & lfa & LGB  |  LGA & LFA & LGB  ;
 mha <=  LGA & lfa & lgb  |  lga & LFA & lgb  |  lga & lfa & LGB  |  lga & lfa & lgb  ;
 MGB <= LFB ; 
 OAH <=  ICH & TSF  |  BAH & TKF  |  AAH & THF  ; 
 OBH <=  ICH & TSF  |  BAH & TKF  |  AAH & THF  ; 
 OAJ <=  ICJ & TSD  |  BAJ & TKD  |  AAJ & THD  ; 
 OBJ <=  ICJ & TSD  |  BAJ & TKD  |  AAJ & THD  ; 
end 
endmodule;
