module ja( IZZ,
 IAA, 
 IAB, 
 IAC, 
 IAD, 
 IAE, 
 IAF, 
 IAG, 
 IAH, 
 IAI, 
 IAJ, 
 IAK, 
 IAL, 
 IAM, 
 IAN, 
 IAO, 
 IAP, 
 IBA, 
 IBB, 
 IBC, 
 IBD, 
 IBE, 
 IBF, 
 IBG, 
 IBH, 
 IBI, 
 IBJ, 
 IBK, 
 IBL, 
 IBM, 
 IBN, 
 IBO, 
 IBP, 
 ICA, 
 ICB, 
 ICC, 
 ICD, 
 ICE, 
 ICF, 
 ICG, 
 ICH, 
 ICI, 
 ICJ, 
 ICK, 
 ICL, 
 ICM, 
 ICN, 
 ICO, 
 ICP, 
 IDA, 
 IDB, 
 IDC, 
 IDD, 
 IDE, 
 IDF, 
 IDG, 
 IDH, 
 IDI, 
 IDJ, 
 IDK, 
 IDL, 
 IDM, 
 IDN, 
 IDO, 
 IDP, 
 IEA, 
 IEB, 
 IEC, 
 IED, 
 IEE, 
 IEF, 
 IEG, 
 IEH, 
 IFA, 
 IFB, 
 IFC, 
 IFD, 
 IGA, 
 IGB, 
 IJA, 
 IJB, 
 IJC, 
 IJD, 
 IJE, 
 IJJ, 
 IJK, 
 IKA, 
 IKB, 
 IKC, 
 IKQ, 
 ILA, 
 OAA, 
 OAB, 
 OAC, 
 OAD, 
 OAE, 
 OAF, 
 OAG, 
 OAH, 
 OAI, 
 OAJ, 
 OAK, 
 OAL, 
 OAM, 
 OAN, 
 OAO, 
 OAP, 
 OBA, 
 OBB, 
 OBC, 
 OBD, 
 OBE, 
 OBF, 
 OBG, 
 OBH, 
 OBI, 
 OBJ, 
 OBK, 
 OBL, 
 OBM, 
 OBN, 
 OBO, 
 OBP, 
 OCA, 
 OCB, 
 OCC, 
 OCD, 
 OCE, 
 OCF, 
 OCG, 
 OCH, 
 OCI, 
 OCJ, 
 OCK, 
 OCL, 
 OCM, 
 OCN, 
 OCO, 
 OCP, 
 ODA, 
 ODB, 
 ODC, 
 ODD, 
 ODE, 
 ODF, 
 ODG, 
 ODH, 
 ODI, 
 ODJ, 
 OEA, 
 OEB, 
 OEC, 
 OED, 
 OEE, 
 OEF, 
 OFA, 
 OFB, 
 OFC, 
 OFD, 
 OFE, 
 OFF, 
 OGA, 
 OGB, 
 OGC, 
 OHA, 
 OHB, 
 OHC, 
 OHD, 
 OHE, 
 OHF, 
 OHG, 
 OIA, 
 OIB, 
 OJA, 
 OJB, 
 OJC, 
 OJD, 
 OKA, 
 OLA, 
 OLB, 
 OLC, 
 OLD, 
 OLE, 
 OLF, 
 OLG, 
 OLH, 
 OMA, 
 OMB, 
 ONA, 
 ONB, 
 OOA, 
 OOB, 
 OOC, 
 OOD, 
 OOE, 
 OOF, 
 OPA, 
 OPB, 
 OPC, 
 OPD, 
 OQA, 
 OQB, 
 OQC, 
 ORA, 
 ORB, 
 ORC, 
 ORD, 
 OSA, 
 OSB, 
 OSC, 
 OSD, 
 OSE, 
 OTA, 
 OTB, 
 OTC, 
 OTD, 
 OTE, 
 OTF, 
 OTG, 
 OUA, 
 OUB, 
 OUC, 
 OUD, 
 OUE, 
 OVA, 
 OVB, 
 OVC, 
 OVD, 
 OVE, 
 OVF, 
 OWA, 
 OWB, 
 OWC, 
 OWD, 
 OWE, 
 OWF, 
 OWG, 
 OWH, 
 OWI, 
 OWJ, 
 OWK, 
 OWL, 
 OWM, 
 OWN, 
 OWO, 
 OWP, 
 OWQ, 
 OWR, 
 OWS, 
 OWT, 
 OWU, 
 OWV, 
 OWW, 
 OWX, 
 OXA, 
 OXB, 
 OXC, 
OZA ); 
    
 input IZZ; 
 input IAA; 
 input IAB; 
 input IAC; 
 input IAD; 
 input IAE; 
 input IAF; 
 input IAG; 
 input IAH; 
 input IAI; 
 input IAJ; 
 input IAK; 
 input IAL; 
 input IAM; 
 input IAN; 
 input IAO; 
 input IAP; 
 input IBA; 
 input IBB; 
 input IBC; 
 input IBD; 
 input IBE; 
 input IBF; 
 input IBG; 
 input IBH; 
 input IBI; 
 input IBJ; 
 input IBK; 
 input IBL; 
 input IBM; 
 input IBN; 
 input IBO; 
 input IBP; 
 input ICA; 
 input ICB; 
 input ICC; 
 input ICD; 
 input ICE; 
 input ICF; 
 input ICG; 
 input ICH; 
 input ICI; 
 input ICJ; 
 input ICK; 
 input ICL; 
 input ICM; 
 input ICN; 
 input ICO; 
 input ICP; 
 input IDA; 
 input IDB; 
 input IDC; 
 input IDD; 
 input IDE; 
 input IDF; 
 input IDG; 
 input IDH; 
 input IDI; 
 input IDJ; 
 input IDK; 
 input IDL; 
 input IDM; 
 input IDN; 
 input IDO; 
 input IDP; 
 input IEA; 
 input IEB; 
 input IEC; 
 input IED; 
 input IEE; 
 input IEF; 
 input IEG; 
 input IEH; 
 input IFA; 
 input IFB; 
 input IFC; 
 input IFD; 
 input IGA; 
 input IGB; 
 input IJA; 
 input IJB; 
 input IJC; 
 input IJD; 
 input IJE; 
 input IJJ; 
 input IJK; 
 input IKA; 
 input IKB; 
 input IKC; 
 input IKQ; 
 input ILA; 
 output OAA; 
 output OAB; 
 output OAC; 
 output OAD; 
 output OAE; 
 output OAF; 
 output OAG; 
 output OAH; 
 output OAI; 
 output OAJ; 
 output OAK; 
 output OAL; 
 output OAM; 
 output OAN; 
 output OAO; 
 output OAP; 
 output OBA; 
 output OBB; 
 output OBC; 
 output OBD; 
 output OBE; 
 output OBF; 
 output OBG; 
 output OBH; 
 output OBI; 
 output OBJ; 
 output OBK; 
 output OBL; 
 output OBM; 
 output OBN; 
 output OBO; 
 output OBP; 
 output OCA; 
 output OCB; 
 output OCC; 
 output OCD; 
 output OCE; 
 output OCF; 
 output OCG; 
 output OCH; 
 output OCI; 
 output OCJ; 
 output OCK; 
 output OCL; 
 output OCM; 
 output OCN; 
 output OCO; 
 output OCP; 
 output ODA; 
 output ODB; 
 output ODC; 
 output ODD; 
 output ODE; 
 output ODF; 
 output ODG; 
 output ODH; 
 output ODI; 
 output ODJ; 
 output OEA; 
 output OEB; 
 output OEC; 
 output OED; 
 output OEE; 
 output OEF; 
 output OFA; 
 output OFB; 
 output OFC; 
 output OFD; 
 output OFE; 
 output OFF; 
 output OGA; 
 output OGB; 
 output OGC; 
 output OHA; 
 output OHB; 
 output OHC; 
 output OHD; 
 output OHE; 
 output OHF; 
 output OHG; 
 output OIA; 
 output OIB; 
 output OJA; 
 output OJB; 
 output OJC; 
 output OJD; 
 output OKA; 
 output OLA; 
 output OLB; 
 output OLC; 
 output OLD; 
 output OLE; 
 output OLF; 
 output OLG; 
 output OLH; 
 output OMA; 
 output OMB; 
 output ONA; 
 output ONB; 
 output OOA; 
 output OOB; 
 output OOC; 
 output OOD; 
 output OOE; 
 output OOF; 
 output OPA; 
 output OPB; 
 output OPC; 
 output OPD; 
 output OQA; 
 output OQB; 
 output OQC; 
 output ORA; 
 output ORB; 
 output ORC; 
 output ORD; 
 output OSA; 
 output OSB; 
 output OSC; 
 output OSD; 
 output OSE; 
 output OTA; 
 output OTB; 
 output OTC; 
 output OTD; 
 output OTE; 
 output OTF; 
 output OTG; 
 output OUA; 
 output OUB; 
 output OUC; 
 output OUD; 
 output OUE; 
 output OVA; 
 output OVB; 
 output OVC; 
 output OVD; 
 output OVE; 
 output OVF; 
 output OWA; 
 output OWB; 
 output OWC; 
 output OWD; 
 output OWE; 
 output OWF; 
 output OWG; 
 output OWH; 
 output OWI; 
 output OWJ; 
 output OWK; 
 output OWL; 
 output OWM; 
 output OWN; 
 output OWO; 
 output OWP; 
 output OWQ; 
 output OWR; 
 output OWS; 
 output OWT; 
 output OWU; 
 output OWV; 
 output OWW; 
 output OWX; 
 output OXA; 
 output OXB; 
 output OXC; 
 output OZA; 
  
  
reg  AAA ;
reg  AAB ;
reg  AAC ;
reg  AAD ;
reg  AAE ;
reg  AAF ;
reg  AAG ;
reg  AAH ;
reg  AAI ;
reg  AAJ ;
reg  AAK ;
reg  AAL ;
reg  AAM ;
reg  AAN ;
reg  AAO ;
reg  AAP ;
reg  ABA ;
reg  ABB ;
reg  ABC ;
reg  ABD ;
reg  ABE ;
reg  ABF ;
reg  ABG ;
reg  ABH ;
reg  ABI ;
reg  ABJ ;
reg  ABK ;
reg  ABL ;
reg  ABM ;
reg  ABN ;
reg  ABO ;
reg  ABP ;
reg  ACA ;
reg  ACB ;
reg  ACC ;
reg  ACD ;
reg  ACE ;
reg  ACF ;
reg  ACG ;
reg  ACH ;
reg  ACI ;
reg  ACJ ;
reg  ACK ;
reg  ACL ;
reg  ACM ;
reg  ACN ;
reg  ACO ;
reg  ACP ;
reg  ADA ;
reg  ADB ;
reg  ADC ;
reg  ADD ;
reg  ADE ;
reg  ADF ;
reg  ADG ;
reg  ADH ;
reg  ADI ;
reg  ADJ ;
reg  ADK ;
reg  ADL ;
reg  ADM ;
reg  ADN ;
reg  ADO ;
reg  ADP ;
reg  cqa ;
reg  cqb ;
reg  cqc ;
reg  cqd ;
reg  cqe ;
reg  cqf ;
reg  cqg ;
reg  cqh ;
reg  cqi ;
reg  cqj ;
reg  cqk ;
reg  cql ;
reg  cqm ;
reg  cqn ;
reg  cqo ;
reg  cqp ;
reg  EAA ;
reg  EAB ;
reg  EAC ;
reg  EAD ;
reg  EAE ;
reg  EAF ;
reg  EAG ;
reg  EAH ;
reg  EAI ;
reg  EAK ;
reg  EAM ;
reg  EAN ;
reg  EAP ;
reg  EBA ;
reg  EBB ;
reg  EBC ;
reg  EBD ;
reg  EBE ;
reg  EBF ;
reg  EBG ;
reg  EBI ;
reg  EBJ ;
reg  EBK ;
reg  EBL ;
reg  EBM ;
reg  EBN ;
reg  ECA ;
reg  ECB ;
reg  ECC ;
reg  ECD ;
reg  ECE ;
reg  ECF ;
reg  ECG ;
reg  ECI ;
reg  ECJ ;
reg  ECK ;
reg  ECL ;
reg  ECM ;
reg  ecn ;
reg  ECO ;
reg  EDA ;
reg  EDB ;
reg  edc ;
reg  EDD ;
reg  ede ;
reg  EDF ;
reg  EDG ;
reg  EDH ;
reg  EDI ;
reg  EDJ ;
reg  EDK ;
reg  EDL ;
reg  EDM ;
reg  EDN ;
reg  EDO ;
reg  EDP ;
reg  EEA ;
reg  eeb ;
reg  EEC ;
reg  EED ;
reg  EEE ;
reg  EEF ;
reg  EEG ;
reg  EEI ;
reg  EEJ ;
reg  EEL ;
reg  EEM ;
reg  EEN ;
reg  EQA ;
reg  EQB ;
reg  EQC ;
reg  EQD ;
reg  EQE ;
reg  EQF ;
reg  EQG ;
reg  EQH ;
reg  EQI ;
reg  EQJ ;
reg  EQK ;
reg  EQL ;
reg  EQM ;
reg  EQN ;
reg  EQO ;
reg  EQP ;
reg  GAA ;
reg  GAB ;
reg  GAC ;
reg  GAD ;
reg  GAE ;
reg  GAF ;
reg  GAG ;
reg  GAH ;
reg  GBA ;
reg  GBB ;
reg  GBC ;
reg  GBD ;
reg  GBE ;
reg  GBF ;
reg  GBG ;
reg  GBH ;
reg  GCA ;
reg  GCB ;
reg  GCC ;
reg  GCD ;
reg  GCE ;
reg  GCF ;
reg  GCG ;
reg  GCH ;
reg  GDA ;
reg  GDB ;
reg  GDC ;
reg  GDD ;
reg  GDE ;
reg  GDF ;
reg  GDG ;
reg  GDH ;
reg  GEA ;
reg  GEB ;
reg  GEC ;
reg  GED ;
reg  GEE ;
reg  GEF ;
reg  GEG ;
reg  GFA ;
reg  GFB ;
reg  GFC ;
reg  GFD ;
reg  GFE ;
reg  GFF ;
reg  GFI ;
reg  GGA ;
reg  GGB ;
reg  GGC ;
reg  GGD ;
reg  GGE ;
reg  GGF ;
reg  GGG ;
reg  GGH ;
reg  GHA ;
reg  GHB ;
reg  GHC ;
reg  GHD ;
reg  GHE ;
reg  GHF ;
reg  GHG ;
reg  GHH ;
reg  GIA ;
reg  GIB ;
reg  GIC ;
reg  GID ;
reg  GIE ;
reg  GIF ;
reg  GIG ;
reg  GIH ;
reg  GJA ;
reg  GJB ;
reg  GJC ;
reg  GJD ;
reg  GJE ;
reg  GJF ;
reg  GJG ;
reg  GJH ;
reg  GKA ;
reg  GKB ;
reg  GKC ;
reg  GKD ;
reg  GKE ;
reg  GKF ;
reg  GKG ;
reg  GLA ;
reg  GLB ;
reg  GLC ;
reg  GLD ;
reg  GLE ;
reg  GLF ;
reg  GLG ;
reg  GLH ;
reg  gqa ;
reg  gqb ;
reg  gqc ;
reg  gqd ;
reg  gqe ;
reg  gqf ;
reg  gqg ;
reg  gqh ;
reg  gqi ;
reg  gqj ;
reg  gqk ;
reg  gql ;
reg  gqm ;
reg  gqn ;
reg  gqo ;
reg  gqp ;
reg  HAA ;
reg  HAB ;
reg  HAC ;
reg  HAD ;
reg  HAE ;
reg  HAF ;
reg  HAG ;
reg  HAH ;
reg  HBA ;
reg  HBB ;
reg  HBC ;
reg  HBD ;
reg  HBE ;
reg  HBF ;
reg  HBG ;
reg  HBH ;
reg  HCA ;
reg  HCB ;
reg  HCC ;
reg  HCD ;
reg  HCE ;
reg  HCF ;
reg  HCG ;
reg  HCH ;
reg  HDA ;
reg  HDB ;
reg  HDC ;
reg  HDD ;
reg  HDE ;
reg  HDF ;
reg  HDG ;
reg  HDH ;
reg  hea ;
reg  heb ;
reg  hec ;
reg  hed ;
reg  hee ;
reg  hef ;
reg  HFA ;
reg  HFB ;
reg  HFC ;
reg  HFD ;
reg  HFE ;
reg  HFF ;
reg  HFG ;
reg  HFH ;
reg  HFI ;
reg  KAA ;
reg  KAB ;
reg  KAC ;
reg  KAD ;
reg  KAF ;
reg  KAG ;
reg  KBA ;
reg  KBB ;
reg  KBC ;
reg  KBD ;
reg  KBF ;
reg  KBG ;
reg  KCA ;
reg  KCB ;
reg  KCC ;
reg  KCD ;
reg  KCF ;
reg  KCG ;
reg  KDA ;
reg  KDB ;
reg  KDC ;
reg  KDD ;
reg  KDF ;
reg  KDG ;
reg  KEA ;
reg  KEB ;
reg  KEC ;
reg  KED ;
reg  KEF ;
reg  KEG ;
reg  KFA ;
reg  KFB ;
reg  KFC ;
reg  KFD ;
reg  KFE ;
reg  KFF ;
reg  KFG ;
reg  KGA ;
reg  KGB ;
reg  KGC ;
reg  KGD ;
reg  KGE ;
reg  KGF ;
reg  KGG ;
reg  KHA ;
reg  KHB ;
reg  KHC ;
reg  KHD ;
reg  KHE ;
reg  KHF ;
reg  KHG ;
reg  KIA ;
reg  KIB ;
reg  KIC ;
reg  KID ;
reg  KIE ;
reg  KIF ;
reg  KIG ;
reg  KJA ;
reg  KJB ;
reg  KJC ;
reg  KJD ;
reg  KJE ;
reg  KJF ;
reg  KJG ;
reg  KKA ;
reg  KKB ;
reg  KKC ;
reg  KKD ;
reg  KKE ;
reg  KKF ;
reg  KLA ;
reg  KLB ;
reg  KLC ;
reg  KLD ;
reg  KLE ;
reg  KLF ;
reg  LAA ;
reg  LAB ;
reg  LAC ;
reg  LBA ;
reg  LBB ;
reg  LBC ;
reg  lbg ;
reg  LCA ;
reg  LCB ;
reg  LCC ;
reg  LCD ;
reg  LCE ;
reg  LCF ;
reg  LCG ;
reg  LDA ;
reg  LDB ;
reg  LDC ;
reg  LDD ;
reg  LDE ;
reg  LDF ;
reg  LDG ;
reg  LEA ;
reg  LEB ;
reg  LEC ;
reg  LED ;
reg  LEE ;
reg  LEF ;
reg  LEG ;
reg  LFA ;
reg  LFB ;
reg  LFC ;
reg  LFD ;
reg  LFE ;
reg  LFF ;
reg  LFG ;
reg  LGA ;
reg  LGB ;
reg  LGC ;
reg  LGD ;
reg  LGE ;
reg  LGF ;
reg  LGG ;
reg  LHA ;
reg  LHB ;
reg  LHC ;
reg  LHD ;
reg  LHE ;
reg  LHF ;
reg  LHG ;
reg  LIA ;
reg  LIB ;
reg  LIC ;
reg  LID ;
reg  LIE ;
reg  LIF ;
reg  LIG ;
reg  LJA ;
reg  LJB ;
reg  LJC ;
reg  LJD ;
reg  LJE ;
reg  LJF ;
reg  LJG ;
reg  LKA ;
reg  LKB ;
reg  LKC ;
reg  LKD ;
reg  LKE ;
reg  LKF ;
reg  LKG ;
reg  LLA ;
reg  LLB ;
reg  LLC ;
reg  LLD ;
reg  LLE ;
reg  LLF ;
reg  LLG ;
reg  LMA ;
reg  LMB ;
reg  LMC ;
reg  LMD ;
reg  LME ;
reg  LMF ;
reg  LMG ;
reg  LNA ;
reg  LNB ;
reg  LNC ;
reg  LND ;
reg  LNE ;
reg  LNF ;
reg  LNG ;
reg  LOA ;
reg  LOB ;
reg  LOC ;
reg  LOD ;
reg  LOE ;
reg  LOF ;
reg  LOG ;
reg  LPA ;
reg  LPB ;
reg  LPC ;
reg  LPD ;
reg  LPE ;
reg  LPF ;
reg  LPG ;
reg  LQA ;
reg  LQB ;
reg  LQC ;
reg  LQD ;
reg  LQE ;
reg  LQF ;
reg  LQG ;
reg  LRA ;
reg  LRB ;
reg  LRC ;
reg  LRD ;
reg  LRE ;
reg  LRF ;
reg  LSA ;
reg  LSB ;
reg  LSC ;
reg  LSD ;
reg  LSE ;
reg  LSF ;
reg  naa ;
reg  nab ;
reg  nac ;
reg  nad ;
reg  NAG ;
reg  nca ;
reg  ncb ;
reg  ncc ;
reg  ncd ;
reg  nce ;
reg  ncf ;
reg  ncg ;
reg  nch ;
reg  nda ;
reg  ndb ;
reg  ndc ;
reg  ndd ;
reg  nde ;
reg  ndf ;
reg  ndg ;
reg  ndh ;
reg  ndi ;
reg  ndj ;
reg  ndk ;
reg  ndl ;
reg  nea ;
reg  neb ;
reg  nec ;
reg  nee ;
reg  nei ;
reg  nia ;
reg  nib ;
reg  nic ;
reg  NKA ;
reg  NKB ;
reg  NKC ;
reg  NKD ;
reg  NKE ;
reg  NKF ;
reg  NKG ;
reg  NKH ;
reg  NKI ;
reg  NKJ ;
reg  NKK ;
reg  NKL ;
reg  NKM ;
reg  NKN ;
reg  NKO ;
reg  NKP ;
reg  NKQ ;
reg  NKR ;
reg  NKS ;
reg  NKT ;
reg  nku ;
reg  NLA ;
reg  NLB ;
reg  NLC ;
reg  NLD ;
reg  NLE ;
reg  NLF ;
reg  NLG ;
reg  NLH ;
reg  oaa ;
reg  oab ;
reg  oac ;
reg  oad ;
reg  oae ;
reg  oaf ;
reg  oag ;
reg  oah ;
reg  oai ;
reg  oaj ;
reg  oak ;
reg  oal ;
reg  oam ;
reg  oan ;
reg  oao ;
reg  oap ;
reg  oba ;
reg  obb ;
reg  obc ;
reg  obd ;
reg  obe ;
reg  obf ;
reg  obg ;
reg  obh ;
reg  obi ;
reg  obj ;
reg  obk ;
reg  obl ;
reg  obm ;
reg  obn ;
reg  obo ;
reg  obp ;
reg  oca ;
reg  ocb ;
reg  occ ;
reg  ocd ;
reg  oce ;
reg  ocf ;
reg  ocg ;
reg  och ;
reg  oci ;
reg  ocj ;
reg  ock ;
reg  ocl ;
reg  ocm ;
reg  ocn ;
reg  oco ;
reg  ocp ;
reg  oda ;
reg  odb ;
reg  odc ;
reg  odd ;
reg  ode ;
reg  odf ;
reg  odg ;
reg  odh ;
reg  odi ;
reg  odj ;
reg  OEA ;
reg  OEB ;
reg  OEC ;
reg  OED ;
reg  OEE ;
reg  OEF ;
reg  OFA ;
reg  OFB ;
reg  OFC ;
reg  OFD ;
reg  OFE ;
reg  OFF ;
reg  OGA ;
reg  OGB ;
reg  OGC ;
reg  OHA ;
reg  OHB ;
reg  OHC ;
reg  OHD ;
reg  OHE ;
reg  OHF ;
reg  OHG ;
reg  OIA ;
reg  OIB ;
reg  oja ;
reg  ojb ;
reg  ojc ;
reg  OJD ;
reg  oka ;
reg  ola ;
reg  olb ;
reg  olc ;
reg  old ;
reg  ole ;
reg  olf ;
reg  olg ;
reg  olh ;
reg  OMA ;
reg  OMB ;
reg  ona ;
reg  onb ;
reg  OOA ;
reg  OOB ;
reg  OOC ;
reg  OOD ;
reg  OOE ;
reg  OOF ;
reg  opa ;
reg  OPB ;
reg  OPC ;
reg  opd ;
reg  oqa ;
reg  OQB ;
reg  OQC ;
reg  ora ;
reg  ORB ;
reg  ORC ;
reg  ORD ;
reg  osa ;
reg  OSB ;
reg  OSC ;
reg  OSD ;
reg  ose ;
reg  ota ;
reg  otb ;
reg  OTC ;
reg  otd ;
reg  OTE ;
reg  OTF ;
reg  OTG ;
reg  oua ;
reg  oub ;
reg  OUC ;
reg  OUD ;
reg  OUE ;
reg  ova ;
reg  OVB ;
reg  OVC ;
reg  OVD ;
reg  OVE ;
reg  OVF ;
reg  OWA ;
reg  OWB ;
reg  OWC ;
reg  OWD ;
reg  OWE ;
reg  OWF ;
reg  owg ;
reg  owh ;
reg  owi ;
reg  owj ;
reg  owk ;
reg  owl ;
reg  OWM ;
reg  OWN ;
reg  OWO ;
reg  owp ;
reg  OWQ ;
reg  owr ;
reg  OWS ;
reg  OWT ;
reg  owu ;
reg  owv ;
reg  oww ;
reg  owx ;
reg  OXA ;
reg  OXB ;
reg  OXC ;
reg  oza ;
reg  ozb ;
reg  PAA ;
reg  PAB ;
reg  PAC ;
reg  PAD ;
reg  PAE ;
reg  PAF ;
reg  PAG ;
reg  PAH ;
reg  PBA ;
reg  PBB ;
reg  PBC ;
reg  PBD ;
reg  PBE ;
reg  PBF ;
reg  PBG ;
reg  PBH ;
reg  PCA ;
reg  PCB ;
reg  PCC ;
reg  PCD ;
reg  PCE ;
reg  PCF ;
reg  PCG ;
reg  PDA ;
reg  PDB ;
reg  PDC ;
reg  PDD ;
reg  PDE ;
reg  PDF ;
reg  PDG ;
reg  PDH ;
reg  PEA ;
reg  PEB ;
reg  PEC ;
reg  PED ;
reg  PEE ;
reg  PEF ;
reg  PFA ;
reg  PFB ;
reg  PFC ;
reg  PFD ;
reg  PFE ;
reg  PFF ;
reg  PFG ;
reg  PFH ;
reg  PGA ;
reg  PGB ;
reg  PGC ;
reg  PGD ;
reg  PGE ;
reg  PGF ;
reg  PGG ;
reg  PHA ;
reg  PHB ;
reg  PHC ;
reg  PHD ;
reg  PHE ;
reg  PHF ;
reg  PHG ;
reg  PHH ;
reg  PIA ;
reg  PIB ;
reg  PIC ;
reg  PID ;
reg  PIE ;
reg  PJA ;
reg  PJC ;
reg  PJD ;
reg  PJE ;
reg  PJF ;
reg  PKA ;
reg  PKB ;
reg  PKC ;
reg  PKD ;
reg  PKE ;
reg  PKF ;
reg  PLA ;
reg  PLB ;
reg  PLC ;
reg  PLD ;
reg  PLE ;
reg  PLF ;
reg  PMA ;
reg  PMB ;
reg  PMC ;
reg  PMD ;
reg  PME ;
reg  PMF ;
reg  PNA ;
reg  PNB ;
reg  PNC ;
reg  PND ;
reg  PNE ;
reg  PNF ;
reg  POA ;
reg  POB ;
reg  POC ;
reg  POD ;
reg  POE ;
reg  POF ;
reg  qaa ;
reg  qab ;
reg  qac ;
reg  qad ;
reg  qae ;
reg  qaf ;
reg  qag ;
reg  qah ;
reg  qba ;
reg  qbb ;
reg  qbc ;
reg  qbd ;
reg  qbe ;
reg  qbf ;
reg  qbg ;
reg  qbh ;
reg  QCA ;
reg  QCB ;
reg  QCC ;
reg  QCD ;
reg  QCE ;
reg  qda ;
reg  qdb ;
reg  qdc ;
reg  qdd ;
reg  qea ;
reg  qeb ;
reg  qec ;
reg  qed ;
reg  qee ;
reg  qfa ;
reg  qfb ;
reg  qfc ;
reg  qfd ;
reg  qfe ;
reg  qff ;
reg  QGA ;
reg  QGB ;
reg  QGC ;
reg  qgd ;
reg  qge ;
reg  QHA ;
reg  QHB ;
reg  QHD ;
reg  QHF ;
reg  QHG ;
reg  QHI ;
reg  QHJ ;
reg  QHK ;
reg  QHL ;
reg  QIA ;
reg  QIB ;
reg  QIC ;
reg  QID ;
reg  qie ;
reg  QJA ;
reg  qka ;
reg  qkb ;
reg  QLA ;
reg  QLB ;
reg  QLC ;
reg  QMA ;
reg  QMB ;
reg  QMC ;
reg  QMD ;
reg  RAA ;
reg  RAB ;
reg  RAC ;
reg  RAD ;
reg  RAE ;
reg  RAF ;
reg  RAG ;
reg  RAH ;
reg  RAI ;
reg  RAJ ;
reg  RAK ;
reg  RAL ;
reg  RAM ;
reg  RAN ;
reg  RAO ;
reg  RAP ;
reg  RAQ ;
reg  RAR ;
reg  RAS ;
reg  RAT ;
reg  RAU ;
reg  RAV ;
reg  RAW ;
reg  RAX ;
reg  WAA ;
reg  WAB ;
reg  WAC ;
reg  WAD ;
reg  WAE ;
reg  WAF ;
reg  WAG ;
reg  WAH ;
reg  WBA ;
reg  WBB ;
reg  WBC ;
reg  WBD ;
reg  WBE ;
reg  WBF ;
reg  WBG ;
reg  WBH ;
reg  WCA ;
reg  WCB ;
reg  WCC ;
reg  WDA ;
reg  WDB ;
reg  WDC ;
wire  aaa ;
wire  aab ;
wire  aac ;
wire  aad ;
wire  aae ;
wire  aaf ;
wire  aag ;
wire  aah ;
wire  aai ;
wire  aaj ;
wire  aak ;
wire  aal ;
wire  aam ;
wire  aan ;
wire  aao ;
wire  aap ;
wire  aba ;
wire  abb ;
wire  abc ;
wire  abd ;
wire  abe ;
wire  abf ;
wire  abg ;
wire  abh ;
wire  abi ;
wire  abj ;
wire  abk ;
wire  abl ;
wire  abm ;
wire  abn ;
wire  abo ;
wire  abp ;
wire  aca ;
wire  acb ;
wire  acc ;
wire  acd ;
wire  ace ;
wire  acf ;
wire  acg ;
wire  ach ;
wire  aci ;
wire  acj ;
wire  ack ;
wire  acl ;
wire  acm ;
wire  acn ;
wire  aco ;
wire  acp ;
wire  ada ;
wire  adb ;
wire  adc ;
wire  add ;
wire  ade ;
wire  adf ;
wire  adg ;
wire  adh ;
wire  adi ;
wire  adj ;
wire  adk ;
wire  adl ;
wire  adm ;
wire  adn ;
wire  ado ;
wire  adp ;
wire  baa ;
wire  BAA ;
wire  bab ;
wire  BAB ;
wire  bac ;
wire  BAC ;
wire  bad ;
wire  BAD ;
wire  bae ;
wire  BAE ;
wire  baf ;
wire  BAF ;
wire  bag ;
wire  BAG ;
wire  bah ;
wire  BAH ;
wire  bba ;
wire  BBA ;
wire  bbb ;
wire  BBB ;
wire  bbc ;
wire  BBC ;
wire  bbd ;
wire  BBD ;
wire  bbe ;
wire  BBE ;
wire  bbf ;
wire  BBF ;
wire  bbg ;
wire  BBG ;
wire  bbh ;
wire  BBH ;
wire  bca ;
wire  BCA ;
wire  bcb ;
wire  BCB ;
wire  bcc ;
wire  BCC ;
wire  bcd ;
wire  BCD ;
wire  bce ;
wire  BCE ;
wire  bcf ;
wire  BCF ;
wire  bcg ;
wire  BCG ;
wire  bch ;
wire  BCH ;
wire  bda ;
wire  BDA ;
wire  bdb ;
wire  BDB ;
wire  bdc ;
wire  BDC ;
wire  bdd ;
wire  BDD ;
wire  bde ;
wire  BDE ;
wire  bdf ;
wire  BDF ;
wire  bdg ;
wire  BDG ;
wire  bdh ;
wire  BDH ;
wire  CQA ;
wire  CQB ;
wire  CQC ;
wire  CQD ;
wire  CQE ;
wire  CQF ;
wire  CQG ;
wire  CQH ;
wire  CQI ;
wire  CQJ ;
wire  CQK ;
wire  CQL ;
wire  CQM ;
wire  CQN ;
wire  CQO ;
wire  CQP ;
wire  daa ;
wire  DAA ;
wire  dab ;
wire  DAB ;
wire  dac ;
wire  DAC ;
wire  dad ;
wire  DAD ;
wire  daf ;
wire  DAF ;
wire  dag ;
wire  DAG ;
wire  dah ;
wire  DAH ;
wire  dai ;
wire  DAI ;
wire  daj ;
wire  DAJ ;
wire  dak ;
wire  DAK ;
wire  dal ;
wire  DAL ;
wire  dam ;
wire  DAM ;
wire  dan ;
wire  DAN ;
wire  dao ;
wire  DAO ;
wire  dap ;
wire  DAP ;
wire  daq ;
wire  DAQ ;
wire  dar ;
wire  DAR ;
wire  das ;
wire  DAS ;
wire  dat ;
wire  DAT ;
wire  dau ;
wire  DAU ;
wire  dav ;
wire  DAV ;
wire  daw ;
wire  DAW ;
wire  dba ;
wire  DBA ;
wire  dbb ;
wire  DBB ;
wire  dbc ;
wire  DBC ;
wire  dbd ;
wire  DBD ;
wire  dbe ;
wire  DBE ;
wire  dbf ;
wire  DBF ;
wire  dbg ;
wire  DBG ;
wire  dbh ;
wire  DBH ;
wire  dbi ;
wire  DBI ;
wire  dbj ;
wire  DBJ ;
wire  dbk ;
wire  DBK ;
wire  dbl ;
wire  DBL ;
wire  dbm ;
wire  DBM ;
wire  dbn ;
wire  DBN ;
wire  dbp ;
wire  DBP ;
wire  dbq ;
wire  DBQ ;
wire  dbs ;
wire  DBS ;
wire  dbt ;
wire  DBT ;
wire  dbu ;
wire  DBU ;
wire  dbv ;
wire  DBV ;
wire  dca ;
wire  DCA ;
wire  dcb ;
wire  DCB ;
wire  dcc ;
wire  DCC ;
wire  dcd ;
wire  DCD ;
wire  dce ;
wire  DCE ;
wire  dcf ;
wire  DCF ;
wire  dci ;
wire  DCI ;
wire  dcj ;
wire  DCJ ;
wire  dck ;
wire  DCK ;
wire  dcl ;
wire  DCL ;
wire  dcm ;
wire  DCM ;
wire  dcn ;
wire  DCN ;
wire  dcq ;
wire  DCQ ;
wire  dct ;
wire  DCT ;
wire  dcu ;
wire  DCU ;
wire  dcv ;
wire  DCV ;
wire  dcw ;
wire  DCW ;
wire  dda ;
wire  DDA ;
wire  ddb ;
wire  DDB ;
wire  ddc ;
wire  DDC ;
wire  ddd ;
wire  DDD ;
wire  dde ;
wire  DDE ;
wire  ddf ;
wire  DDF ;
wire  ddg ;
wire  DDG ;
wire  ddh ;
wire  DDH ;
wire  ddi ;
wire  DDI ;
wire  ddj ;
wire  DDJ ;
wire  ddk ;
wire  DDK ;
wire  ddl ;
wire  DDL ;
wire  ddm ;
wire  DDM ;
wire  ddn ;
wire  DDN ;
wire  ddo ;
wire  DDO ;
wire  ddp ;
wire  DDP ;
wire  dea ;
wire  DEA ;
wire  deb ;
wire  DEB ;
wire  dec ;
wire  DEC ;
wire  ded ;
wire  DED ;
wire  dee ;
wire  DEE ;
wire  def ;
wire  DEF ;
wire  dei ;
wire  DEI ;
wire  dej ;
wire  DEJ ;
wire  dek ;
wire  DEK ;
wire  del ;
wire  DEL ;
wire  dem ;
wire  DEM ;
wire  den ;
wire  DEN ;
wire  dfb ;
wire  DFB ;
wire  dfc ;
wire  DFC ;
wire  dfd ;
wire  DFD ;
wire  dfe ;
wire  DFE ;
wire  dff ;
wire  DFF ;
wire  dfg ;
wire  DFG ;
wire  dfj ;
wire  DFJ ;
wire  dfk ;
wire  DFK ;
wire  dfm ;
wire  DFM ;
wire  dfn ;
wire  DFN ;
wire  dgc ;
wire  DGC ;
wire  dge ;
wire  DGE ;
wire  dgk ;
wire  DGK ;
wire  dgm ;
wire  DGM ;
wire  eaa ;
wire  eab ;
wire  eac ;
wire  ead ;
wire  eae ;
wire  eaf ;
wire  eag ;
wire  eah ;
wire  eai ;
wire  eak ;
wire  eam ;
wire  ean ;
wire  eap ;
wire  eba ;
wire  ebb ;
wire  ebc ;
wire  ebd ;
wire  ebe ;
wire  ebf ;
wire  ebg ;
wire  ebi ;
wire  ebj ;
wire  ebk ;
wire  ebl ;
wire  ebm ;
wire  ebn ;
wire  eca ;
wire  ecb ;
wire  ecc ;
wire  ecd ;
wire  ece ;
wire  ecf ;
wire  ecg ;
wire  eci ;
wire  ecj ;
wire  eck ;
wire  ecl ;
wire  ecm ;
wire  ECN ;
wire  eco ;
wire  eda ;
wire  edb ;
wire  EDC ;
wire  edd ;
wire  EDE ;
wire  edf ;
wire  edg ;
wire  edh ;
wire  edi ;
wire  edj ;
wire  edk ;
wire  edl ;
wire  edm ;
wire  edn ;
wire  edo ;
wire  edp ;
wire  eea ;
wire  EEB ;
wire  eec ;
wire  eed ;
wire  eee ;
wire  eef ;
wire  eeg ;
wire  eei ;
wire  eej ;
wire  eel ;
wire  eem ;
wire  een ;
wire  eqa ;
wire  eqb ;
wire  eqc ;
wire  eqd ;
wire  eqe ;
wire  eqf ;
wire  eqg ;
wire  eqh ;
wire  eqi ;
wire  eqj ;
wire  eqk ;
wire  eql ;
wire  eqm ;
wire  eqn ;
wire  eqo ;
wire  eqp ;
wire  FAA ;
wire  FAB ;
wire  FAC ;
wire  FAD ;
wire  FAE ;
wire  FAF ;
wire  FAG ;
wire  FAH ;
wire  FBA ;
wire  FBB ;
wire  FBC ;
wire  FBD ;
wire  FBE ;
wire  FBF ;
wire  FBG ;
wire  FBH ;
wire  FCA ;
wire  FCB ;
wire  FCC ;
wire  FCD ;
wire  FCE ;
wire  FCF ;
wire  FCG ;
wire  FCH ;
wire  fda ;
wire  FDA ;
wire  fdb ;
wire  FDB ;
wire  fdc ;
wire  FDC ;
wire  fdd ;
wire  FDD ;
wire  fde ;
wire  FDE ;
wire  fdf ;
wire  FDF ;
wire  fdg ;
wire  FDG ;
wire  fdh ;
wire  FDH ;
wire  fdi ;
wire  FDI ;
wire  fdj ;
wire  FDJ ;
wire  fdk ;
wire  FDK ;
wire  fdl ;
wire  FDL ;
wire  fdm ;
wire  FDM ;
wire  fdn ;
wire  FDN ;
wire  fdo ;
wire  FDO ;
wire  fdp ;
wire  FDP ;
wire  fdq ;
wire  FDQ ;
wire  fdr ;
wire  FDR ;
wire  fds ;
wire  FDS ;
wire  fdt ;
wire  FDT ;
wire  fdu ;
wire  FDU ;
wire  fdv ;
wire  FDV ;
wire  fdw ;
wire  FDW ;
wire  fdx ;
wire  FDX ;
wire  fdy ;
wire  FDY ;
wire  fdz ;
wire  FDZ ;
wire  fea ;
wire  FEA ;
wire  gaa ;
wire  gab ;
wire  gac ;
wire  gad ;
wire  gae ;
wire  gaf ;
wire  gag ;
wire  gah ;
wire  gba ;
wire  gbb ;
wire  gbc ;
wire  gbd ;
wire  gbe ;
wire  gbf ;
wire  gbg ;
wire  gbh ;
wire  gca ;
wire  gcb ;
wire  gcc ;
wire  gcd ;
wire  gce ;
wire  gcf ;
wire  gcg ;
wire  gch ;
wire  gda ;
wire  gdb ;
wire  gdc ;
wire  gdd ;
wire  gde ;
wire  gdf ;
wire  gdg ;
wire  gdh ;
wire  gea ;
wire  geb ;
wire  gec ;
wire  ged ;
wire  gee ;
wire  gef ;
wire  geg ;
wire  gfa ;
wire  gfb ;
wire  gfc ;
wire  gfd ;
wire  gfe ;
wire  gff ;
wire  gfi ;
wire  gga ;
wire  ggb ;
wire  ggc ;
wire  ggd ;
wire  gge ;
wire  ggf ;
wire  ggg ;
wire  ggh ;
wire  gha ;
wire  ghb ;
wire  ghc ;
wire  ghd ;
wire  ghe ;
wire  ghf ;
wire  ghg ;
wire  ghh ;
wire  gia ;
wire  gib ;
wire  gic ;
wire  gid ;
wire  gie ;
wire  gif ;
wire  gig ;
wire  gih ;
wire  gja ;
wire  gjb ;
wire  gjc ;
wire  gjd ;
wire  gje ;
wire  gjf ;
wire  gjg ;
wire  gjh ;
wire  gka ;
wire  gkb ;
wire  gkc ;
wire  gkd ;
wire  gke ;
wire  gkf ;
wire  gkg ;
wire  gla ;
wire  glb ;
wire  glc ;
wire  gld ;
wire  gle ;
wire  glf ;
wire  glg ;
wire  glh ;
wire  GQA ;
wire  GQB ;
wire  GQC ;
wire  GQD ;
wire  GQE ;
wire  GQF ;
wire  GQG ;
wire  GQH ;
wire  GQI ;
wire  GQJ ;
wire  GQK ;
wire  GQL ;
wire  GQM ;
wire  GQN ;
wire  GQO ;
wire  GQP ;
wire  haa ;
wire  hab ;
wire  hac ;
wire  had ;
wire  hae ;
wire  haf ;
wire  hag ;
wire  hah ;
wire  hba ;
wire  hbb ;
wire  hbc ;
wire  hbd ;
wire  hbe ;
wire  hbf ;
wire  hbg ;
wire  hbh ;
wire  hca ;
wire  hcb ;
wire  hcc ;
wire  hcd ;
wire  hce ;
wire  hcf ;
wire  hcg ;
wire  hch ;
wire  hda ;
wire  hdb ;
wire  hdc ;
wire  hdd ;
wire  hde ;
wire  hdf ;
wire  hdg ;
wire  hdh ;
wire  HEA ;
wire  HEB ;
wire  HEC ;
wire  HED ;
wire  HEE ;
wire  HEF ;
wire  hfa ;
wire  hfb ;
wire  hfc ;
wire  hfd ;
wire  hfe ;
wire  hff ;
wire  hfg ;
wire  hfh ;
wire  hfi ;
wire  iaa ;
wire  iab ;
wire  iac ;
wire  iad ;
wire  iae ;
wire  iaf ;
wire  iag ;
wire  iah ;
wire  iai ;
wire  iaj ;
wire  iak ;
wire  ial ;
wire  iam ;
wire  ian ;
wire  iao ;
wire  iap ;
wire  iba ;
wire  ibb ;
wire  ibc ;
wire  ibd ;
wire  ibe ;
wire  ibf ;
wire  ibg ;
wire  ibh ;
wire  ibi ;
wire  ibj ;
wire  ibk ;
wire  ibl ;
wire  ibm ;
wire  ibn ;
wire  ibo ;
wire  ibp ;
wire  ica ;
wire  icb ;
wire  icc ;
wire  icd ;
wire  ice ;
wire  icf ;
wire  icg ;
wire  ich ;
wire  ici ;
wire  icj ;
wire  ick ;
wire  icl ;
wire  icm ;
wire  icn ;
wire  ico ;
wire  icp ;
wire  ida ;
wire  idb ;
wire  idc ;
wire  idd ;
wire  ide ;
wire  idf ;
wire  idg ;
wire  idh ;
wire  idi ;
wire  idj ;
wire  idk ;
wire  idl ;
wire  idm ;
wire  idn ;
wire  ido ;
wire  idp ;
wire  iea ;
wire  ieb ;
wire  iec ;
wire  ied ;
wire  iee ;
wire  ief ;
wire  ieg ;
wire  ieh ;
wire  ifa ;
wire  ifb ;
wire  ifc ;
wire  ifd ;
wire  iga ;
wire  igb ;
wire  ija ;
wire  ijb ;
wire  ijc ;
wire  ijd ;
wire  ije ;
wire  ijj ;
wire  ijk ;
wire  ika ;
wire  ikb ;
wire  ikc ;
wire  ikq ;
wire  ila ;
wire  izz ;
wire  jaa ;
wire  JAA ;
wire  jab ;
wire  JAB ;
wire  jac ;
wire  JAC ;
wire  jad ;
wire  JAD ;
wire  jae ;
wire  JAE ;
wire  jaf ;
wire  JAF ;
wire  jag ;
wire  JAG ;
wire  jah ;
wire  JAH ;
wire  jba ;
wire  JBA ;
wire  jbb ;
wire  JBB ;
wire  jbc ;
wire  JBC ;
wire  jbd ;
wire  JBD ;
wire  jbe ;
wire  JBE ;
wire  JCA ;
wire  JCB ;
wire  JCC ;
wire  JCD ;
wire  JCE ;
wire  JCF ;
wire  JCG ;
wire  JCH ;
wire  jda ;
wire  JDA ;
wire  jdb ;
wire  JDB ;
wire  jdc ;
wire  JDC ;
wire  jdi ;
wire  JDI ;
wire  jfa ;
wire  JFA ;
wire  jfb ;
wire  JFB ;
wire  jfc ;
wire  JFC ;
wire  jfd ;
wire  JFD ;
wire  jfi ;
wire  JFI ;
wire  jga ;
wire  JGA ;
wire  jgb ;
wire  JGB ;
wire  jgc ;
wire  JGC ;
wire  jgd ;
wire  JGD ;
wire  jge ;
wire  JGE ;
wire  jgf ;
wire  JGF ;
wire  jgg ;
wire  JGG ;
wire  jgi ;
wire  JGI ;
wire  jka ;
wire  JKA ;
wire  jkb ;
wire  JKB ;
wire  jkc ;
wire  JKC ;
wire  jkd ;
wire  JKD ;
wire  jke ;
wire  JKE ;
wire  jkf ;
wire  JKF ;
wire  jkg ;
wire  JKG ;
wire  jkh ;
wire  JKH ;
wire  jki ;
wire  JKI ;
wire  jla ;
wire  JLA ;
wire  jlb ;
wire  JLB ;
wire  jlc ;
wire  JLC ;
wire  jld ;
wire  JLD ;
wire  jle ;
wire  JLE ;
wire  jlf ;
wire  JLF ;
wire  jlg ;
wire  JLG ;
wire  jma ;
wire  JMA ;
wire  jmb ;
wire  JMB ;
wire  jmc ;
wire  JMC ;
wire  jmd ;
wire  JMD ;
wire  jme ;
wire  JME ;
wire  jmf ;
wire  JMF ;
wire  jna ;
wire  JNA ;
wire  jnb ;
wire  JNB ;
wire  joa ;
wire  JOA ;
wire  job ;
wire  JOB ;
wire  joc ;
wire  JOC ;
wire  jpa ;
wire  JPA ;
wire  jwa ;
wire  JWA ;
wire  jwb ;
wire  JWB ;
wire  jwc ;
wire  JWC ;
wire  jwd ;
wire  JWD ;
wire  jwe ;
wire  JWE ;
wire  jwf ;
wire  JWF ;
wire  jwg ;
wire  JWG ;
wire  jwh ;
wire  JWH ;
wire  jxa ;
wire  JXA ;
wire  kaa ;
wire  kab ;
wire  kac ;
wire  kad ;
wire  kaf ;
wire  kag ;
wire  kba ;
wire  kbb ;
wire  kbc ;
wire  kbd ;
wire  kbf ;
wire  kbg ;
wire  kca ;
wire  kcb ;
wire  kcc ;
wire  kcd ;
wire  kcf ;
wire  kcg ;
wire  kda ;
wire  kdb ;
wire  kdc ;
wire  kdd ;
wire  kdf ;
wire  kdg ;
wire  kea ;
wire  keb ;
wire  kec ;
wire  ked ;
wire  kef ;
wire  keg ;
wire  kfa ;
wire  kfb ;
wire  kfc ;
wire  kfd ;
wire  kfe ;
wire  kff ;
wire  kfg ;
wire  kga ;
wire  kgb ;
wire  kgc ;
wire  kgd ;
wire  kge ;
wire  kgf ;
wire  kgg ;
wire  kha ;
wire  khb ;
wire  khc ;
wire  khd ;
wire  khe ;
wire  khf ;
wire  khg ;
wire  kia ;
wire  kib ;
wire  kic ;
wire  kid ;
wire  kie ;
wire  kif ;
wire  kig ;
wire  kja ;
wire  kjb ;
wire  kjc ;
wire  kjd ;
wire  kje ;
wire  kjf ;
wire  kjg ;
wire  kka ;
wire  kkb ;
wire  kkc ;
wire  kkd ;
wire  kke ;
wire  kkf ;
wire  kla ;
wire  klb ;
wire  klc ;
wire  kld ;
wire  kle ;
wire  klf ;
wire  laa ;
wire  lab ;
wire  lac ;
wire  lba ;
wire  lbb ;
wire  lbc ;
wire  LBG ;
wire  lca ;
wire  lcb ;
wire  lcc ;
wire  lcd ;
wire  lce ;
wire  lcf ;
wire  lcg ;
wire  lda ;
wire  ldb ;
wire  ldc ;
wire  ldd ;
wire  lde ;
wire  ldf ;
wire  ldg ;
wire  lea ;
wire  leb ;
wire  lec ;
wire  led ;
wire  lee ;
wire  lef ;
wire  leg ;
wire  lfa ;
wire  lfb ;
wire  lfc ;
wire  lfd ;
wire  lfe ;
wire  lff ;
wire  lfg ;
wire  lga ;
wire  lgb ;
wire  lgc ;
wire  lgd ;
wire  lge ;
wire  lgf ;
wire  lgg ;
wire  lha ;
wire  lhb ;
wire  lhc ;
wire  lhd ;
wire  lhe ;
wire  lhf ;
wire  lhg ;
wire  lia ;
wire  lib ;
wire  lic ;
wire  lid ;
wire  lie ;
wire  lif ;
wire  lig ;
wire  lja ;
wire  ljb ;
wire  ljc ;
wire  ljd ;
wire  lje ;
wire  ljf ;
wire  ljg ;
wire  lka ;
wire  lkb ;
wire  lkc ;
wire  lkd ;
wire  lke ;
wire  lkf ;
wire  lkg ;
wire  lla ;
wire  llb ;
wire  llc ;
wire  lld ;
wire  lle ;
wire  llf ;
wire  llg ;
wire  lma ;
wire  lmb ;
wire  lmc ;
wire  lmd ;
wire  lme ;
wire  lmf ;
wire  lmg ;
wire  lna ;
wire  lnb ;
wire  lnc ;
wire  lnd ;
wire  lne ;
wire  lnf ;
wire  lng ;
wire  loa ;
wire  lob ;
wire  loc ;
wire  lod ;
wire  loe ;
wire  lof ;
wire  log ;
wire  lpa ;
wire  lpb ;
wire  lpc ;
wire  lpd ;
wire  lpe ;
wire  lpf ;
wire  lpg ;
wire  lqa ;
wire  lqb ;
wire  lqc ;
wire  lqd ;
wire  lqe ;
wire  lqf ;
wire  lqg ;
wire  lra ;
wire  lrb ;
wire  lrc ;
wire  lrd ;
wire  lre ;
wire  lrf ;
wire  lsa ;
wire  lsb ;
wire  lsc ;
wire  lsd ;
wire  lse ;
wire  lsf ;
wire  maa ;
wire  MAA ;
wire  mab ;
wire  MAB ;
wire  mac ;
wire  MAC ;
wire  mad ;
wire  MAD ;
wire  mae ;
wire  MAE ;
wire  maf ;
wire  MAF ;
wire  mag ;
wire  MAG ;
wire  mah ;
wire  MAH ;
wire  mba ;
wire  MBA ;
wire  mbb ;
wire  MBB ;
wire  mbc ;
wire  MBC ;
wire  mbd ;
wire  MBD ;
wire  mbe ;
wire  MBE ;
wire  mbf ;
wire  MBF ;
wire  mbg ;
wire  MBG ;
wire  mbh ;
wire  MBH ;
wire  NAA ;
wire  NAB ;
wire  NAC ;
wire  NAD ;
wire  nag ;
wire  NCA ;
wire  NCB ;
wire  NCC ;
wire  NCD ;
wire  NCE ;
wire  NCF ;
wire  NCG ;
wire  NCH ;
wire  NDA ;
wire  NDB ;
wire  NDC ;
wire  NDD ;
wire  NDE ;
wire  NDF ;
wire  NDG ;
wire  NDH ;
wire  NDI ;
wire  NDJ ;
wire  NDK ;
wire  NDL ;
wire  NEA ;
wire  NEB ;
wire  NEC ;
wire  NEE ;
wire  NEI ;
wire  NIA ;
wire  NIB ;
wire  NIC ;
wire  nka ;
wire  nkb ;
wire  nkc ;
wire  nkd ;
wire  nke ;
wire  nkf ;
wire  nkg ;
wire  nkh ;
wire  nki ;
wire  nkj ;
wire  nkk ;
wire  nkl ;
wire  nkm ;
wire  nkn ;
wire  nko ;
wire  nkp ;
wire  nkq ;
wire  nkr ;
wire  nks ;
wire  nkt ;
wire  NKU ;
wire  nla ;
wire  nlb ;
wire  nlc ;
wire  nld ;
wire  nle ;
wire  nlf ;
wire  nlg ;
wire  nlh ;
wire  OAA ;
wire  OAB ;
wire  OAC ;
wire  OAD ;
wire  OAE ;
wire  OAF ;
wire  OAG ;
wire  OAH ;
wire  OAI ;
wire  OAJ ;
wire  OAK ;
wire  OAL ;
wire  OAM ;
wire  OAN ;
wire  OAO ;
wire  OAP ;
wire  OBA ;
wire  OBB ;
wire  OBC ;
wire  OBD ;
wire  OBE ;
wire  OBF ;
wire  OBG ;
wire  OBH ;
wire  OBI ;
wire  OBJ ;
wire  OBK ;
wire  OBL ;
wire  OBM ;
wire  OBN ;
wire  OBO ;
wire  OBP ;
wire  OCA ;
wire  OCB ;
wire  OCC ;
wire  OCD ;
wire  OCE ;
wire  OCF ;
wire  OCG ;
wire  OCH ;
wire  OCI ;
wire  OCJ ;
wire  OCK ;
wire  OCL ;
wire  OCM ;
wire  OCN ;
wire  OCO ;
wire  OCP ;
wire  ODA ;
wire  ODB ;
wire  ODC ;
wire  ODD ;
wire  ODE ;
wire  ODF ;
wire  ODG ;
wire  ODH ;
wire  ODI ;
wire  ODJ ;
wire  oea ;
wire  oeb ;
wire  oec ;
wire  oed ;
wire  oee ;
wire  oef ;
wire  ofa ;
wire  ofb ;
wire  ofc ;
wire  ofd ;
wire  ofe ;
wire  off ;
wire  oga ;
wire  ogb ;
wire  ogc ;
wire  oha ;
wire  ohb ;
wire  ohc ;
wire  ohd ;
wire  ohe ;
wire  ohf ;
wire  ohg ;
wire  oia ;
wire  oib ;
wire  OJA ;
wire  OJB ;
wire  OJC ;
wire  ojd ;
wire  OKA ;
wire  OLA ;
wire  OLB ;
wire  OLC ;
wire  OLD ;
wire  OLE ;
wire  OLF ;
wire  OLG ;
wire  OLH ;
wire  oma ;
wire  omb ;
wire  ONA ;
wire  ONB ;
wire  ooa ;
wire  oob ;
wire  ooc ;
wire  ood ;
wire  ooe ;
wire  oof ;
wire  OPA ;
wire  opb ;
wire  opc ;
wire  OPD ;
wire  OQA ;
wire  oqb ;
wire  oqc ;
wire  ORA ;
wire  orb ;
wire  orc ;
wire  ord ;
wire  OSA ;
wire  osb ;
wire  osc ;
wire  osd ;
wire  OSE ;
wire  OTA ;
wire  OTB ;
wire  otc ;
wire  OTD ;
wire  ote ;
wire  otf ;
wire  otg ;
wire  OUA ;
wire  OUB ;
wire  ouc ;
wire  oud ;
wire  oue ;
wire  OVA ;
wire  ovb ;
wire  ovc ;
wire  ovd ;
wire  ove ;
wire  ovf ;
wire  owa ;
wire  owb ;
wire  owc ;
wire  owd ;
wire  owe ;
wire  owf ;
wire  OWG ;
wire  OWH ;
wire  OWI ;
wire  OWJ ;
wire  OWK ;
wire  OWL ;
wire  owm ;
wire  own ;
wire  owo ;
wire  OWP ;
wire  owq ;
wire  OWR ;
wire  ows ;
wire  owt ;
wire  OWU ;
wire  OWV ;
wire  OWW ;
wire  OWX ;
wire  oxa ;
wire  oxb ;
wire  oxc ;
wire  OZA ;
wire  OZB ;
wire  paa ;
wire  pab ;
wire  pac ;
wire  pad ;
wire  pae ;
wire  paf ;
wire  pag ;
wire  pah ;
wire  pba ;
wire  pbb ;
wire  pbc ;
wire  pbd ;
wire  pbe ;
wire  pbf ;
wire  pbg ;
wire  pbh ;
wire  pca ;
wire  pcb ;
wire  pcc ;
wire  pcd ;
wire  pce ;
wire  pcf ;
wire  pcg ;
wire  pda ;
wire  pdb ;
wire  pdc ;
wire  pdd ;
wire  pde ;
wire  pdf ;
wire  pdg ;
wire  pdh ;
wire  pea ;
wire  peb ;
wire  pec ;
wire  ped ;
wire  pee ;
wire  pef ;
wire  pfa ;
wire  pfb ;
wire  pfc ;
wire  pfd ;
wire  pfe ;
wire  pff ;
wire  pfg ;
wire  pfh ;
wire  pga ;
wire  pgb ;
wire  pgc ;
wire  pgd ;
wire  pge ;
wire  pgf ;
wire  pgg ;
wire  pha ;
wire  phb ;
wire  phc ;
wire  phd ;
wire  phe ;
wire  phf ;
wire  phg ;
wire  phh ;
wire  pia ;
wire  pib ;
wire  pic ;
wire  pid ;
wire  pie ;
wire  pja ;
wire  pjc ;
wire  pjd ;
wire  pje ;
wire  pjf ;
wire  pka ;
wire  pkb ;
wire  pkc ;
wire  pkd ;
wire  pke ;
wire  pkf ;
wire  pla ;
wire  plb ;
wire  plc ;
wire  pld ;
wire  ple ;
wire  plf ;
wire  pma ;
wire  pmb ;
wire  pmc ;
wire  pmd ;
wire  pme ;
wire  pmf ;
wire  pna ;
wire  pnb ;
wire  pnc ;
wire  pnd ;
wire  pne ;
wire  pnf ;
wire  poa ;
wire  pob ;
wire  poc ;
wire  pod ;
wire  poe ;
wire  pof ;
wire  QAA ;
wire  QAB ;
wire  QAC ;
wire  QAD ;
wire  QAE ;
wire  QAF ;
wire  QAG ;
wire  QAH ;
wire  QBA ;
wire  QBB ;
wire  QBC ;
wire  QBD ;
wire  QBE ;
wire  QBF ;
wire  QBG ;
wire  QBH ;
wire  qca ;
wire  qcb ;
wire  qcc ;
wire  qcd ;
wire  qce ;
wire  QDA ;
wire  QDB ;
wire  QDC ;
wire  QDD ;
wire  QEA ;
wire  QEB ;
wire  QEC ;
wire  QED ;
wire  QEE ;
wire  QFA ;
wire  QFB ;
wire  QFC ;
wire  QFD ;
wire  QFE ;
wire  QFF ;
wire  qga ;
wire  qgb ;
wire  qgc ;
wire  QGD ;
wire  QGE ;
wire  qha ;
wire  qhb ;
wire  qhd ;
wire  qhf ;
wire  qhg ;
wire  qhi ;
wire  qhj ;
wire  qhk ;
wire  qhl ;
wire  qia ;
wire  qib ;
wire  qic ;
wire  qid ;
wire  QIE ;
wire  qja ;
wire  QKA ;
wire  QKB ;
wire  qla ;
wire  qlb ;
wire  qlc ;
wire  qma ;
wire  qmb ;
wire  qmc ;
wire  qmd ;
wire  raa ;
wire  rab ;
wire  rac ;
wire  rad ;
wire  rae ;
wire  raf ;
wire  rag ;
wire  rah ;
wire  rai ;
wire  raj ;
wire  rak ;
wire  ral ;
wire  ram ;
wire  ran ;
wire  rao ;
wire  rap ;
wire  raq ;
wire  rar ;
wire  ras ;
wire  rat ;
wire  rau ;
wire  rav ;
wire  raw ;
wire  rax ;
wire  tca ;
wire  TCA ;
wire  tcb ;
wire  TCB ;
wire  tcc ;
wire  TCC ;
wire  tcd ;
wire  TCD ;
wire  tce ;
wire  TCE ;
wire  tcf ;
wire  TCF ;
wire  tcg ;
wire  TCG ;
wire  tch ;
wire  TCH ;
wire  tci ;
wire  TCI ;
wire  tcj ;
wire  TCJ ;
wire  tck ;
wire  TCK ;
wire  tcl ;
wire  TCL ;
wire  tcm ;
wire  TCM ;
wire  tcn ;
wire  TCN ;
wire  tco ;
wire  TCO ;
wire  tcp ;
wire  TCP ;
wire  tcq ;
wire  TCQ ;
wire  tcr ;
wire  TCR ;
wire  tcs ;
wire  TCS ;
wire  tct ;
wire  TCT ;
wire  tcu ;
wire  TCU ;
wire  tcv ;
wire  TCV ;
wire  tcw ;
wire  TCW ;
wire  tcx ;
wire  TCX ;
wire  tea ;
wire  TEA ;
wire  teb ;
wire  TEB ;
wire  tec ;
wire  TEC ;
wire  ted ;
wire  TED ;
wire  tee ;
wire  TEE ;
wire  tef ;
wire  TEF ;
wire  teg ;
wire  TEG ;
wire  teh ;
wire  TEH ;
wire  tei ;
wire  TEI ;
wire  tej ;
wire  TEJ ;
wire  tek ;
wire  TEK ;
wire  tel ;
wire  TEL ;
wire  tem ;
wire  TEM ;
wire  ten ;
wire  TEN ;
wire  teo ;
wire  TEO ;
wire  tep ;
wire  TEP ;
wire  teq ;
wire  TEQ ;
wire  tes ;
wire  TES ;
wire  tga ;
wire  TGA ;
wire  tgb ;
wire  TGB ;
wire  tgc ;
wire  TGC ;
wire  tgd ;
wire  TGD ;
wire  tge ;
wire  TGE ;
wire  tgf ;
wire  TGF ;
wire  tgg ;
wire  TGG ;
wire  tgh ;
wire  TGH ;
wire  tgi ;
wire  TGI ;
wire  tgq ;
wire  TGQ ;
wire  tgr ;
wire  TGR ;
wire  tgs ;
wire  TGS ;
wire  tgt ;
wire  TGT ;
wire  tha ;
wire  THA ;
wire  thb ;
wire  THB ;
wire  thc ;
wire  THC ;
wire  thd ;
wire  THD ;
wire  the ;
wire  THE ;
wire  thf ;
wire  THF ;
wire  thg ;
wire  THG ;
wire  thh ;
wire  THH ;
wire  thi ;
wire  THI ;
wire  thj ;
wire  THJ ;
wire  thk ;
wire  THK ;
wire  thl ;
wire  THL ;
wire  thm ;
wire  THM ;
wire  tia ;
wire  TIA ;
wire  tib ;
wire  TIB ;
wire  tic ;
wire  TIC ;
wire  tid ;
wire  TID ;
wire  tie ;
wire  TIE ;
wire  tif ;
wire  TIF ;
wire  tig ;
wire  TIG ;
wire  tii ;
wire  TII ;
wire  tij ;
wire  TIJ ;
wire  tja ;
wire  TJA ;
wire  tjb ;
wire  TJB ;
wire  tjc ;
wire  TJC ;
wire  tjd ;
wire  TJD ;
wire  tje ;
wire  TJE ;
wire  tjf ;
wire  TJF ;
wire  tjg ;
wire  TJG ;
wire  tjh ;
wire  TJH ;
wire  tji ;
wire  TJI ;
wire  tjj ;
wire  TJJ ;
wire  tjk ;
wire  TJK ;
wire  tjl ;
wire  TJL ;
wire  tjm ;
wire  TJM ;
wire  tjn ;
wire  TJN ;
wire  tjo ;
wire  TJO ;
wire  tjp ;
wire  TJP ;
wire  tjq ;
wire  TJQ ;
wire  tjr ;
wire  TJR ;
wire  tjs ;
wire  TJS ;
wire  tjt ;
wire  TJT ;
wire  waa ;
wire  wab ;
wire  wac ;
wire  wad ;
wire  wae ;
wire  waf ;
wire  wag ;
wire  wah ;
wire  wba ;
wire  wbb ;
wire  wbc ;
wire  wbd ;
wire  wbe ;
wire  wbf ;
wire  wbg ;
wire  wbh ;
wire  wca ;
wire  wcb ;
wire  wcc ;
wire  wda ;
wire  wdb ;
wire  wdc ;
wire  yyy ;
wire  YYY ;
wire  ZZI ;
wire  ZZO ;
assign ZZI = 1'b1;
assign ZZO = 1'b0;
assign yyy =  ZZO  ; 
assign YYY = ~yyy;  //complement 
assign pia = ~PIA;  //complement 
assign pib = ~PIB;  //complement 
assign pic = ~PIC;  //complement 
assign pea = ~PEA;  //complement 
assign peb = ~PEB;  //complement 
assign pec = ~PEC;  //complement 
assign paa = ~PAA;  //complement 
assign pab = ~PAB;  //complement 
assign pac = ~PAC;  //complement 
assign DAA =  PAA & PHA & pna  ; 
assign daa = ~DAA;  //complement 
assign DAI =  PCA & PHA & PJA  ; 
assign dai = ~DAI;  //complement 
assign DAQ =  PAA & PJA  ; 
assign daq = ~DAQ;  //complement 
assign DBA =  PDA & PGA & pna  ; 
assign dba = ~DBA;  //complement 
assign DBI =  PDA & PEA  ; 
assign dbi = ~DBI;  //complement 
assign DBQ =  PAA & PGA  ; 
assign dbq = ~DBQ;  //complement 
assign DCA =  pba & paa  ; 
assign dca = ~DCA;  //complement 
assign DCI =  PDA & PGA & PKA  ; 
assign dci = ~DCI;  //complement 
assign DCQ =  PBA & pea & PKA  ; 
assign dcq = ~DCQ;  //complement 
assign ped = ~PED;  //complement 
assign pee = ~PEE;  //complement 
assign DDA =  PAA & PEA & PJA & pma  ; 
assign dda = ~DDA;  //complement  
assign DDI =  PBA & PEA & PNA & PMB  ; 
assign ddi = ~DDI;  //complement 
assign DEA =  PAA & PHA & PKA & pma  ; 
assign dea = ~DEA;  //complement  
assign DEI =  PBA & poa & PKA & pma  ; 
assign dei = ~DEI;  //complement 
assign CQA = ~cqa;  //complement 
assign CQI = ~cqi;  //complement 
assign eca = ~ECA;  //complement 
assign eci = ~ECI;  //complement 
assign eda = ~EDA;  //complement 
assign edi = ~EDI;  //complement 
assign teq =  WAA & QFB  |  WBA & QFC  ; 
assign TEQ = ~teq;  //complement 
assign tea =  WAA & QFB  |  WBA & QFC  ; 
assign TEA = ~tea; //complement 
assign tei =  WAA & QFB  |  WBA & QFC  ; 
assign TEI = ~tei;  //complement 
assign eba = ~EBA;  //complement 
assign ebi = ~EBI;  //complement 
assign eaa = ~EAA;  //complement 
assign eai = ~EAI;  //complement 
assign thi =  WAB  |  WBB  ; 
assign THI = ~thi;  //complement 
assign thb =  WAB  |  WBB  ; 
assign THB = ~thb; //complement 
assign tha =  WAB  |  WBB  ; 
assign THA = ~tha;  //complement 
assign eea = ~EEA;  //complement 
assign eei = ~EEI;  //complement 
assign eqa = ~EQA;  //complement 
assign eqi = ~EQI;  //complement 
assign FCA = ~EQC & ~EQB & ~EQA  ; 
assign FCB = ~EQC & ~EQB &  EQA  ; 
assign FCC = ~EQC &  EQB & ~EQA  ; 
assign FCD = ~EQC &  EQB &  EQA  ; 
assign FCE =  EQC & ~EQB & ~EQA  ; 
assign FCF =  EQC & ~EQB &  EQA ; 
assign FCG =  EQC &  EQB & ~EQA  ; 
assign FCH =  EQC &  EQB &  EQA ; 
assign gla = ~GLA;  //complement 
assign fdb =  eba & edi & ebg & ebj & ebe  ; 
assign FDB = ~fdb;  //complement  
assign fdj =  eca & ecl & eda & eci  ; 
assign FDJ = ~fdj;  //complement 
assign fdn =  eca & eda  ; 
assign FDN = ~fdn;  //complement  
assign fdy =  ebe & eba  ; 
assign FDY = ~fdy;  //complement 
assign FDZ =  EDO & eea  ; 
assign fdz = ~FDZ;  //complement  
assign BAA =  AAI & RAA  |  ABI & RAB  |  ACI & RAC  |  ADI & RAD  ; 
assign baa = ~BAA;  //complement 
assign BBA =  AAI & RAA  |  ABI & RAB  |  ACI & RAC  |  ADI & RAD  ; 
assign bba = ~BBA; //complement 
assign BCA =  AAI & RAA  |  ABI & RAB  |  ACI & RAC  |  ADI & RAD  ; 
assign bca = ~BCA;  //complement 
assign aaa = ~AAA;  //complement 
assign aai = ~AAI;  //complement 
assign aba = ~ABA;  //complement 
assign abi = ~ABI;  //complement 
assign BDA =  AAA & RAI  |  ABA & RAJ  |  ACA & RAK  |  ADA & RAL  ; 
assign bda = ~BDA;  //complement 
assign aca = ~ACA;  //complement 
assign aci = ~ACI;  //complement 
assign ada = ~ADA;  //complement 
assign adi = ~ADI;  //complement 
assign raa = ~RAA;  //complement 
assign rai = ~RAI;  //complement 
assign raq = ~RAQ;  //complement 
assign JAA =  rai & raj & rak & ral & QCB  ; 
assign jaa = ~JAA;  //complement  
assign JBA =  RAQ & qce  ; 
assign jba = ~JBA;  //complement 
assign JAH =  rai & raj & rak & ral & QCB  ; 
assign jah = ~JAH;  //complement  
assign TCA =  wac & wbc  |  ZZO  |  ZZI & qeb  |  ZZI & qfc  ; 
assign tca = ~TCA;  //complement 
assign TCI =  wac & wbc  |  ZZO  |  ZZI & qeb  |  ZZI & qfc  ; 
assign tci = ~TCI; //complement 
assign TCQ =  wac & wbc  |  ZZO  |  ZZI & qeb  |  ZZI & qfc  ; 
assign tcq = ~TCQ;  //complement 
assign MBA =  GAA & HAA  |  GBA & HBA  |  GCA & HCA  |  GDA & HDA  |  GEA & HEA  |  GFA & HFA  ;
assign mba = ~MBA;  //complement 
assign ODA = ~oda;  //complement 
assign ODB = ~odb;  //complement 
assign tja =  ZZO  |  ZZO  |  ZZI & WCA  |  ZZI & WDA  ; 
assign TJA = ~tja;  //complement 
assign tji =  ZZO  |  ZZO  |  ZZI & WCA  |  ZZI & WDA  ; 
assign TJI = ~tji; //complement 
assign tjq =  ZZO  |  ZZO  |  ZZI & WCA  |  ZZI & WDA  ; 
assign TJQ = ~tjq;  //complement 
assign TGI =  waa & wba & eai  ; 
assign tgi = ~TGI;  //complement  
assign TGA =  waa & wba & eaa  ; 
assign tga = ~TGA;  //complement 
assign MAA =  GAA & HAA  |  GBA & HBA  |  GCA & HCA  |  GDA & HDA  |  GEA & HEA  |  GFA & HFA  ;
assign maa = ~MAA;  //complement 
assign waa = ~WAA;  //complement 
assign wab = ~WAB;  //complement 
assign TGQ =  waf & wbf  ; 
assign tgq = ~TGQ;  //complement  
assign TIA =  wca & wda & NAA  ; 
assign tia = ~TIA;  //complement 
assign gaa = ~GAA;  //complement 
assign gda = ~GDA;  //complement 
assign gea = ~GEA;  //complement 
assign gha = ~GHA;  //complement 
assign gia = ~GIA;  //complement 
assign gba = ~GBA;  //complement 
assign gfa = ~GFA;  //complement 
assign gga = ~GGA;  //complement 
assign gja = ~GJA;  //complement 
assign gka = ~GKA;  //complement 
assign gca = ~GCA;  //complement 
assign lca = ~LCA;  //complement 
assign lfa = ~LFA;  //complement 
assign lma = ~LMA;  //complement 
assign lna = ~LNA;  //complement 
assign nla = ~NLA;  //complement 
assign nlb = ~NLB;  //complement 
assign nlc = ~NLC;  //complement 
assign nld = ~NLD;  //complement 
assign QAA = ~qaa;  //complement 
assign QBA = ~qba;  //complement 
assign kba = ~KBA;  //complement 
assign kca = ~KCA;  //complement 
assign kda = ~KDA;  //complement 
assign kea = ~KEA;  //complement 
assign OAA = ~oaa;  //complement 
assign OBA = ~oba;  //complement 
assign OCA = ~oca;  //complement 
assign owa = ~OWA;  //complement 
assign jgf =  gee  ; 
assign JGF = ~jgf;  //complement 
assign kaa = ~KAA;  //complement 
assign kfa = ~KFA;  //complement 
assign lqa = ~LQA;  //complement 
assign lra = ~LRA;  //complement 
assign OAI = ~oai;  //complement 
assign OBI = ~obi;  //complement 
assign OCI = ~oci;  //complement 
assign ofa = ~OFA;  //complement 
assign GQA = ~gqa;  //complement 
assign GQI = ~gqi;  //complement 
assign kia = ~KIA;  //complement 
assign kja = ~KJA;  //complement 
assign kla = ~KLA;  //complement 
assign lsa = ~LSA;  //complement 
assign kga = ~KGA;  //complement 
assign kha = ~KHA;  //complement 
assign kka = ~KKA;  //complement 
assign oea = ~OEA;  //complement 
assign haa = ~HAA;  //complement 
assign hba = ~HBA;  //complement 
assign OTD = ~otd;  //complement 
assign QGD = ~qgd;  //complement 
assign oga = ~OGA;  //complement 
assign oha = ~OHA;  //complement 
assign hca = ~HCA;  //complement 
assign hda = ~HDA;  //complement 
assign hfa = ~HFA;  //complement 
assign OTA = ~ota;  //complement 
assign OTB = ~otb;  //complement 
assign OLA = ~ola;  //complement 
assign JCH = ~nic & ~nib & ~nia  ; 
assign JCG = ~nic & ~nib &  nia  ; 
assign JCF = ~nic &  nib & ~nia  ; 
assign JCE = ~nic &  nib &  nia  ; 
assign JCD =  nic & ~nib & ~nia  ; 
assign JCC =  nic & ~nib &  nia ; 
assign JCB =  nic &  nib & ~nia  ; 
assign JCA =  nic &  nib &  nia ; 
assign jfa =  nea & neb & nei  ; 
assign JFA = ~jfa;  //complement 
assign jda =  hfa  ; 
assign JDA = ~jda;  //complement 
assign JWA =  qga  ; 
assign jwa = ~JWA;  //complement 
assign qhf = ~QHF;  //complement 
assign qhk = ~QHK;  //complement 
assign HEA = ~hea;  //complement 
assign ooa = ~OOA;  //complement 
assign ood = ~OOD;  //complement 
assign owd = ~OWD;  //complement 
assign NAA = ~naa;  //complement 
assign NIA = ~nia;  //complement 
assign NCA = ~nca;  //complement 
assign NDJ = ~ndj;  //complement 
assign qhj = ~QHJ;  //complement 
assign qhl = ~QHL;  //complement 
assign NDA = ~nda;  //complement 
assign ONA = ~ona;  //complement 
assign OWG = ~owg;  //complement 
assign OPD = ~opd;  //complement 
assign OSE = ~ose;  //complement 
assign NEA = ~nea;  //complement 
assign lba = ~LBA;  //complement 
assign lda = ~LDA;  //complement 
assign lea = ~LEA;  //complement 
assign lga = ~LGA;  //complement 
assign lia = ~LIA;  //complement 
assign lja = ~LJA;  //complement 
assign lka = ~LKA;  //complement 
assign lla = ~LLA;  //complement 
assign loa = ~LOA;  //complement 
assign lpa = ~LPA;  //complement 
assign laa = ~LAA;  //complement 
assign pja = ~PJA;  //complement 
assign pjc = ~PJC;  //complement 
assign pfa = ~PFA;  //complement 
assign pfb = ~PFB;  //complement 
assign pfc = ~PFC;  //complement 
assign pba = ~PBA;  //complement 
assign pbb = ~PBB;  //complement 
assign pbc = ~PBC;  //complement 
assign DAB =  PAB & PGB & pnb  ; 
assign dab = ~DAB;  //complement 
assign DAJ =  PBB & POB & PIB  ; 
assign daj = ~DAJ;  //complement 
assign DAR =  PAB & pob & PIB  ; 
assign dar = ~DAR;  //complement 
assign DBB =  PAB & PGB & PIB  ; 
assign dbb = ~DBB;  //complement 
assign DBJ =  PCB & PEB & PLB  ; 
assign dbj = ~DBJ;  //complement 
assign DCB =  PCB & PFB & pnb  ; 
assign dcb = ~DCB;  //complement 
assign DCJ =  PDB & PFB & pnb  ; 
assign dcj = ~DCJ;  //complement 
assign pfd = ~PFD;  //complement 
assign pfe = ~PFE;  //complement 
assign DDB =  PBB & PEB & PLB & PMD  ; 
assign ddb = ~DDB;  //complement  
assign DDJ =  PDB & PGB & plb  ; 
assign ddj = ~DDJ;  //complement 
assign DEB =  PBB & PEB & PKB & pmb  ; 
assign deb = ~DEB;  //complement  
assign DEJ =  PBB & pob & PNB  ; 
assign dej = ~DEJ;  //complement 
assign DFB =  PBB & PHB & PKB  ; 
assign dfb = ~DFB;  //complement  
assign DFJ =  PAB & PEB & PLB  ; 
assign dfj = ~DFJ;  //complement 
assign CQB = ~cqb;  //complement 
assign CQJ = ~cqj;  //complement 
assign DEN =  PBB & poa & PLA  ; 
assign den = ~DEN;  //complement  
assign ecb = ~ECB;  //complement 
assign ecj = ~ECJ;  //complement 
assign edb = ~EDB;  //complement 
assign edj = ~EDJ;  //complement 
assign teb =  WAA & QFB  |  WBA & QFC  ; 
assign TEB = ~teb; //complement 
assign tej =  WAA & QFB  |  WBA & QFC  ; 
assign TEJ = ~tej;  //complement 
assign ebb = ~EBB;  //complement 
assign ebj = ~EBJ;  //complement 
assign eab = ~EAB;  //complement 
assign thj =  WAB  |  WBB  ; 
assign THJ = ~thj;  //complement 
assign thd =  WAB  |  WBB  ; 
assign THD = ~thd; //complement 
assign thc =  WAB  |  WBB  ; 
assign THC = ~thc;  //complement 
assign EEB = ~eeb;  //complement 
assign eej = ~EEJ;  //complement 
assign eqb = ~EQB;  //complement 
assign eqj = ~EQJ;  //complement 
assign glb = ~GLB;  //complement 
assign fdc =  ebb & ebj  ; 
assign FDC = ~fdc;  //complement  
assign fdk =  ecj & edb & edh  ; 
assign FDK = ~fdk;  //complement 
assign fdr =  eeg & edj  ; 
assign FDR = ~fdr;  //complement  
assign BAB =  AAJ & RAA  |  ABJ & RAB  |  ACJ & RAC  |  ADJ & RAD  ; 
assign bab = ~BAB;  //complement 
assign BBB =  AAJ & RAA  |  ABJ & RAB  |  ACJ & RAC  |  ADJ & RAD  ; 
assign bbb = ~BBB; //complement 
assign BCB =  AAJ & RAA  |  ABJ & RAB  |  ACJ & RAC  |  ADJ & RAD  ; 
assign bcb = ~BCB;  //complement 
assign aab = ~AAB;  //complement 
assign aaj = ~AAJ;  //complement 
assign abb = ~ABB;  //complement 
assign abj = ~ABJ;  //complement 
assign BDB =  AAB & RAI  |  ABB & RAJ  |  ACB & RAK  |  ADB & RAL  ; 
assign bdb = ~BDB;  //complement 
assign acb = ~ACB;  //complement 
assign acj = ~ACJ;  //complement 
assign adb = ~ADB;  //complement 
assign adj = ~ADJ;  //complement 
assign rab = ~RAB;  //complement 
assign raj = ~RAJ;  //complement 
assign rar = ~RAR;  //complement 
assign JAB =  rai & raj & rak & ral & QCB  ; 
assign jab = ~JAB;  //complement  
assign JBB =  RAR & qce  ; 
assign jbb = ~JBB;  //complement 
assign GQB = ~gqb;  //complement 
assign GQJ = ~gqj;  //complement 
assign TCB =  wac & wbc  |  ZZO  |  ZZI & qeb  |  ZZI & qfc  ; 
assign tcb = ~TCB;  //complement 
assign TCJ =  wac & wbc  |  ZZO  |  ZZI & qeb  |  ZZI & qfc  ; 
assign tcj = ~TCJ; //complement 
assign TCR =  wac & wbc  |  ZZO  |  ZZI & qeb  |  ZZI & qfc  ; 
assign tcr = ~TCR;  //complement 
assign MBB =  GAB & HAB  |  GBB & HBB  |  GCB & HCB  |  GDB & HDB  |  GEB & HEB  |  GFB & HFB  ;
assign mbb = ~MBB;  //complement 
assign ODC = ~odc;  //complement 
assign wca = ~WCA;  //complement 
assign tjb =  ZZO  |  ZZO  |  ZZI & WCA  |  ZZI & WDA  ; 
assign TJB = ~tjb;  //complement 
assign tjj =  ZZO  |  ZZO  |  ZZI & WCA  |  ZZI & WDA  ; 
assign TJJ = ~tjj; //complement 
assign tjr =  ZZO  |  ZZO  |  ZZI & WCA  |  ZZI & WDA  ; 
assign TJR = ~tjr;  //complement 
assign TGB =  waa & wba & eab  ; 
assign tgb = ~TGB;  //complement  
assign MAB =  GAB & HAB  |  GBB & HBB  |  GCB & HCB  |  GDB & HDB  |  GEB & HEB  |  GFB & HFB  ;
assign mab = ~MAB;  //complement 
assign wac = ~WAC;  //complement 
assign wad = ~WAD;  //complement 
assign TGR =  waf & wbf  ; 
assign tgr = ~TGR;  //complement  
assign TIB =  wca & wda & NAB  ; 
assign tib = ~TIB;  //complement 
assign gab = ~GAB;  //complement 
assign gdb = ~GDB;  //complement 
assign geb = ~GEB;  //complement 
assign ghb = ~GHB;  //complement 
assign gib = ~GIB;  //complement 
assign gbb = ~GBB;  //complement 
assign gfb = ~GFB;  //complement 
assign ggb = ~GGB;  //complement 
assign gjb = ~GJB;  //complement 
assign gkb = ~GKB;  //complement 
assign gcb = ~GCB;  //complement 
assign lcb = ~LCB;  //complement 
assign lfb = ~LFB;  //complement 
assign lmb = ~LMB;  //complement 
assign lnb = ~LNB;  //complement 
assign nle = ~NLE;  //complement 
assign nlf = ~NLF;  //complement 
assign nlg = ~NLG;  //complement 
assign nlh = ~NLH;  //complement 
assign QAB = ~qab;  //complement 
assign QBB = ~qbb;  //complement 
assign kbb = ~KBB;  //complement 
assign kcb = ~KCB;  //complement 
assign kdb = ~KDB;  //complement 
assign keb = ~KEB;  //complement 
assign OAB = ~oab;  //complement 
assign OBB = ~obb;  //complement 
assign OCB = ~ocb;  //complement 
assign owb = ~OWB;  //complement 
assign jgg =  gef  ; 
assign JGG = ~jgg;  //complement 
assign kab = ~KAB;  //complement 
assign kfb = ~KFB;  //complement 
assign lqb = ~LQB;  //complement 
assign lrb = ~LRB;  //complement 
assign OAJ = ~oaj;  //complement 
assign OBJ = ~obj;  //complement 
assign OCJ = ~ocj;  //complement 
assign ofb = ~OFB;  //complement 
assign JKA = KJA; 
assign jka = ~JKA; //complement 
assign JKB = KJB; 
assign jkb = ~JKB;  //complement 
assign JKC = KJG & kjc ; 
assign jkc = ~JKC ;  //complement 
assign JKD = KJG & KJC; 
assign jkd = ~JKD; 
assign kib = ~KIB;  //complement 
assign kjb = ~KJB;  //complement 
assign klb = ~KLB;  //complement 
assign lsb = ~LSB;  //complement 
assign kgb = ~KGB;  //complement 
assign khb = ~KHB;  //complement 
assign kkb = ~KKB;  //complement 
assign oeb = ~OEB;  //complement 
assign hab = ~HAB;  //complement 
assign hbb = ~HBB;  //complement 
assign qha = ~QHA;  //complement 
assign qhb = ~QHB;  //complement 
assign ogb = ~OGB;  //complement 
assign oob = ~OOB;  //complement 
assign ooe = ~OOE;  //complement 
assign owe = ~OWE;  //complement 
assign hcb = ~HCB;  //complement 
assign hdb = ~HDB;  //complement 
assign HEB = ~heb;  //complement 
assign hfb = ~HFB;  //complement 
assign ORA = ~ora;  //complement 
assign OSA = ~osa;  //complement 
assign OLB = ~olb;  //complement 
assign qhd = ~QHD;  //complement 
assign qhi = ~QHI;  //complement 
assign jfb =  nea  ; 
assign JFB = ~jfb;  //complement 
assign jdb =  hfb  ; 
assign JDB = ~jdb;  //complement 
assign JWB =  qga  ; 
assign jwb = ~JWB;  //complement 
assign jfc =  neb & nei  ; 
assign JFC = ~jfc;  //complement 
assign jfi =  nei  ; 
assign JFI = ~jfi;  //complement 
assign ohb = ~OHB;  //complement 
assign qhg = ~QHG;  //complement 
assign NIB = ~nib;  //complement 
assign NCB = ~ncb;  //complement 
assign NDK = ~ndk;  //complement 
assign NEB = ~neb;  //complement 
assign OZA = ~oza;  //complement 
assign OZB = ~ozb;  //complement 
assign NDB = ~ndb;  //complement 
assign OWH = ~owh;  //complement 
assign oxa = ~OXA;  //complement 
assign oxb = ~OXB;  //complement 
assign lha = ~LHA;  //complement 
assign lhb = ~LHB;  //complement 
assign lbb = ~LBB;  //complement 
assign ldb = ~LDB;  //complement 
assign leb = ~LEB;  //complement 
assign lgb = ~LGB;  //complement 
assign lib = ~LIB;  //complement 
assign ljb = ~LJB;  //complement 
assign lkb = ~LKB;  //complement 
assign llb = ~LLB;  //complement 
assign lob = ~LOB;  //complement 
assign lpb = ~LPB;  //complement 
assign lab = ~LAB;  //complement 
assign poa = ~POA;  //complement 
assign pob = ~POB;  //complement 
assign poc = ~POC;  //complement 
assign pka = ~PKA;  //complement 
assign pkb = ~PKB;  //complement 
assign pkc = ~PKC;  //complement 
assign pga = ~PGA;  //complement 
assign pgb = ~PGB;  //complement 
assign pgc = ~PGC;  //complement 
assign pca = ~PCA;  //complement 
assign pcb = ~PCB;  //complement 
assign pcc = ~PCC;  //complement 
assign DAC =  PBC & poc  ; 
assign dac = ~DAC;  //complement 
assign DAK =  PBC & pob & PLB  ; 
assign dak = ~DAK;  //complement 
assign DAS =  PAC & PEC & PLB  ; 
assign das = ~DAS;  //complement 
assign DBC =  PAC & PGC & PNC  ; 
assign dbc = ~DBC;  //complement 
assign DBK =  PAC & PHC & plc  ; 
assign dbk = ~DBK;  //complement 
assign DBS =  PBC & PGC & plc  ; 
assign dbs = ~DBS;  //complement 
assign DCC =  PCC & PFC & PJC  ; 
assign dcc = ~DCC;  //complement 
assign DCK =  PCC & PHC & PIC  ; 
assign dck = ~DCK;  //complement 
assign pgd = ~PGD;  //complement 
assign pge = ~PGE;  //complement 
assign DDC =  PBC & PEC & PKC & PMD  ; 
assign ddc = ~DDC;  //complement  
assign DDK =  PDC & PFC & pnc  ; 
assign ddk = ~DDK;  //complement 
assign DEC =  PBC & POC & PLC  ; 
assign dec = ~DEC;  //complement  
assign DEK =  PAC & PFC & PNC  ; 
assign dek = ~DEK;  //complement 
assign DFC =  PBC & PFC & PLC & pmc  ; 
assign dfc = ~DFC;  //complement  
assign DFK =  PCC & PGC & pnc  ; 
assign dfk = ~DFK;  //complement 
assign CQC = ~cqc;  //complement 
assign CQK = ~cqk;  //complement 
assign DGC =  PDC & PHC & plc  ; 
assign dgc = ~DGC;  //complement  
assign DGK =  PBC & PHC & pnc  ; 
assign dgk = ~DGK;  //complement 
assign ecc = ~ECC;  //complement 
assign eck = ~ECK;  //complement 
assign EDC = ~edc;  //complement 
assign edk = ~EDK;  //complement 
assign tes =  WAC & QFB  |  WBC & QFC  ; 
assign TES = ~tes;  //complement 
assign tec =  WAC & QFB  |  WBC & QFC  ; 
assign TEC = ~tec; //complement 
assign tek =  WAC & QFB  |  WBC & QFC  ; 
assign TEK = ~tek;  //complement 
assign ebc = ~EBC;  //complement 
assign ebk = ~EBK;  //complement 
assign eac = ~EAC;  //complement 
assign eak = ~EAK;  //complement 
assign QFA = ~qfa;  //complement 
assign QFB = ~qfb;  //complement 
assign QFC = ~qfc;  //complement 
assign eec = ~EEC;  //complement 
assign eqc = ~EQC;  //complement 
assign eqk = ~EQK;  //complement 
assign glc = ~GLC;  //complement 
assign fdf =  ebk  ; 
assign FDF = ~fdf;  //complement  
assign fdl =  edc & eck  ; 
assign FDL = ~fdl;  //complement 
assign fds =  eec & edk  ; 
assign FDS = ~fds;  //complement  
assign fea =  ecd & ebk  ; 
assign FEA = ~fea;  //complement 
assign BAC =  AAK & RAA  |  ABK & RAB  |  ACK & RAC  |  ADK & RAD  ; 
assign bac = ~BAC;  //complement 
assign BBC =  AAK & RAA  |  ABK & RAB  |  ACK & RAC  |  ADK & RAD  ; 
assign bbc = ~BBC; //complement 
assign BCC =  AAK & RAA  |  ABK & RAB  |  ACK & RAC  |  ADK & RAD  ; 
assign bcc = ~BCC;  //complement 
assign aac = ~AAC;  //complement 
assign aak = ~AAK;  //complement 
assign abc = ~ABC;  //complement 
assign abk = ~ABK;  //complement 
assign BDC =  AAC & RAI  |  ABC & RAJ  |  ACC & RAK  |  ADC & RAL  ; 
assign bdc = ~BDC;  //complement 
assign acc = ~ACC;  //complement 
assign ack = ~ACK;  //complement 
assign adc = ~ADC;  //complement 
assign adk = ~ADK;  //complement 
assign rac = ~RAC;  //complement 
assign rak = ~RAK;  //complement 
assign ras = ~RAS;  //complement 
assign JAC =  raa & rab & rac & rad & QCB  ; 
assign jac = ~JAC;  //complement  
assign JBC =  RAS & qce  ; 
assign jbc = ~JBC;  //complement 
assign GQC = ~gqc;  //complement 
assign GQK = ~gqk;  //complement 
assign TCC =  wac & wbc  |  ZZO  |  ZZI & qeb  |  ZZI & qfc  ; 
assign tcc = ~TCC;  //complement 
assign TCK =  wac & wbc  |  ZZO  |  ZZI & qeb  |  ZZI & qfc  ; 
assign tck = ~TCK; //complement 
assign TCS =  wac & wbc  |  ZZO  |  ZZI & qeb  |  ZZI & qfc  ; 
assign tcs = ~TCS;  //complement 
assign MBC =  GAC & HAC  |  GBC & HBC  |  GCC & HCC  |  GDC & HDC  |  GEC & HEC  |  GFC & HFC  ;
assign mbc = ~MBC;  //complement 
assign ODD = ~odd;  //complement 
assign wcb = ~WCB;  //complement 
assign tjc =  ZZO  |  ZZO  |  ZZI & WCA  |  ZZI & WDA  ; 
assign TJC = ~tjc;  //complement 
assign tjk =  ZZO  |  ZZO  |  ZZI & WCA  |  ZZI & WDA  ; 
assign TJK = ~tjk; //complement 
assign tjs =  ZZO  |  ZZO  |  ZZI & WCA  |  ZZI & WDA  ; 
assign TJS = ~tjs;  //complement 
assign TGC =  wab & wbb & eac & eak  ; 
assign tgc = ~TGC;  //complement  
assign MAC =  GAC & HAC  |  GBC & HBC  |  GCC & HCC  |  GDC & HDC  |  GEC & HEC  |  GFC & HFC  ;
assign mac = ~MAC;  //complement 
assign wae = ~WAE;  //complement 
assign waf = ~WAF;  //complement 
assign TGS =  waf & wbf  ; 
assign tgs = ~TGS;  //complement  
assign TIC =  wca & wda & NAC  ; 
assign tic = ~TIC;  //complement 
assign gac = ~GAC;  //complement 
assign gdc = ~GDC;  //complement 
assign gec = ~GEC;  //complement 
assign ghc = ~GHC;  //complement 
assign gic = ~GIC;  //complement 
assign gbc = ~GBC;  //complement 
assign gfc = ~GFC;  //complement 
assign ggc = ~GGC;  //complement 
assign gjc = ~GJC;  //complement 
assign gkc = ~GKC;  //complement 
assign gcc = ~GCC;  //complement 
assign lcc = ~LCC;  //complement 
assign lfc = ~LFC;  //complement 
assign lmc = ~LMC;  //complement 
assign lnc = ~LNC;  //complement 
assign QAC = ~qac;  //complement 
assign QBC = ~qbc;  //complement 
assign kbc = ~KBC;  //complement 
assign kcc = ~KCC;  //complement 
assign kdc = ~KDC;  //complement 
assign kec = ~KEC;  //complement 
assign OAC = ~oac;  //complement 
assign OBC = ~obc;  //complement 
assign OCC = ~occ;  //complement 
assign owc = ~OWC;  //complement 
assign kac = ~KAC;  //complement 
assign kfc = ~KFC;  //complement 
assign lqc = ~LQC;  //complement 
assign lrc = ~LRC;  //complement 
assign OAK = ~oak;  //complement 
assign OBK = ~obk;  //complement 
assign OCK = ~ock;  //complement 
assign ofc = ~OFC;  //complement 
assign JLA = LQA; 
assign jla = ~JLA; //complement 
assign JLB = LQB; 
assign jlb = ~JLB;  //complement 
assign JLC = LQG & lqc ; 
assign jlc = ~JLC ;  //complement 
assign JLD = LQG & LQC; 
assign jld = ~JLD; 
assign kic = ~KIC;  //complement 
assign kjc = ~KJC;  //complement 
assign klc = ~KLC;  //complement 
assign lsc = ~LSC;  //complement 
assign kgc = ~KGC;  //complement 
assign khc = ~KHC;  //complement 
assign kkc = ~KKC;  //complement 
assign oec = ~OEC;  //complement 
assign hac = ~HAC;  //complement 
assign hbc = ~HBC;  //complement 
assign OUA = ~oua;  //complement 
assign OUB = ~oub;  //complement 
assign ogc = ~OGC;  //complement 
assign ohc = ~OHC;  //complement 
assign hcc = ~HCC;  //complement 
assign hdc = ~HDC;  //complement 
assign hfc = ~HFC;  //complement 
assign OPA = ~opa;  //complement 
assign OQA = ~oqa;  //complement 
assign OLC = ~olc;  //complement 
assign HEC = ~hec;  //complement 
assign owf = ~OWF;  //complement 
assign NIC = ~nic;  //complement 
assign jdi =  hfi  ; 
assign JDI = ~jdi;  //complement 
assign jdc =  hfc  ; 
assign JDC = ~jdc;  //complement 
assign JWC =  qga  ; 
assign jwc = ~JWC;  //complement 
assign hfi = ~HFI;  //complement 
assign ooc = ~OOC;  //complement 
assign oof = ~OOF;  //complement 
assign owt = ~OWT;  //complement 
assign NAC = ~nac;  //complement 
assign NCC = ~ncc;  //complement 
assign NDL = ~ndl;  //complement 
assign NEC = ~nec;  //complement 
assign NDC = ~ndc;  //complement 
assign OWI = ~owi;  //complement 
assign lhc = ~LHC;  //complement 
assign lbc = ~LBC;  //complement 
assign ldc = ~LDC;  //complement 
assign lec = ~LEC;  //complement 
assign lgc = ~LGC;  //complement 
assign lic = ~LIC;  //complement 
assign ljc = ~LJC;  //complement 
assign lkc = ~LKC;  //complement 
assign llc = ~LLC;  //complement 
assign loc = ~LOC;  //complement 
assign lpc = ~LPC;  //complement 
assign lac = ~LAC;  //complement 
assign pod = ~POD;  //complement 
assign poe = ~POE;  //complement 
assign pof = ~POF;  //complement 
assign pla = ~PLA;  //complement 
assign plb = ~PLB;  //complement 
assign plc = ~PLC;  //complement 
assign pha = ~PHA;  //complement 
assign phb = ~PHB;  //complement 
assign phc = ~PHC;  //complement 
assign pda = ~PDA;  //complement 
assign pdb = ~PDB;  //complement 
assign pdc = ~PDC;  //complement 
assign DAD =  PBD & pfc & pgc  ; 
assign dad = ~DAD;  //complement 
assign DAL =  PCD & PHD & PND  ; 
assign dal = ~DAL;  //complement 
assign DAT =  PDD & PND  ; 
assign dat = ~DAT;  //complement 
assign DBD =  PAD & PGD & PJD  ; 
assign dbd = ~DBD;  //complement 
assign DBL =  PCD & PED & PKD  ; 
assign dbl = ~DBL;  //complement 
assign DBT =  PAD & PFD & PKD  ; 
assign dbt = ~DBT;  //complement 
assign DCD =  PCD & PFD & PKD  ; 
assign dcd = ~DCD;  //complement 
assign DCL =  PDD & PFD & PND  ; 
assign dcl = ~DCL;  //complement 
assign DCT =  pbb & pca & PND  ; 
assign dct = ~DCT;  //complement 
assign phd = ~PHD;  //complement 
assign phe = ~PHE;  //complement 
assign DDD =  PBD & PFD & PKD & PMD  ; 
assign ddd = ~DDD;  //complement  
assign DDL =  PBD & PFD & PKD & pmb  ; 
assign ddl = ~DDL;  //complement 
assign DED =  PDD & PGD & PLD  ; 
assign ded = ~DED;  //complement  
assign DEL =  PDD & PGD & PKF  ; 
assign del = ~DEL;  //complement 
assign DFD =  PCD & ped & pgd & PJD  ; 
assign dfd = ~DFD;  //complement  
assign CQD = ~cqd;  //complement 
assign CQL = ~cql;  //complement 
assign ecd = ~ECD;  //complement 
assign ecl = ~ECL;  //complement 
assign edd = ~EDD;  //complement 
assign edl = ~EDL;  //complement 
assign ted =  WAC & QFB  |  WBC & QFF  ; 
assign TED = ~ted; //complement 
assign tel =  WAC & QFB  |  WBC & QFF  ; 
assign TEL = ~tel;  //complement 
assign ebd = ~EBD;  //complement 
assign ebl = ~EBL;  //complement 
assign ead = ~EAD;  //complement 
assign QFD = ~qfd;  //complement 
assign QFE = ~qfe;  //complement 
assign QFF = ~qff;  //complement 
assign eed = ~EED;  //complement 
assign eel = ~EEL;  //complement 
assign eqd = ~EQD;  //complement 
assign eql = ~EQL;  //complement 
assign FBA = ~EQF & ~EQE & ~EQD  ; 
assign FBB = ~EQF & ~EQE &  EQD  ; 
assign FBC = ~EQF &  EQE & ~EQD  ; 
assign FBD = ~EQF &  EQE &  EQD  ; 
assign FBE =  EQF & ~EQE & ~EQD  ; 
assign FBF =  EQF & ~EQE &  EQD ; 
assign FBG =  EQF &  EQE & ~EQD  ; 
assign FBH =  EQF &  EQE &  EQD ; 
assign gld = ~GLD;  //complement 
assign fdg =  ebc & ecd & ecc  ; 
assign FDG = ~fdg;  //complement  
assign fdm =  edd & ebi & edl & eed  ; 
assign FDM = ~fdm;  //complement 
assign fdo =  ebi & edl & eed  ; 
assign FDO = ~fdo;  //complement  
assign BAD =  AAL & RAA  |  ABL & RAB  |  ACL & RAC  |  ADL & RAD  ; 
assign bad = ~BAD;  //complement 
assign BBD =  AAL & RAA  |  ABL & RAB  |  ACL & RAC  |  ADL & RAD  ; 
assign bbd = ~BBD; //complement 
assign BCD =  AAL & RAA  |  ABL & RAB  |  ACL & RAC  |  ADL & RAD  ; 
assign bcd = ~BCD;  //complement 
assign aad = ~AAD;  //complement 
assign aal = ~AAL;  //complement 
assign abd = ~ABD;  //complement 
assign abl = ~ABL;  //complement 
assign BDD =  AAD & RAI  |  ABD & RAJ  |  ACD & RAK  |  ADD & RAL  ; 
assign bdd = ~BDD;  //complement 
assign acd = ~ACD;  //complement 
assign acl = ~ACL;  //complement 
assign add = ~ADD;  //complement 
assign adl = ~ADL;  //complement 
assign rad = ~RAD;  //complement 
assign ral = ~RAL;  //complement 
assign rat = ~RAT;  //complement 
assign JAD =  raa & rab & rac & rad & QCC  ; 
assign jad = ~JAD;  //complement  
assign JBD =  RAT & qce  ; 
assign jbd = ~JBD;  //complement 
assign GQD = ~gqd;  //complement 
assign GQL = ~gql;  //complement 
assign TCD =  wad & wbd  |  ZZO  |  ZZI & qec  |  ZZI & qfd  ; 
assign tcd = ~TCD;  //complement 
assign TCL =  wad & wbd  |  ZZO  |  ZZI & qec  |  ZZI & qfd  ; 
assign tcl = ~TCL; //complement 
assign TCT =  wad & wbd  |  ZZO  |  ZZI & qec  |  ZZI & qfd  ; 
assign tct = ~TCT;  //complement 
assign MBD =  GAD & HAD  |  GBD & HBD  |  GCD & HCD  |  GDD & HDD  |  GED & HED  |  GFD & HFD  ;
assign mbd = ~MBD;  //complement 
assign ODE = ~ode;  //complement 
assign wcc = ~WCC;  //complement 
assign tjd =  ZZO  |  ZZO  |  ZZI & WCB  |  ZZI & WDB  ; 
assign TJD = ~tjd;  //complement 
assign tjl =  ZZO  |  ZZO  |  ZZI & WCB  |  ZZI & WDB  ; 
assign TJL = ~tjl; //complement 
assign tjt =  ZZO  |  ZZO  |  ZZI & WCB  |  ZZI & WDB  ; 
assign TJT = ~tjt;  //complement 
assign TGD =  wab & wbb & ead  ; 
assign tgd = ~TGD;  //complement  
assign MAD =  GAD & HAD  |  GBD & HBD  |  GCD & HCD  |  GDD & HDD  |  GED & HED  |  GFD & HFD  ;
assign mad = ~MAD;  //complement 
assign wag = ~WAG;  //complement 
assign wah = ~WAH;  //complement 
assign TGT =  waf & wbf  ; 
assign tgt = ~TGT;  //complement  
assign TID =  wcb & wdb & NAD  ; 
assign tid = ~TID;  //complement 
assign gad = ~GAD;  //complement 
assign gdd = ~GDD;  //complement 
assign ged = ~GED;  //complement 
assign ghd = ~GHD;  //complement 
assign gid = ~GID;  //complement 
assign gbd = ~GBD;  //complement 
assign gfd = ~GFD;  //complement 
assign ggd = ~GGD;  //complement 
assign gjd = ~GJD;  //complement 
assign gkd = ~GKD;  //complement 
assign gcd = ~GCD;  //complement 
assign lcd = ~LCD;  //complement 
assign lmd = ~LMD;  //complement 
assign nka = ~NKA;  //complement 
assign nkb = ~NKB;  //complement 
assign nkc = ~NKC;  //complement 
assign nkd = ~NKD;  //complement 
assign QAD = ~qad;  //complement 
assign QBD = ~qbd;  //complement 
assign kbd = ~KBD;  //complement 
assign kcd = ~KCD;  //complement 
assign kdd = ~KDD;  //complement 
assign ked = ~KED;  //complement 
assign OAD = ~oad;  //complement 
assign OBD = ~obd;  //complement 
assign OCD = ~ocd;  //complement 
assign OWJ = ~owj;  //complement 
assign jga =  ggd  ; 
assign JGA = ~jga;  //complement 
assign JLE =  gid & ghd & NLD  ; 
assign jle = ~JLE;  //complement 
assign kad = ~KAD;  //complement 
assign kfd = ~KFD;  //complement 
assign lqd = ~LQD;  //complement 
assign lrd = ~LRD;  //complement 
assign OAL = ~oal;  //complement 
assign OBL = ~obl;  //complement 
assign OCL = ~ocl;  //complement 
assign ofd = ~OFD;  //complement 
assign JKE =  GGA & NKH  ; 
assign jke = ~JKE;  //complement 
assign JKH =  GGF & NKT  ; 
assign jkh = ~JKH;  //complement 
assign JMD =  gqk & gqj  ; 
assign jmd = ~JMD;  //complement 
assign kid = ~KID;  //complement 
assign kjd = ~KJD;  //complement 
assign kld = ~KLD;  //complement 
assign lsd = ~LSD;  //complement 
assign kgd = ~KGD;  //complement 
assign khd = ~KHD;  //complement 
assign kkd = ~KKD;  //complement 
assign oed = ~OED;  //complement 
assign had = ~HAD;  //complement 
assign hbd = ~HBD;  //complement 
assign OVA = ~ova;  //complement 
assign QGE = ~qge;  //complement 
assign qgc = ~QGC;  //complement 
assign ohd = ~OHD;  //complement 
assign jxa =  qgc & qge  ; 
assign JXA = ~jxa;  //complement 
assign hcd = ~HCD;  //complement 
assign hdd = ~HDD;  //complement 
assign HED = ~hed;  //complement 
assign hfd = ~HFD;  //complement 
assign qja = ~QJA;  //complement 
assign otc = ~OTC;  //complement 
assign OLD = ~old;  //complement 
assign osd = ~OSD;  //complement 
assign jma =  gdb & gfc & gdd & gie  ; 
assign JMA = ~jma;  //complement  
assign joc =  gql  ; 
assign JOC = ~joc;  //complement 
assign jpa =  ndd & nde & ndf  ; 
assign JPA = ~jpa;  //complement 
assign JWD =  qga & ndf  ; 
assign jwd = ~JWD;  //complement 
assign ojd = ~OJD;  //complement 
assign otg = ~OTG;  //complement 
assign oue = ~OUE;  //complement 
assign NAD = ~nad;  //complement 
assign NCD = ~ncd;  //complement 
assign NDD = ~ndd;  //complement 
assign lfd = ~LFD;  //complement 
assign NDG = ~ndg;  //complement 
assign OWK = ~owk;  //complement 
assign OWL = ~owl;  //complement 
assign lnd = ~LND;  //complement 
assign ldd = ~LDD;  //complement 
assign led = ~LED;  //complement 
assign lgd = ~LGD;  //complement 
assign lhd = ~LHD;  //complement 
assign lid = ~LID;  //complement 
assign ljd = ~LJD;  //complement 
assign lkd = ~LKD;  //complement 
assign lld = ~LLD;  //complement 
assign lod = ~LOD;  //complement 
assign lpd = ~LPD;  //complement 
assign pna = ~PNA;  //complement 
assign pnb = ~PNB;  //complement 
assign pnc = ~PNC;  //complement 
assign pid = ~PID;  //complement 
assign pie = ~PIE;  //complement 
assign pef = ~PEF;  //complement 
assign pad = ~PAD;  //complement 
assign pae = ~PAE;  //complement 
assign paf = ~PAF;  //complement 
assign DAM =  PCE & PGE & PIE  ; 
assign dam = ~DAM;  //complement 
assign DAU =  pce & pde & PIE  ; 
assign dau = ~DAU;  //complement 
assign DBE =  PCE & PGE & PNE  ; 
assign dbe = ~DBE;  //complement 
assign DBM =  PAE & PHE & PLE  ; 
assign dbm = ~DBM;  //complement 
assign DBU =  PCE & pee & PLE  ; 
assign dbu = ~DBU;  //complement 
assign DCE =  PDE & PHE & PKC  ; 
assign dce = ~DCE;  //complement 
assign DCM =  PCE & PEE & pne  ; 
assign dcm = ~DCM;  //complement 
assign DCU =  PDE & PGE & pne  ; 
assign dcu = ~DCU;  //complement 
assign pag = ~PAG;  //complement 
assign pah = ~PAH;  //complement 
assign DDE =  PAE & POE & PKE & pme  ; 
assign dde = ~DDE;  //complement  
assign DDM =  PBE & PEE & PLE & pme  ; 
assign ddm = ~DDM;  //complement 
assign DEE =  PDE & PEE & PME  ; 
assign dee = ~DEE;  //complement  
assign DEM =  PDE & PFE & PKE & pme  ; 
assign dem = ~DEM;  //complement 
assign DFE =  PBE & PFE & PJE & PME  ; 
assign dfe = ~DFE;  //complement  
assign DFM =  PAE & PEE & pie & ple  ; 
assign dfm = ~DFM;  //complement 
assign CQE = ~cqe;  //complement 
assign CQM = ~cqm;  //complement 
assign DGE =  PBE & PGE & PNE  ; 
assign dge = ~DGE;  //complement  
assign DGM =  PBE & PEE & PJE  ; 
assign dgm = ~DGM;  //complement 
assign ece = ~ECE;  //complement 
assign ecm = ~ECM;  //complement 
assign EDE = ~ede;  //complement 
assign edm = ~EDM;  //complement 
assign tee =  WAE & QFD  |  WBE & QFE  ; 
assign TEE = ~tee; //complement 
assign tem =  WAE & QFD  |  WBE & QFE  ; 
assign TEM = ~tem;  //complement 
assign ebe = ~EBE;  //complement 
assign ebm = ~EBM;  //complement 
assign eae = ~EAE;  //complement 
assign eam = ~EAM;  //complement 
assign QEA = ~qea;  //complement 
assign QEB = ~qeb;  //complement 
assign QEC = ~qec;  //complement 
assign eee = ~EEE;  //complement 
assign eem = ~EEM;  //complement 
assign eqe = ~EQE;  //complement 
assign eqm = ~EQM;  //complement 
assign gle = ~GLE;  //complement 
assign fdh =  ebm & ebl & ecm & ece & ecl  ; 
assign FDH = ~fdh;  //complement  
assign fde =  ebm & ece  ; 
assign FDE = ~fde;  //complement 
assign fdt =  ede & edm & eee & ecn & eem  ; 
assign FDT = ~fdt;  //complement  
assign fdv =  ede & edn & edm & eee  ; 
assign FDV = ~fdv;  //complement 
assign fdw =  ede & edm & eem & een & eee  ; 
assign FDW = ~fdw;  //complement  
assign BAE =  AAM & RAU  |  ABM & RAV  |  ACM & RAG  |  ADM & RAH  ; 
assign bae = ~BAE;  //complement 
assign BBE =  AAM & RAU  |  ABM & RAV  |  ACM & RAG  |  ADM & RAH  ; 
assign bbe = ~BBE; //complement 
assign BCE =  AAM & RAU  |  ABM & RAV  |  ACM & RAG  |  ADM & RAH  ; 
assign bce = ~BCE;  //complement 
assign aae = ~AAE;  //complement 
assign aam = ~AAM;  //complement 
assign abe = ~ABE;  //complement 
assign abm = ~ABM;  //complement 
assign BDE =  AAE & RAM  |  ABE & RAN  |  ACE & RAO  |  ADE & RAP  ; 
assign bde = ~BDE;  //complement 
assign ace = ~ACE;  //complement 
assign acm = ~ACM;  //complement 
assign ade = ~ADE;  //complement 
assign adm = ~ADM;  //complement 
assign rae = ~RAE;  //complement 
assign ram = ~RAM;  //complement 
assign rau = ~RAU;  //complement 
assign JAE =  rae & raf & rag & rah & QCC  ; 
assign jae = ~JAE;  //complement  
assign JBE =  QCA & QCE  ; 
assign jbe = ~JBE;  //complement 
assign GQE = ~gqe;  //complement 
assign GQM = ~gqm;  //complement 
assign TCE =  wad & wbd  |  ZZO  |  ZZI & qec  |  ZZI & qfe  ; 
assign tce = ~TCE;  //complement 
assign TCM =  wad & wbd  |  ZZO  |  ZZI & qec  |  ZZI & qfe  ; 
assign tcm = ~TCM; //complement 
assign TCU =  wad & wbd  |  ZZO  |  ZZI & qec  |  ZZI & qfe  ; 
assign tcu = ~TCU;  //complement 
assign MBE =  GAE & HAE  |  GBE & HBE  |  GCE & HCE  |  GDE & HDE  |  GEE & HEE  |  GFE & HFE  ;
assign mbe = ~MBE;  //complement 
assign ODF = ~odf;  //complement 
assign wda = ~WDA;  //complement 
assign tje =  ZZO  |  ZZO  |  ZZI & WCB  |  ZZI & WDB  ; 
assign TJE = ~tje;  //complement 
assign tjm =  ZZO  |  ZZO  |  ZZI & WCB  |  ZZI & WDB  ; 
assign TJM = ~tjm; //complement 
assign TGE =  wag & wbg & eae & eam  ; 
assign tge = ~TGE;  //complement  
assign MAE =  GAE & HAE  |  GBE & HBE  |  GCE & HCE  |  GDE & HDE  |  GEE & HEE  |  GFE & HFE  ;
assign mae = ~MAE;  //complement 
assign wba = ~WBA;  //complement 
assign wbb = ~WBB;  //complement 
assign TII =  wcc & wdc & GHE  ; 
assign tii = ~TII;  //complement  
assign TIE =  wcb & wdb  ; 
assign tie = ~TIE;  //complement 
assign gae = ~GAE;  //complement 
assign gde = ~GDE;  //complement 
assign gee = ~GEE;  //complement 
assign ghe = ~GHE;  //complement 
assign gie = ~GIE;  //complement 
assign gbe = ~GBE;  //complement 
assign gfe = ~GFE;  //complement 
assign gge = ~GGE;  //complement 
assign gje = ~GJE;  //complement 
assign gke = ~GKE;  //complement 
assign gce = ~GCE;  //complement 
assign lce = ~LCE;  //complement 
assign lfe = ~LFE;  //complement 
assign lme = ~LME;  //complement 
assign lne = ~LNE;  //complement 
assign nke = ~NKE;  //complement 
assign nkf = ~NKF;  //complement 
assign nkg = ~NKG;  //complement 
assign nkh = ~NKH;  //complement 
assign QAE = ~qae;  //complement 
assign QBE = ~qbe;  //complement 
assign OAE = ~oae;  //complement 
assign OBE = ~obe;  //complement 
assign OCE = ~oce;  //complement 
assign owm = ~OWM;  //complement 
assign jgb =  gde  ; 
assign JGB = ~jgb;  //complement 
assign JLF =  gge & ZZI & NLD  ; 
assign jlf = ~JLF;  //complement 
assign kfe = ~KFE;  //complement 
assign lqe = ~LQE;  //complement 
assign lre = ~LRE;  //complement 
assign OAM = ~oam;  //complement 
assign OBM = ~obm;  //complement 
assign OCM = ~ocm;  //complement 
assign ofe = ~OFE;  //complement 
assign JKF =  gga & NKH  ; 
assign jkf = ~JKF;  //complement 
assign JNB =  GQJ  ; 
assign jnb = ~JNB;  //complement 
assign JME =  GQK & GQJ  ; 
assign jme = ~JME;  //complement 
assign kie = ~KIE;  //complement 
assign kje = ~KJE;  //complement 
assign kle = ~KLE;  //complement 
assign lse = ~LSE;  //complement 
assign kge = ~KGE;  //complement 
assign khe = ~KHE;  //complement 
assign kke = ~KKE;  //complement 
assign oee = ~OEE;  //complement 
assign hae = ~HAE;  //complement 
assign hbe = ~HBE;  //complement 
assign ovb = ~OVB;  //complement 
assign ohe = ~OHE;  //complement 
assign hce = ~HCE;  //complement 
assign hde = ~HDE;  //complement 
assign HEE = ~hee;  //complement 
assign hfe = ~HFE;  //complement 
assign OJA = ~oja;  //complement 
assign OJB = ~ojb;  //complement 
assign OLE = ~ole;  //complement 
assign oma = ~OMA;  //complement 
assign jmb =  gfb & gfc & gda & gie  ; 
assign JMB = ~jmb;  //complement  
assign JNA =  GIE  ; 
assign jna = ~JNA;  //complement 
assign JWE =  qgb  ; 
assign jwe = ~JWE;  //complement 
assign NCE = ~nce;  //complement 
assign NDE = ~nde;  //complement 
assign NDH = ~ndh;  //complement 
assign lde = ~LDE;  //complement 
assign lee = ~LEE;  //complement 
assign lge = ~LGE;  //complement 
assign lhe = ~LHE;  //complement 
assign lie = ~LIE;  //complement 
assign lje = ~LJE;  //complement 
assign lke = ~LKE;  //complement 
assign lle = ~LLE;  //complement 
assign loe = ~LOE;  //complement 
assign lpe = ~LPE;  //complement 
assign OWU = ~owu;  //complement 
assign pnd = ~PND;  //complement 
assign pne = ~PNE;  //complement 
assign pnf = ~PNF;  //complement 
assign pjd = ~PJD;  //complement 
assign pje = ~PJE;  //complement 
assign pjf = ~PJF;  //complement 
assign pff = ~PFF;  //complement 
assign pfg = ~PFG;  //complement 
assign pfh = ~PFH;  //complement 
assign pbd = ~PBD;  //complement 
assign pbe = ~PBE;  //complement 
assign pbf = ~PBF;  //complement 
assign DAF =  PCF & PEF & plf  ; 
assign daf = ~DAF;  //complement 
assign DAN =  PBF & PFF & pnf  ; 
assign dan = ~DAN;  //complement 
assign DAV =  PCF & PGF & pnf  ; 
assign dav = ~DAV;  //complement 
assign DBF =  PCF & PHF & pnf  ; 
assign dbf = ~DBF;  //complement 
assign DBN =  PAF & PGF & PLF  ; 
assign dbn = ~DBN;  //complement 
assign DBV =  PCF & phf & PLF  ; 
assign dbv = ~DBV;  //complement 
assign DCF =  PBF & PEF & pnf  ; 
assign dcf = ~DCF;  //complement 
assign DCN =  PCF & PFF & PLF  ; 
assign dcn = ~DCN;  //complement 
assign DCV =  PDF & PFF & PLF  ; 
assign dcv = ~DCV;  //complement 
assign pbg = ~PBG;  //complement 
assign pbh = ~PBH;  //complement 
assign DDF =  PAF & PGF & PKF & PMF  ; 
assign ddf = ~DDF;  //complement  
assign DDN =  PBF & pef & phf & pmf  ; 
assign ddn = ~DDN;  //complement 
assign DEF =  PDF & POF & pnf & pmf  ; 
assign def = ~DEF;  //complement  
assign DCW =  PDF & PHF & PMF & plf  ; 
assign dcw = ~DCW;  //complement 
assign DFF =  PBF & pof & plf  ; 
assign dff = ~DFF;  //complement  
assign DFN =  PBF & PEF & PIE  ; 
assign dfn = ~DFN;  //complement 
assign CQF = ~cqf;  //complement 
assign CQN = ~cqn;  //complement 
assign ecf = ~ECF;  //complement 
assign ECN = ~ecn;  //complement 
assign edf = ~EDF;  //complement 
assign edn = ~EDN;  //complement 
assign tef =  WAE & QFD  |  WBE & QFE  ; 
assign TEF = ~tef; //complement 
assign ten =  WAE & QFD  |  WBE & QFE  ; 
assign TEN = ~ten;  //complement 
assign ebf = ~EBF;  //complement 
assign ebn = ~EBN;  //complement 
assign eaf = ~EAF;  //complement 
assign ean = ~EAN;  //complement 
assign QED = ~qed;  //complement 
assign QEE = ~qee;  //complement 
assign eef = ~EEF;  //complement 
assign een = ~EEN;  //complement 
assign eqf = ~EQF;  //complement 
assign eqn = ~EQN;  //complement 
assign glf = ~GLF;  //complement 
assign eeg = ~EEG;  //complement 
assign FDX =  EDN & EEB  ; 
assign fdx = ~FDX;  //complement  
assign fdd =  ebf & ebn & ecf  ; 
assign FDD = ~fdd;  //complement 
assign fdi =  ecn & edf  ; 
assign FDI = ~fdi;  //complement  
assign fdu =  eef & edo  ; 
assign FDU = ~fdu;  //complement 
assign BAF =  AAN & RAU  |  ABN & RAV  |  ACN & RAG  |  ADN & RAH  ; 
assign baf = ~BAF;  //complement 
assign BBF =  AAN & RAU  |  ABN & RAV  |  ACN & RAG  |  ADN & RAH  ; 
assign bbf = ~BBF; //complement 
assign BCF =  AAN & RAU  |  ABN & RAV  |  ACN & RAG  |  ADN & RAH  ; 
assign bcf = ~BCF;  //complement 
assign aaf = ~AAF;  //complement 
assign aan = ~AAN;  //complement 
assign abf = ~ABF;  //complement 
assign abn = ~ABN;  //complement 
assign BDF =  AAF & RAM  |  ABF & RAN  |  ACF & RAO  |  ADF & RAP  ; 
assign bdf = ~BDF;  //complement 
assign acf = ~ACF;  //complement 
assign acn = ~ACN;  //complement 
assign adf = ~ADF;  //complement 
assign adn = ~ADN;  //complement 
assign raf = ~RAF;  //complement 
assign ran = ~RAN;  //complement 
assign rav = ~RAV;  //complement 
assign JAG =  rae & raf & rag & rah & QCC  ; 
assign jag = ~JAG;  //complement  
assign jaf =  rae & raf & rag & rah  ; 
assign JAF = ~jaf;  //complement 
assign GQF = ~gqf;  //complement 
assign GQN = ~gqn;  //complement 
assign TCF =  wad & wbd  |  ZZO  |  ZZI & qec  |  ZZI & qfe  ; 
assign tcf = ~TCF;  //complement 
assign TCN =  wad & wbd  |  ZZO  |  ZZI & qec  |  ZZI & qfe  ; 
assign tcn = ~TCN; //complement 
assign TCV =  wad & wbd  |  ZZO  |  ZZI & qec  |  ZZI & qfe  ; 
assign tcv = ~TCV;  //complement 
assign MBF =  GAF & HAF  |  GBF & HBF  |  GCF & HCF  |  GDF & HDF  |  GEF & HEF  |  GFF & HFF  ;
assign mbf = ~MBF;  //complement 
assign ODG = ~odg;  //complement 
assign wdb = ~WDB;  //complement 
assign tjf =  ZZO  |  ZZO  |  ZZI & WCC  |  ZZI & WDC  ; 
assign TJF = ~tjf;  //complement 
assign tjn =  ZZO  |  ZZO  |  ZZI & WCC  |  ZZI & WDC  ; 
assign TJN = ~tjn; //complement 
assign TGF =  wag & wbg & eaf  ; 
assign tgf = ~TGF;  //complement  
assign MAF =  GAF & HAF  |  GBF & HBF  |  GCF & HCF  |  GDF & HDF  |  GEF & HEF  |  GFF & HFF  ;
assign maf = ~MAF;  //complement 
assign wbc = ~WBC;  //complement 
assign wbd = ~WBD;  //complement 
assign TIJ =  wcc & wdc & GHF  ; 
assign tij = ~TIJ;  //complement  
assign TIF =  wcb & wdb  ; 
assign tif = ~TIF;  //complement 
assign gaf = ~GAF;  //complement 
assign gdf = ~GDF;  //complement 
assign gef = ~GEF;  //complement 
assign ghf = ~GHF;  //complement 
assign gif = ~GIF;  //complement 
assign gbf = ~GBF;  //complement 
assign gff = ~GFF;  //complement 
assign ggf = ~GGF;  //complement 
assign gjf = ~GJF;  //complement 
assign gkf = ~GKF;  //complement 
assign gcf = ~GCF;  //complement 
assign lcf = ~LCF;  //complement 
assign lff = ~LFF;  //complement 
assign lmf = ~LMF;  //complement 
assign nki = ~NKI;  //complement 
assign nkj = ~NKJ;  //complement 
assign nkk = ~NKK;  //complement 
assign nkl = ~NKL;  //complement 
assign QAF = ~qaf;  //complement 
assign QBF = ~qbf;  //complement 
assign kbf = ~KBF;  //complement 
assign kcf = ~KCF;  //complement 
assign kdf = ~KDF;  //complement 
assign kef = ~KEF;  //complement 
assign OAF = ~oaf;  //complement 
assign OBF = ~obf;  //complement 
assign OCF = ~ocf;  //complement 
assign own = ~OWN;  //complement 
assign jgc =  gdf  ; 
assign JGC = ~jgc;  //complement 
assign JLG =  gid & gge & NLD  ; 
assign jlg = ~JLG;  //complement 
assign kaf = ~KAF;  //complement 
assign kff = ~KFF;  //complement 
assign lqf = ~LQF;  //complement 
assign lrf = ~LRF;  //complement 
assign OAN = ~oan;  //complement 
assign OBN = ~obn;  //complement 
assign OCN = ~ocn;  //complement 
assign off = ~OFF;  //complement 
assign JKG =  gib & NKL  ; 
assign jkg = ~JKG;  //complement 
assign JKI =  ggf & NKT  ; 
assign jki = ~JKI;  //complement 
assign JMF =  GQK  ; 
assign jmf = ~JMF;  //complement 
assign kif = ~KIF;  //complement 
assign kjf = ~KJF;  //complement 
assign klf = ~KLF;  //complement 
assign lsf = ~LSF;  //complement 
assign kgf = ~KGF;  //complement 
assign khf = ~KHF;  //complement 
assign kkf = ~KKF;  //complement 
assign oef = ~OEF;  //complement 
assign haf = ~HAF;  //complement 
assign hbf = ~HBF;  //complement 
assign ovc = ~OVC;  //complement 
assign ohf = ~OHF;  //complement 
assign hcf = ~HCF;  //complement 
assign hdf = ~HDF;  //complement 
assign HEF = ~hef;  //complement 
assign hff = ~HFF;  //complement 
assign qia = ~QIA;  //complement 
assign qib = ~QIB;  //complement 
assign OLF = ~olf;  //complement 
assign omb = ~OMB;  //complement 
assign jmc =  gdc & gdd & gda & gie  ; 
assign JMC = ~jmc;  //complement  
assign jfd =  qia & qic & qid & qie  ; 
assign JFD = ~jfd;  //complement 
assign JWF =  qgb  ; 
assign jwf = ~JWF;  //complement 
assign qic = ~QIC;  //complement 
assign qid = ~QID;  //complement 
assign QIE = ~qie;  //complement 
assign ONB = ~onb;  //complement 
assign ows = ~OWS;  //complement 
assign NCF = ~ncf;  //complement 
assign NDF = ~ndf;  //complement 
assign NDI = ~ndi;  //complement 
assign lnf = ~LNF;  //complement 
assign ldf = ~LDF;  //complement 
assign lef = ~LEF;  //complement 
assign lgf = ~LGF;  //complement 
assign lif = ~LIF;  //complement 
assign ljf = ~LJF;  //complement 
assign lkf = ~LKF;  //complement 
assign llf = ~LLF;  //complement 
assign lof = ~LOF;  //complement 
assign lpf = ~LPF;  //complement 
assign OWV = ~owv;  //complement 
assign pma = ~PMA;  //complement 
assign pmb = ~PMB;  //complement 
assign pmc = ~PMC;  //complement 
assign pkd = ~PKD;  //complement 
assign pke = ~PKE;  //complement 
assign pkf = ~PKF;  //complement 
assign pgf = ~PGF;  //complement 
assign pgg = ~PGG;  //complement 
assign pcd = ~PCD;  //complement 
assign pce = ~PCE;  //complement 
assign pcf = ~PCF;  //complement 
assign DAG =  PBG & PHG & plf  ; 
assign dag = ~DAG;  //complement 
assign DAO =  PDG & PHG & PLA  ; 
assign dao = ~DAO;  //complement 
assign DAW =  pdg & PLA  ; 
assign daw = ~DAW;  //complement 
assign DBG =  PBG & POD & PMF  ; 
assign dbg = ~DBG;  //complement 
assign pcg = ~PCG;  //complement 
assign DDG =  PAG & PGG & PKF & pmf  ; 
assign ddg = ~DDG;  //complement  
assign DDO =  PBG & PFG & PLA & PMF  ; 
assign ddo = ~DDO;  //complement 
assign DFG =  PBG & pof & PKC  ; 
assign dfg = ~DFG;  //complement  
assign CQG = ~cqg;  //complement 
assign CQO = ~cqo;  //complement 
assign ecg = ~ECG;  //complement 
assign eco = ~ECO;  //complement 
assign edg = ~EDG;  //complement 
assign edo = ~EDO;  //complement 
assign teg =  WAG & QFD  |  WBG & QFE  ; 
assign TEG = ~teg; //complement 
assign teo =  WAG & QFD  |  WBG & QFE  ; 
assign TEO = ~teo;  //complement 
assign ebg = ~EBG;  //complement 
assign eag = ~EAG;  //complement 
assign thk =  WAH  |  WBH  ; 
assign THK = ~thk;  //complement 
assign thf =  WAH  |  WBH  ; 
assign THF = ~thf; //complement 
assign the =  WAH  |  WBH  ; 
assign THE = ~the;  //complement 
assign eqg = ~EQG;  //complement 
assign eqo = ~EQO;  //complement 
assign glg = ~GLG;  //complement 
assign fdq =  ecc & ecg & edg  ; 
assign FDQ = ~fdq;  //complement  
assign FDA =  EAN & ecn & edf  ; 
assign fda = ~FDA;  //complement  
assign BAG =  AAO & RAE  |  ABO & RAF  |  ACO & RAW  |  ADO & RAX  ; 
assign bag = ~BAG;  //complement 
assign BBG =  AAO & RAE  |  ABO & RAF  |  ACO & RAW  |  ADO & RAX  ; 
assign bbg = ~BBG; //complement 
assign BCG =  AAO & RAE  |  ABO & RAF  |  ACO & RAW  |  ADO & RAX  ; 
assign bcg = ~BCG;  //complement 
assign aag = ~AAG;  //complement 
assign aao = ~AAO;  //complement 
assign abg = ~ABG;  //complement 
assign abo = ~ABO;  //complement 
assign BDG =  AAG & RAM  |  ABG & RAN  |  ACG & RAO  |  ADG & RAP  ; 
assign bdg = ~BDG;  //complement 
assign acg = ~ACG;  //complement 
assign aco = ~ACO;  //complement 
assign adg = ~ADG;  //complement 
assign ado = ~ADO;  //complement 
assign rag = ~RAG;  //complement 
assign rao = ~RAO;  //complement 
assign raw = ~RAW;  //complement 
assign qcd = ~QCD;  //complement 
assign qce = ~QCE;  //complement 
assign GQG = ~gqg;  //complement 
assign GQO = ~gqo;  //complement 
assign TCG =  wae & wbe  |  ZZO  |  ZZI & qed  |  ZZI & qff  ; 
assign tcg = ~TCG;  //complement 
assign TCO =  wae & wbe  |  ZZO  |  ZZI & qed  |  ZZI & qff  ; 
assign tco = ~TCO; //complement 
assign TCW =  wae & wbe  |  ZZO  |  ZZI & qed  |  ZZI & qff  ; 
assign tcw = ~TCW;  //complement 
assign MBG =  GAG & HAG  |  GBG & HBG  |  GCG & HCG  |  GDG & HDG  |  GFI & HFI  |  ZZI & HFG  ;
assign mbg = ~MBG;  //complement 
assign ODH = ~odh;  //complement 
assign wdc = ~WDC;  //complement 
assign tjg =  ZZO  |  ZZO  |  ZZI & WCC  |  ZZI & WDC  ; 
assign TJG = ~tjg;  //complement 
assign tjo =  ZZO  |  ZZO  |  ZZI & WCC  |  ZZI & WDC  ; 
assign TJO = ~tjo; //complement 
assign TGG =  wah & wbh & eag  ; 
assign tgg = ~TGG;  //complement  
assign MAG =  GAG & HAG  |  GBG & HBG  |  GCG & HCG  |  GDG & HDG  |  GFI & HFI  |  ZZI & HFG  ;
assign mag = ~MAG;  //complement 
assign wbe = ~WBE;  //complement 
assign wbf = ~WBF;  //complement 
assign NEI = ~nei;  //complement 
assign NKU = ~nku;  //complement 
assign gag = ~GAG;  //complement 
assign gdg = ~GDG;  //complement 
assign geg = ~GEG;  //complement 
assign ghg = ~GHG;  //complement 
assign gig = ~GIG;  //complement 
assign gbg = ~GBG;  //complement 
assign gfi = ~GFI;  //complement 
assign ggg = ~GGG;  //complement 
assign gjg = ~GJG;  //complement 
assign gkg = ~GKG;  //complement 
assign gcg = ~GCG;  //complement 
assign lcg = ~LCG;  //complement 
assign lfg = ~LFG;  //complement 
assign lmg = ~LMG;  //complement 
assign lng = ~LNG;  //complement 
assign nkm = ~NKM;  //complement 
assign nkn = ~NKN;  //complement 
assign nko = ~NKO;  //complement 
assign nkp = ~NKP;  //complement 
assign QAG = ~qag;  //complement 
assign QBG = ~qbg;  //complement 
assign kbg = ~KBG;  //complement 
assign kcg = ~KCG;  //complement 
assign kdg = ~KDG;  //complement 
assign keg = ~KEG;  //complement 
assign OAG = ~oag;  //complement 
assign OBG = ~obg;  //complement 
assign OCG = ~ocg;  //complement 
assign owo = ~OWO;  //complement 
assign jgd =  gdg  ; 
assign JGD = ~jgd;  //complement 
assign kag = ~KAG;  //complement 
assign kfg = ~KFG;  //complement 
assign lqg = ~LQG;  //complement 
assign OAO = ~oao;  //complement 
assign OBO = ~obo;  //complement 
assign OCO = ~oco;  //complement 
assign JOA =  GQJ  ; 
assign joa = ~JOA;  //complement 
assign kig = ~KIG;  //complement 
assign kjg = ~KJG;  //complement 
assign kgg = ~KGG;  //complement 
assign khg = ~KHG;  //complement 
assign hag = ~HAG;  //complement 
assign hbg = ~HBG;  //complement 
assign ovd = ~OVD;  //complement 
assign ohg = ~OHG;  //complement 
assign hcg = ~HCG;  //complement 
assign hdg = ~HDG;  //complement 
assign hfg = ~HFG;  //complement 
assign OJC = ~ojc;  //complement 
assign OWR = ~owr;  //complement 
assign OLG = ~olg;  //complement 
assign ord = ~ORD;  //complement 
assign nag = ~NAG;  //complement 
assign NAB = ~nab;  //complement 
assign JWG =  qgb  ; 
assign jwg = ~JWG;  //complement 
assign QKA = ~qka;  //complement 
assign QKB = ~qkb;  //complement 
assign NCG = ~ncg;  //complement 
assign TIG =  wcc & wdc & NAG  ; 
assign tig = ~TIG;  //complement  
assign ote = ~OTE;  //complement 
assign ouc = ~OUC;  //complement 
assign ove = ~OVE;  //complement 
assign opb = ~OPB;  //complement 
assign oqb = ~OQB;  //complement 
assign orb = ~ORB;  //complement 
assign osb = ~OSB;  //complement 
assign lhf = ~LHF;  //complement 
assign lhg = ~LHG;  //complement 
assign LBG = ~lbg;  //complement 
assign ldg = ~LDG;  //complement 
assign leg = ~LEG;  //complement 
assign lgg = ~LGG;  //complement 
assign lig = ~LIG;  //complement 
assign ljg = ~LJG;  //complement 
assign lkg = ~LKG;  //complement 
assign llg = ~LLG;  //complement 
assign log = ~LOG;  //complement 
assign lpg = ~LPG;  //complement 
assign OWW = ~oww;  //complement 
assign pmd = ~PMD;  //complement 
assign pme = ~PME;  //complement 
assign pmf = ~PMF;  //complement 
assign pld = ~PLD;  //complement 
assign ple = ~PLE;  //complement 
assign plf = ~PLF;  //complement 
assign phf = ~PHF;  //complement 
assign phg = ~PHG;  //complement 
assign phh = ~PHH;  //complement 
assign pdd = ~PDD;  //complement 
assign pde = ~PDE;  //complement 
assign pdf = ~PDF;  //complement 
assign DAH =  PBH & PHH & PJF  ; 
assign dah = ~DAH;  //complement 
assign DAP =  PDH & pfh & pme  ; 
assign dap = ~DAP;  //complement 
assign DBH =  PDH & POD & PNF  ; 
assign dbh = ~DBH;  //complement 
assign DBP =  PDH & PHH & PLF  ; 
assign dbp = ~DBP;  //complement 
assign pdg = ~PDG;  //complement 
assign pdh = ~PDH;  //complement 
assign DDH =  PBH & PHH & pld & pme  ; 
assign ddh = ~DDH;  //complement  
assign DDP =  PAH & PHH & PKE & PMF  ; 
assign ddp = ~DDP;  //complement 
assign CQH = ~cqh;  //complement 
assign CQP = ~cqp;  //complement 
assign edh = ~EDH;  //complement 
assign edp = ~EDP;  //complement 
assign teh =  WAG & QFD  |  WBG & QFE  ; 
assign TEH = ~teh; //complement 
assign tep =  WAG & QFD  |  WBG & QFE  ; 
assign TEP = ~tep;  //complement 
assign eah = ~EAH;  //complement 
assign eap = ~EAP;  //complement 
assign thl =  WAH  |  WBH  ; 
assign THL = ~thl;  //complement 
assign thh =  WAH  |  WBH  ; 
assign THH = ~thh; //complement 
assign thg =  WAH  |  WBH  ; 
assign THG = ~thg;  //complement 
assign eqh = ~EQH;  //complement 
assign eqp = ~EQP;  //complement 
assign FAA = ~EQI & ~EQH & ~EQG  ; 
assign FAB = ~EQI & ~EQH &  EQG  ; 
assign FAC = ~EQI &  EQH & ~EQG  ; 
assign FAD = ~EQI &  EQH &  EQG  ; 
assign FAE =  EQI & ~EQH & ~EQG  ; 
assign FAF =  EQI & ~EQH &  EQG ; 
assign FAG =  EQI &  EQH & ~EQG  ; 
assign FAH =  EQI &  EQH &  EQG ; 
assign glh = ~GLH;  //complement 
assign fdp =  eap  ; 
assign FDP = ~fdp;  //complement  
assign BAH =  AAP & RAE  |  ABP & RAF  |  ACP & RAW  |  ADP & RAX  ; 
assign bah = ~BAH;  //complement 
assign BBH =  AAP & RAE  |  ABP & RAF  |  ACP & RAW  |  ADP & RAX  ; 
assign bbh = ~BBH; //complement 
assign BCH =  AAP & RAE  |  ABP & RAF  |  ACP & RAW  |  ADP & RAX  ; 
assign bch = ~BCH;  //complement 
assign aah = ~AAH;  //complement 
assign aap = ~AAP;  //complement 
assign abh = ~ABH;  //complement 
assign abp = ~ABP;  //complement 
assign BDH =  AAH & RAM  |  ABH & RAN  |  ACH & RAO  |  ADH & RAP  ; 
assign bdh = ~BDH;  //complement 
assign ach = ~ACH;  //complement 
assign acp = ~ACP;  //complement 
assign adh = ~ADH;  //complement 
assign adp = ~ADP;  //complement 
assign rah = ~RAH;  //complement 
assign rap = ~RAP;  //complement 
assign rax = ~RAX;  //complement 
assign qca = ~QCA;  //complement 
assign qcb = ~QCB;  //complement 
assign qcc = ~QCC;  //complement 
assign GQH = ~gqh;  //complement 
assign GQP = ~gqp;  //complement 
assign TCH =  wae & wbe  |  ZZO  |  ZZI & qed  |  ZZI & qff  ; 
assign tch = ~TCH;  //complement 
assign TCP =  wae & wbe  |  ZZO  |  ZZI & qed  |  ZZI & qff  ; 
assign tcp = ~TCP; //complement 
assign TCX =  wae & wbe  |  ZZO  |  ZZI & qed  |  ZZI & qff  ; 
assign tcx = ~TCX;  //complement 
assign MBH =  GAH & HAH  |  GBH & HBH  |  GCH & HCH  |  GDH & HDH  |  GIG & QKB  |  ZZI & HFH  ;
assign mbh = ~MBH;  //complement 
assign ODI = ~odi;  //complement 
assign ODJ = ~odj;  //complement 
assign tjh =  ZZO  |  ZZO  |  ZZI & WCC  |  ZZI & WDC  ; 
assign TJH = ~tjh;  //complement 
assign tjp =  ZZO  |  ZZO  |  ZZI & WCC  |  ZZI & WDC  ; 
assign TJP = ~tjp; //complement 
assign TGH =  wah & wbh & eah  ; 
assign tgh = ~TGH;  //complement  
assign MAH =  GAH & HAH  |  GBH & HBH  |  GCH & HCH  |  GDH & HDH  |  GIG & QKB  |  ZZI & HFH  ;
assign mah = ~MAH;  //complement 
assign wbg = ~WBG;  //complement 
assign wbh = ~WBH;  //complement 
assign gah = ~GAH;  //complement 
assign gdh = ~GDH;  //complement 
assign ghh = ~GHH;  //complement 
assign gih = ~GIH;  //complement 
assign gbh = ~GBH;  //complement 
assign ggh = ~GGH;  //complement 
assign gjh = ~GJH;  //complement 
assign gch = ~GCH;  //complement 
assign jgi =  GQP  ; 
assign JGI = ~jgi;  //complement 
assign nkq = ~NKQ;  //complement 
assign nkr = ~NKR;  //complement 
assign nks = ~NKS;  //complement 
assign nkt = ~NKT;  //complement 
assign QAH = ~qah;  //complement 
assign QBH = ~qbh;  //complement 
assign qma = ~QMA;  //complement 
assign qmb = ~QMB;  //complement 
assign qmc = ~QMC;  //complement 
assign qmd = ~QMD;  //complement 
assign OAH = ~oah;  //complement 
assign OBH = ~obh;  //complement 
assign OCH = ~och;  //complement 
assign jge =  gdh  ; 
assign JGE = ~jge;  //complement 
assign OAP = ~oap;  //complement 
assign OBP = ~obp;  //complement 
assign OCP = ~ocp;  //complement 
assign JOB =  GQK  ; 
assign job = ~JOB;  //complement 
assign QDA = ~qda;  //complement 
assign QDB = ~qdb;  //complement 
assign QDC = ~qdc;  //complement 
assign QDD = ~qdd;  //complement 
assign OKA = ~oka;  //complement 
assign hah = ~HAH;  //complement 
assign hbh = ~HBH;  //complement 
assign qla = ~QLA;  //complement 
assign qlb = ~QLB;  //complement 
assign qlc = ~QLC;  //complement 
assign hch = ~HCH;  //complement 
assign hdh = ~HDH;  //complement 
assign hfh = ~HFH;  //complement 
assign qga = ~QGA;  //complement 
assign qgb = ~QGB;  //complement 
assign OLH = ~olh;  //complement 
assign oxc = ~OXC;  //complement 
assign thm =  WAF  |  WBF  ; 
assign THM = ~thm;  //complement 
assign JWH =  qgb  ; 
assign jwh = ~JWH;  //complement 
assign oia = ~OIA;  //complement 
assign oib = ~OIB;  //complement 
assign OWP = ~owp;  //complement 
assign owq = ~OWQ;  //complement 
assign NEE = ~nee;  //complement 
assign NCH = ~nch;  //complement 
assign otf = ~OTF;  //complement 
assign oud = ~OUD;  //complement 
assign ovf = ~OVF;  //complement 
assign OWX = ~owx;  //complement 
assign opc = ~OPC;  //complement 
assign oqc = ~OQC;  //complement 
assign orc = ~ORC;  //complement 
assign osc = ~OSC;  //complement 
assign iaa = ~IAA; //complement 
assign iab = ~IAB; //complement 
assign iac = ~IAC; //complement 
assign iad = ~IAD; //complement 
assign iae = ~IAE; //complement 
assign iaf = ~IAF; //complement 
assign iag = ~IAG; //complement 
assign iah = ~IAH; //complement 
assign iai = ~IAI; //complement 
assign iaj = ~IAJ; //complement 
assign iak = ~IAK; //complement 
assign ial = ~IAL; //complement 
assign iam = ~IAM; //complement 
assign ian = ~IAN; //complement 
assign iao = ~IAO; //complement 
assign iap = ~IAP; //complement 
assign iba = ~IBA; //complement 
assign ibb = ~IBB; //complement 
assign ibc = ~IBC; //complement 
assign ibd = ~IBD; //complement 
assign ibe = ~IBE; //complement 
assign ibf = ~IBF; //complement 
assign ibg = ~IBG; //complement 
assign ibh = ~IBH; //complement 
assign ibi = ~IBI; //complement 
assign ibj = ~IBJ; //complement 
assign ibk = ~IBK; //complement 
assign ibl = ~IBL; //complement 
assign ibm = ~IBM; //complement 
assign ibn = ~IBN; //complement 
assign ibo = ~IBO; //complement 
assign ibp = ~IBP; //complement 
assign ica = ~ICA; //complement 
assign icb = ~ICB; //complement 
assign icc = ~ICC; //complement 
assign icd = ~ICD; //complement 
assign ice = ~ICE; //complement 
assign icf = ~ICF; //complement 
assign icg = ~ICG; //complement 
assign ich = ~ICH; //complement 
assign ici = ~ICI; //complement 
assign icj = ~ICJ; //complement 
assign ick = ~ICK; //complement 
assign icl = ~ICL; //complement 
assign icm = ~ICM; //complement 
assign icn = ~ICN; //complement 
assign ico = ~ICO; //complement 
assign icp = ~ICP; //complement 
assign ida = ~IDA; //complement 
assign idb = ~IDB; //complement 
assign idc = ~IDC; //complement 
assign idd = ~IDD; //complement 
assign ide = ~IDE; //complement 
assign idf = ~IDF; //complement 
assign idg = ~IDG; //complement 
assign idh = ~IDH; //complement 
assign idi = ~IDI; //complement 
assign idj = ~IDJ; //complement 
assign idk = ~IDK; //complement 
assign idl = ~IDL; //complement 
assign idm = ~IDM; //complement 
assign idn = ~IDN; //complement 
assign ido = ~IDO; //complement 
assign idp = ~IDP; //complement 
assign iea = ~IEA; //complement 
assign ieb = ~IEB; //complement 
assign iec = ~IEC; //complement 
assign ied = ~IED; //complement 
assign iee = ~IEE; //complement 
assign ief = ~IEF; //complement 
assign ieg = ~IEG; //complement 
assign ieh = ~IEH; //complement 
assign ifa = ~IFA; //complement 
assign ifb = ~IFB; //complement 
assign ifc = ~IFC; //complement 
assign ifd = ~IFD; //complement 
assign iga = ~IGA; //complement 
assign igb = ~IGB; //complement 
assign ija = ~IJA; //complement 
assign ijb = ~IJB; //complement 
assign ijc = ~IJC; //complement 
assign ijd = ~IJD; //complement 
assign ije = ~IJE; //complement 
assign ijj = ~IJJ; //complement 
assign ijk = ~IJK; //complement 
assign ika = ~IKA; //complement 
assign ikb = ~IKB; //complement 
assign ikc = ~IKC; //complement 
assign ikq = ~IKQ; //complement 
assign ila = ~ILA; //complement 
assign izz = ~IZZ; //complement 
always@(posedge IZZ )
   begin 
 PIA <=  bbd & bbc & TCQ  |  PIA & tcq  ; 
 PIB <=  bbd & bbc & TCQ  |  PIA & tcq  ; 
 PIC <=  bbd & bbc & TCQ  |  PIA & tcq  ; 
 PEA <=  bbf & bbe & TCI  |  PEA & tci  ; 
 PEB <=  bbf & bbe & TCI  |  PEA & tci  ; 
 PEC <=  bbf & bbe & TCI  |  PEA & tci  ; 
 PAA <=  bbh & bbg & TCI  |  PAA & tci  ; 
 PAB <=  bbh & bbg & TCI  |  PAA & tci  ; 
 PAC <=  bbh & bbg & TCI  |  PAA & tci  ; 
 PED <=  bcf & bce & TCI  |  PED & tci  ; 
 PEE <=  bcf & bce & TCI  |  PED & tci  ; 
 cqa <=  bda & TCA  |  cqa & tca  ; 
 cqi <=  baa & TCA  |  cqi & tca  ; 
 ECA <=  DAA & TEI  |  ECA & tei  ; 
 ECI <=  DEA & TEI  |  ECI & tei  ; 
 EDA <=  DBI & TEI  |  EDA & tei  ; 
 EDI <=  DAB & TEI  |  EDI & tei  ; 
 EBA <=  DDA & TEI  |  EBA & tei  ; 
 EBI <=  DAI & TEI  |  EBI & tei  ; 
 EAA <=  DAQ & dbq & dda & ZZI & TEQ  |  DDI & dda & ZZI & TEQ  |  DCQ & ZZI & TEQ  |  DCA & TEQ  |  EAA & teq  ; 
 EAI <=  DAW & daa & ZZI & ZZI & TEQ  |  DDK & ZZI & ZZI & TEQ  |  DAO & ZZI & TEQ  |  DCI & TEQ  |  EAI & teq  ; 
 EEA <=  DEI & TEA  |  EEA & tea  ; 
 EEI <=  DBA & TEA  |  EEI & tea  ; 
 EQA <=  CQA & TEA  |  EQA & tea  ; 
 EQI <=  CQI & TEA  |  EQI & tea  ; 
 GLA <=  FAA & EAP & THA  |  GLA & tha  ; 
 AAA <=  IAA & JAA  |  AAA & jaa  ; 
 AAI <=  IAI & JAA  |  AAI & jaa  ; 
 ABA <=  IBA & JAB  |  ABA & jab  ; 
 ABI <=  IBI & JAB  |  ABI & jab  ; 
 ACA <=  ICA & JAC  |  ACA & jac  ; 
 ACI <=  ICI & JAC  |  ACI & jac  ; 
 ADA <=  IDA & JAD  |  ADA & jad  ; 
 ADI <=  IDI & JAD  |  ADI & jad  ; 
 RAA <=  JAE & jbe  |  QDA & JBE  |  JBA & tca  ; 
 RAI <=  JAE & jbe  |  QDA & JBE  |  JBA & tca  ; 
 RAQ <=  JAE & jbe  |  QDA & JBE  |  JBA & tca  ; 
 oda <=  MBA  |  MBB  |  MBC  |  MBD  |  TJQ  ; 
 odb <=  MBA  |  MBB  |  MBC  |  MBD  |  TJQ  ; 
 WAA <=  MAA & JWA  |  MAB & JWA  |  MAC & JWA  |  MAD & JWA  |  TJQ  ; 
 WAB <=  MAA & JWA  |  MAB & JWA  |  MAC & JWA  |  MAD & JWA  |  TJQ  ; 
 GAA <=  FAA & TGA  |  FBA & TGB  |  FCA & TGC  |  GAA & tha  ; 
 GDA <=  FDJ & TGQ  |  GDA & tgq  ; 
 GEA <=  EBI & TGQ  |  GEA & tgq  ; 
 GHA <=  ECA & TGS  |  GHA & tgs  ; 
 GIA <=  ECI & TGS  |  GIA & tgs  ; 
 GBA <=  FAA & TGD  |  FBA & TGE  |  FCA & TGF  |  GBA & tha  ; 
 GFA <=  EEA & TGR  |  GFA & tgr  ; 
 GGA <=  EBA & TGR  |  GGA & tgr  ; 
 GJA <=  FDN & TGT  |  GJA & tgt  ; 
 GKA <=  EDA & TGT  |  GKA & tgt  ; 
 GCA <=  FAA & TGG  |  FBA & TGH  |  FCA & TGI  |  GCA & tha  ; 
 LCA <=  TIA & NIA  |  ZZO  |  LBA & LBG  ; 
 LFA <=  TIB & NIA  |  LEA  |  ZZO & LBG  ; 
 LMA <=  TIC & NIA  |  LLA  ; 
 LNA <=  TID & NIA  |  LMA  ; 
 NLA <= JGF & GQG ; 
 NLB <= JGF & GQH ; 
 NLC <= JGF & GQI ; 
 NLD <= JGF & ZZI ; 
 qaa <=  jkc & qma  |  JKB & qmb  |  JKA & qmc  ; 
 qba <=  jlc & qma  |  JLB & qmb  |  JLA & qmc  ; 
 KBA <= KAA ; 
 KCA <= KBA ; 
 KDA <= KCA ; 
 KEA <= KDA ; 
 oaa <= eqa ; 
 oba <= eqa ; 
 oca <= eqa ; 
 OWA <= GQA ; 
 KAA <=  NKA & TIE  ; 
 KFA <=  NKE & TIE  |  KEA  ; 
 LQA <=  NLA & TJI  |  LPA  ; 
 LRA <=  LQA & TJI  ; 
 oai <= eqi ; 
 obi <= eqi ; 
 oci <= eqi ; 
 OFA <= LSA ; 
 gqa <=  eqa & THI  |  gqa & thi  ; 
 gqi <=  eqi & THI  |  gqi & thi  ; 
 KIA <=  NKI & TIF  |  KHA  ; 
 KJA <=  NKM & TIF  |  KIA  ; 
 KLA <=  NKQ & TJI  |  KKA  ; 
 LSA <=  NLE & TJI  |  LRA  ; 
 KGA <= KFA ; 
 KHA <= KGA ; 
 KKA <= KJA ; 
 OEA <= KLA ; 
 HAA <=  TII & JCA  |  HAA & qaa  ; 
 HBA <=  TIJ & JCA  |  HBA & qaa  ; 
 otd <=  gka  |  tji  ; 
 qgd <=  tji  ; 
 OGA <=  GQA & TJI  |  ZZO & QGC  |  NDJ & QGD  ; 
 OHA <=  GQD & TJI  |  NDA & JXA  |  ZZO & QGD  ; 
 HCA <=  NCA & TJA  |  HCA & iea  ; 
 HDA <=  GJA & TJA  |  HDA & iea  ; 
 HFA <=  JFA & TJA  |  JDA & qhg  |  QHJ  |  QHL  ; 
 ota <=  gha  |  tja  ; 
 otb <=  gia  |  tja  ; 
 ola <=  gla & TJA  |  gca & tja  |  GLA & tja  ; 
 QHF <= IJE ; 
 QHK <= QHJ ; 
 hea <= ifd ; 
 OOA <= GQA ; 
 OOD <= GQD ; 
 OWD <= GQD ; 
 naa <= gea ; 
 nia <= gqg ; 
 nca <= gca ; 
 ndj <= gqd ; 
 QHJ <=  JFI & TJJ  ; 
 QHL <=  NEB & TJJ  ; 
 nda <=  gqg & GGG  |  gqa & ggg  ; 
 ona <= gfa ; 
 owg <= gqg ; 
 opd <= gqa ; 
 ose <= gqa ; 
 nea <= gfa ; 
 LBA <= LAA ; 
 LDA <= LCA ; 
 LEA <= LDA ; 
 LGA <= LFA ; 
 LIA <= LHA ; 
 LJA <= LIA ; 
 LKA <= LJA ; 
 LLA <= LKA ; 
 LOA <= LNA ; 
 LPA <= LOA ; 
 LAA <= IFA ; 
 PJA <=  bbd & BAC & TCR  |  PJA & tcr  ; 
 PJC <=  bbd & BAC & TCR  |  PJA & tcr  ; 
 PFA <=  bbf & BBE & TCJ  |  PFA & tcj  ; 
 PFB <=  bbf & BBE & TCJ  |  PFA & tcj  ; 
 PFC <=  bbf & BBE & TCJ  |  PFA & tcj  ; 
 PBA <=  bbh & BBG & TCJ  |  PBA & tcj  ; 
 PBB <=  bbh & BBG & TCJ  |  PBA & tcj  ; 
 PBC <=  bbh & BBG & TCJ  |  PBA & tcj  ; 
 PFD <=  bcf & BCE & TCJ  |  PFD & tcj  ; 
 PFE <=  bcf & BCE & TCJ  |  PFD & tcj  ; 
 cqb <=  bdb & TCB  |  cqb & tcb  ; 
 cqj <=  bab & TCB  |  cqj & tcb  ; 
 ECB <=  DAV & TEJ  |  ECB & tej  ; 
 ECJ <=  DCJ & TEJ  |  ECJ & tej  ; 
 EDB <=  DDJ & TEJ  |  EDB & tej  ; 
 EDJ <=  DFB & TEJ  |  EDJ & tej  ; 
 EBB <=  DBB & TEJ  |  EBB & tej  ; 
 EBJ <=  DEB & TEJ  |  EBJ & tej  ; 
 EAB <=  dab & ddb & daj & ZZI & TEB  |  ZZO & daj & ZZI & TEB  |  ZZO & ZZI & TEB  |  ZZO & TEB  |  EAB & teb  ; 
 eeb <=  dej & TEB  |  DEI & TEB  |  eeb & teb  ; 
 EEJ <=  DAR & TEB  |  ZZO & TEB  |  EEJ & teb  ; 
 EQB <=  CQB & TEB  |  EQB & teb  ; 
 EQJ <=  CQJ & TEB  |  EQJ & teb  ; 
 GLB <=  FAB & EAP & THB  |  GLB & thb  ; 
 AAB <=  IAB & JAA  |  AAB & jaa  ; 
 AAJ <=  IAJ & JAA  |  AAJ & jaa  ; 
 ABB <=  IBB & JAB  |  ABB & jab  ; 
 ABJ <=  IBJ & JAB  |  ABJ & jab  ; 
 ACB <=  ICB & JAC  |  ACB & jac  ; 
 ACJ <=  ICJ & JAC  |  ACJ & jac  ; 
 ADB <=  IDB & JAD  |  ADB & jad  ; 
 ADJ <=  IDJ & JAD  |  ADJ & jad  ; 
 RAB <=  JBA & TCB  |  QDB & JBE  |  JBB & tcb  ; 
 RAJ <=  JBA & TCB  |  QDB & JBE  |  JBB & tcb  ; 
 RAR <=  JBA & TCB  |  QDB & JBE  |  JBB & tcb  ; 
 gqb <=  eqb & THJ  |  gqb & thj  ; 
 gqj <=  eqj & THJ  |  gqj & thj  ; 
 odc <=  MBA  |  MBB  |  MBC  |  MBD  |  TJR  ; 
 WCA <=  MBA  |  MBB  |  MBC  |  MBD  |  TJR  ; 
 WAC <=  MAA & JWB  |  MAB & JWB  |  MAC & JWB  |  MAD & JWB  |  TJR  ; 
 WAD <=  MAA & JWB  |  MAB & JWB  |  MAC & JWB  |  MAD & JWB  |  TJR  ; 
 GAB <=  FAB & TGA  |  FBB & TGB  |  FCB & TGC  |  GAB & thb  ; 
 GDB <=  FDK & TGQ  |  GDB & tgq  ; 
 GEB <=  ECB & TGQ  |  GEB & tgq  ; 
 GHB <=  EEI & TGS  |  GHB & tgs  ; 
 GIB <=  EBJ & TGS  |  GIB & tgs  ; 
 GBB <=  FAB & TGD  |  FBB & TGE  |  FCB & TGF  |  GBB & thb  ; 
 GFB <=  FDR & TGR  |  GFB & tgr  ; 
 GGB <=  EBB & TGR  |  GGB & tgr  ; 
 GJB <=  FDK & TGT  |  GJB & tgt  ; 
 GKB <=  ECJ & TGT  |  GKB & tgt  ; 
 GCB <=  FAB & TGG  |  FBB & TGH  |  FCB & TGI  |  GCB & thb  ; 
 LCB <=  TIA & NIB  |  ZZO  |  LBB & LBG  ; 
 LFB <=  TIB & NIB  |  LEB  |  ZZO & LBG  ; 
 LMB <=  TIC & NIB  |  LLB  ; 
 LNB <=  TID & NIB  |  LMB  ; 
 NLE <= JGG & GQG ; 
 NLF <= JGG & GQH ; 
 NLG <= JGG & GQI ; 
 NLH <= JGG & ZZI ; 
 qab <=  jkc & qma  |  JKB & qmb  |  jka & qmc  ; 
 qbb <=  jlc & qma  |  JLB & qmb  |  jla & qmc  ; 
 KBB <= KAB ; 
 KCB <= KBB ; 
 KDB <= KCB ; 
 KEB <= KDB ; 
 oab <= eqb ; 
 obb <= eqb ; 
 ocb <= eqb ; 
 OWB <= GQB ; 
 KAB <=  NKB & TIE  ; 
 KFB <=  NKF & TIE  |  KEB  ; 
 LQB <=  NLB & TJJ  |  LPB  ; 
 LRB <=  LQB & TJJ  ; 
 oaj <= eqj ; 
 obj <= eqj ; 
 ocj <= eqj ; 
 OFB <= LSB ; 
 KIB <=  NKJ & TIF  |  KHB  ; 
 KJB <=  NKN & TIF  |  KIB  ; 
 KLB <=  NKR & TJJ  |  KKB  ; 
 LSB <=  NLF & TJJ  |  LRB  ; 
 KGB <= KFB ; 
 KHB <= KGB ; 
 KKB <= KJB ; 
 OEB <= KLB ; 
 HAB <=  TII & JCB  |  HAB & qab  ; 
 HBB <=  TIJ & JCB  |  HBB & qab  ; 
 QHA <=  QHF & TJJ  |  QHK  ; 
 QHB <=  JFB & TJJ  |  QHA  ; 
 OGB <=  GQB & TJJ  |  ZZO & QGC  |  NDK & QGD  ; 
 OOB <= GQB ; 
 OOE <= GQE ; 
 OWE <= GQE ; 
 HCB <=  NCB & TJB  |  HCB & ieb  ; 
 HDB <=  GJB & TJB  |  HDB & ieb  ; 
 heb <=  lcg & TJB  ; 
 HFB <=  JFC & TJB  |  JDB & qhd  |  QHJ  ; 
 ora <=  ghb  |  tjb  ; 
 osa <=  gkb  |  tjb  ; 
 olb <=  glb & TJB  |  gcb & tjb  |  GLB & tjb  ; 
 QHD <=  QHJ  |  QHF  ; 
 QHI <=  QHF  |  QHJ  ; 
 OHB <=  GQE & TJJ  |  NDB & JXA  |  ZZO & QGD  ; 
 QHG <= QHB ; 
 nib <= gqh ; 
 ncb <= gcb ; 
 ndk <= gqe ; 
 neb <= gfb ; 
 oza <= hfb ; 
 ozb <= hfb ; 
 ndb <=  gqh & GGG  |  gqb & ggg  ; 
 owh <= gqh ; 
 OXA <= GQA ; 
 OXB <= GQB ; 
 LHA <=  NIA & TIG  |  LGA  ; 
 LHB <=  NIB & TIG  |  LGB  ; 
 LBB <= LAB ; 
 LDB <= LCB ; 
 LEB <= LDB ; 
 LGB <= LFB ; 
 LIB <= LHB ; 
 LJB <= LIB ; 
 LKB <= LJB ; 
 LLB <= LKB ; 
 LOB <= LNB ; 
 LPB <= LOB ; 
 LAB <= IFB ; 
 POA <=  BAF & TCS  |  POA & tcs  ; 
 POB <=  BAF & TCS  |  POA & tcs  ; 
 POC <=  BAF & TCS  |  POA & tcs  ; 
 PKA <=  BBD & bbc & TCS  |  PKA & tcs  ; 
 PKB <=  BBD & bbc & TCS  |  PKA & tcs  ; 
 PKC <=  BBD & bbc & TCS  |  PKA & tcs  ; 
 PGA <=  BBF & bbe & TCK  |  PGA & tck  ; 
 PGB <=  BBF & bbe & TCK  |  PGA & tck  ; 
 PGC <=  BBF & bbe & TCK  |  PGA & tck  ; 
 PCA <=  BBH & bbg & TCK  |  PCA & tck  ; 
 PCB <=  BBH & bbg & TCK  |  PCA & tck  ; 
 PCC <=  BBH & bbg & TCK  |  PCA & tck  ; 
 PGD <=  BCF & bce & TCK  |  PGD & tck  ; 
 PGE <=  BCF & bce & TCK  |  PGD & tck  ; 
 cqc <=  bdc & TCC  |  cqc & tcc  ; 
 cqk <=  bac & TCC  |  cqk & tcc  ; 
 ECC <=  DCB & TEK  |  ECC & tek  ; 
 ECK <=  DGC & TEK  |  ECK & tek  ; 
 edc <=  dfk & TEK  |  edc & tek  ; 
 EDK <=  DGK & TEK  |  EDK & tek  ; 
 EBC <=  DFC & TEK  |  EBC & tek  ; 
 EBK <=  DBJ & TEK  |  EBK & tek  ; 
 EAC <=  DAC & ddc & dak & ZZI & TEC  |  DBC & dak & ZZI & TEC  |  DBK & ZZI & TEC  |  ZZO & TEC  |  EAC & tec  ; 
 EAK <=  DCA & dcc & dck & ddk & TES  |  DEC & dck & ddk & TES  |  DEK & ddk & TES  |  DAS & dda & TES  |  EAK & tes  ; 
 qfa <=  qea & TES  |  qfb & tes  |  QCD  ; 
 qfb <=  qea & TES  |  qfb & tes  |  QCD  ; 
 qfc <=  qea & TES  |  qfb & tes  |  QCD  ; 
 EEC <=  DBS & TEC  |  EEC & tec  ; 
 EQC <=  CQC & TEC  |  EQC & tec  ; 
 EQK <=  CQK & TEC  |  EQK & tec  ; 
 GLC <=  FAC & EAP & THC  |  GLC & thc  ; 
 AAC <=  IAC & JAA  |  AAC & jaa  ; 
 AAK <=  IAK & JAA  |  AAK & jaa  ; 
 ABC <=  IBC & JAB  |  ABC & jab  ; 
 ABK <=  IBK & JAB  |  ABK & jab  ; 
 ACC <=  ICC & JAC  |  ACC & jac  ; 
 ACK <=  ICK & JAC  |  ACK & jac  ; 
 ADC <=  IDC & JAD  |  ADC & jad  ; 
 ADK <=  IDK & JAD  |  ADK & jad  ; 
 RAC <=  JBB & TCC  |  QDC & JBE  |  JBC & tcc  ; 
 RAK <=  JBB & TCC  |  QDC & JBE  |  JBC & tcc  ; 
 RAS <=  JBB & TCC  |  QDC & JBE  |  JBC & tcc  ; 
 gqc <=  eqc & THJ  |  gqc & thj  ; 
 gqk <=  eqk & THJ  |  gqk & thj  ; 
 odd <=  MBA  |  MBB  |  MBC  |  MBD  |  TJS  ; 
 WCB <=  MBA  |  MBB  |  MBC  |  MBD  |  TJS  ; 
 WAE <=  MAA & JWC  |  MAB & JWC  |  MAC & JWC  |  MAD & JWC  |  TJS  ; 
 WAF <=  MAA & JWC  |  MAB & JWC  |  MAC & JWC  |  MAD & JWC  |  TJS  ; 
 GAC <=  FAC & TGA  |  FBC & TGB  |  FCC & TGC  |  GAC & thc  ; 
 GDC <=  FDL & TGQ  |  GDC & tgq  ; 
 GEC <=  FDF & TGQ  |  GEC & tgq  ; 
 GHC <=  ECC & TGS  |  GHC & tgs  ; 
 GIC <=  FEA & TGS  |  GIC & tgs  ; 
 GBC <=  FAC & TGD  |  FBC & TGE  |  FCC & TGF  |  GBC & thc  ; 
 GFC <=  FDS & TGR  |  GFC & tgr  ; 
 GGC <=  EDK & TGR  |  GGC & tgr  ; 
 GJC <=  ECK & TGT  |  GJC & tgt  ; 
 GKC <=  EDC & TGT  |  GKC & tgt  ; 
 GCC <=  FAC & TGG  |  FBC & TGH  |  FCC & TGI  |  GCC & thc  ; 
 LCC <=  TIA & NIC  |  ZZO  |  LBC & LBG  ; 
 LFC <=  TIB & NIC  |  LEC  |  ZZO & LBG  ; 
 LMC <=  TIC & NIC  |  LLC  ; 
 LNC <=  TID & NIC  |  LMC  ; 
 qac <=  jkc & qma  |  jkb & qmb  |  JKA & qmc  ; 
 qbc <=  jlc & qma  |  jlb & qmb  |  JLA & qmc  ; 
 KBC <= KAC ; 
 KCC <= KBC ; 
 KDC <= KCC ; 
 KEC <= KDC ; 
 oac <= eqc ; 
 obc <= eqc ; 
 occ <= eqc ; 
 OWC <= GQC ; 
 KAC <=  NKC & TIE  ; 
 KFC <=  NKG & TIE  |  KEC  ; 
 LQC <=  NLC & TJK  |  LPC  ; 
 LRC <=  LQC & TJK  ; 
 oak <= eqk ; 
 obk <= eqk ; 
 ock <= eqk ; 
 OFC <= LSC ; 
 KIC <=  NKK & TIF  |  KHC  ; 
 KJC <=  NKO & TIF  |  KIC  ; 
 KLC <=  NKS & TJK  |  KKC  ; 
 LSC <=  NLG & TJK  |  LRC  ; 
 KGC <= KFC ; 
 KHC <= KGC ; 
 KKC <= KJC ; 
 OEC <= KLC ; 
 HAC <=  TII & JCC  |  HAC & qac  ; 
 HBC <=  TIJ & JCC  |  HBC & qac  ; 
 oua <=  gjc  |  tjk  ; 
 oub <=  gkc  |  tjk  ; 
 OGC <=  GQC & TJK  |  ZZO & QGC  |  NDL & QGD  ; 
 OHC <=  GQF & TJK  |  NDC & JXA  |  ZZO & QGD  ; 
 HCC <=  NCC & TJC  |  HCC & iec  ; 
 HDC <=  GJC & TJC  |  HDC & iec  ; 
 HFC <=  GGC & TJC  |  JDC & nec  |  IJJ  |  IJK  ; 
 opa <=  gic  |  tjc  ; 
 oqa <=  ghc  |  tjc  ; 
 olc <=  glc & TJC  |  gcc & tjc  |  GLC & tjc  ; 
 hec <= ljg ; 
 OWF <= GQF ; 
 nic <= gqi ; 
 HFI <=  JFC & TJC  |  JDI & qhi  ; 
 OOC <= GQC ; 
 OOF <= GQF ; 
 OWT <= QFA ; 
 nac <= gec ; 
 ncc <= gcc ; 
 ndl <= gqf ; 
 nec <= qmd & ijj ; 
 ndc <=  gqi & GGG  |  gqc & ggg  ; 
 owi <= gqi ; 
 LHC <=  NIC & TIG  |  LGC  ; 
 LBC <= LAC ; 
 LDC <= LCC ; 
 LEC <= LDC ; 
 LGC <= LFC ; 
 LIC <= LHC ; 
 LJC <= LIC ; 
 LKC <= LJC ; 
 LLC <= LKC ; 
 LOC <= LNC ; 
 LPC <= LOC ; 
 LAC <= IFC ; 
 POD <=  BAF & TCT  |  POD & tct  ; 
 POE <=  BAF & TCT  |  POD & tct  ; 
 POF <=  BAF & TCT  |  POD & tct  ; 
 PLA <=  BBD & BAC & TCT  |  PLA & tct  ; 
 PLB <=  BBD & BAC & TCT  |  PLA & tct  ; 
 PLC <=  BBD & BAC & TCT  |  PLA & tct  ; 
 PHA <=  BBF & BBE & TCL  |  PHA & tcl  ; 
 PHB <=  BBF & BBE & TCL  |  PHA & tcl  ; 
 PHC <=  BBF & BBE & TCL  |  PHA & tcl  ; 
 PDA <=  BBH & BBG & TCL  |  PDA & tcl  ; 
 PDB <=  BBH & BBG & TCL  |  PDA & tcl  ; 
 PDC <=  BBH & BBG & TCL  |  PDA & tcl  ; 
 PHD <=  BCF & BCE & TCL  |  PHD & tcl  ; 
 PHE <=  BCF & BCE & TCL  |  PHD & tcl  ; 
 cqd <=  bdd & TCD  |  cqd & tcd  ; 
 cql <=  bad & TCD  |  cql & tcd  ; 
 ECD <=  DBL & TEL  |  ECD & tel  ; 
 ECL <=  DCD & TEL  |  ECL & tel  ; 
 EDD <=  DBE & TEL  |  EDD & tel  ; 
 EDL <=  DCL & TEL  |  EDL & tel  ; 
 EBD <=  DBD & TEL  |  EBD & tel  ; 
 EBL <=  DDL & TEL  |  EBL & tel  ; 
 EAD <=  DCT & ZZI & ZZI & ZZI & TED  |  DAD & ZZI & ZZI & TED  |  DDD & ZZI & TED  |  DAL & TED  |  EAD & ted  ; 
 qfd <=  qea & TED  |  qfb & ted  |  QCD  ; 
 qfe <=  qea & TED  |  qfb & ted  |  QCD  ; 
 qff <=  qea & TED  |  qfb & ted  |  QCD  ; 
 EED <=  DED & TEL  |  EED & tel  ; 
 EEL <=  DEL & TEL  |  EEL & tel  ; 
 EQD <=  CQD & TED  |  EQD & ted  ; 
 EQL <=  CQL & TED  |  EQL & ted  ; 
 GLD <=  FAD & EAP & THD  |  GLD & thd  ; 
 AAD <=  IAD & JAA  |  AAD & jaa  ; 
 AAL <=  IAL & JAA  |  AAL & jaa  ; 
 ABD <=  IBD & JAB  |  ABD & jab  ; 
 ABL <=  IBL & JAB  |  ABL & jab  ; 
 ACD <=  ICD & JAC  |  ACD & jac  ; 
 ACL <=  ICL & JAC  |  ACL & jac  ; 
 ADD <=  IDD & JAD  |  ADD & jad  ; 
 ADL <=  IDL & JAD  |  ADL & jad  ; 
 RAD <=  JBC & TCD  |  QDD & JBE  |  JBD & tcd  ; 
 RAL <=  JBC & TCD  |  QDD & JBE  |  JBD & tcd  ; 
 RAT <=  JBC & TCD  |  QDD & JBE  |  JBD & tcd  ; 
 gqd <=  eqd & THJ  |  gqd & thj  ; 
 gql <=  eql & THJ  |  gql & thj  ; 
 ode <=  MBA  |  MBB  |  MBC  |  MBD  |  TJT  ; 
 WCC <=  MBA  |  MBB  |  MBC  |  MBD  |  TJT  ; 
 WAG <=  MAA & JWD  |  MAB & JWD  |  MAC & JWD  |  MAD & JWD  |  TJT  ; 
 WAH <=  MAA & JWD  |  MAB & JWD  |  MAC & JWD  |  MAD & JWD  |  TJT  ; 
 GAD <=  FAD & TGA  |  FBD & TGB  |  FCD & TGC  |  GAD & thd  ; 
 GDD <=  FDM & TGQ  |  GDD & tgq  ; 
 GED <=  FDG & TGQ  |  GED & tgq  ; 
 GHD <=  ECL & TGS  |  GHD & tgs  ; 
 GID <=  EBL & TGS  |  GID & tgs  ; 
 GBD <=  FAD & TGD  |  FBD & TGE  |  FCD & TGF  |  GBD & thd  ; 
 GFD <=  EBM & TGR  |  GFD & tgr  ; 
 GGD <=  EBD & TGR  |  GGD & tgr  ; 
 GJD <=  FDO & TGT  |  GJD & tgt  ; 
 GKD <=  EDD & TGT  |  GKD & tgt  ; 
 GCD <=  FAD & TGG  |  FBD & TGH  |  FCD & TGI  |  GCD & thd  ; 
 LCD <=  TIA & ZZI  |  LBG  ; 
 LMD <=  TIC & ZZI  |  LLD  ; 
 NKA <= JGA & GQG ; 
 NKB <= JGA & GQH ; 
 NKC <= JGA & GQI ; 
 NKD <= JGA & ZZI ; 
 qad <=  jkc & qma  |  jkb & qmb  |  jka & qmc  ; 
 qbd <=  jlc & qma  |  jlb & qmb  |  jla & qmc  ; 
 KBD <= KAD ; 
 KCD <= KBD ; 
 KDD <= KCD ; 
 KED <= KDD ; 
 oad <= eqd ; 
 obd <= eqd ; 
 ocd <= eqd ; 
 owj <= gqj ; 
 KAD <=  NKD & TIE  ; 
 KFD <=  JKE & TIE  |  KED  ; 
 LQD <=  JLE & TJL  |  LPD  ; 
 LRD <=  LQD & TJL  ; 
 oal <= eql ; 
 obl <= eql ; 
 ocl <= eql ; 
 OFD <= LSD ; 
 KID <=  ZZO & TIF  |  KHD  ; 
 KJD <=  NKP & TIF  |  KID  ; 
 KLD <=  JKH & TJL  |  KKD  ; 
 LSD <=  NLH & TJL  |  LRD  ; 
 KGD <= KFD ; 
 KHD <= KGD ; 
 KKD <= KJD ; 
 OED <= KLD ; 
 HAD <=  TII & JCD  |  HAD & qad  ; 
 HBD <=  TIJ & JCD  |  HBD & qad  ; 
 ova <=  gkd  |  tjl  ; 
 qge <=  ged  |  tjl  ; 
 QGC <=  JPA & TJL  ; 
 OHD <=  NDD & TJL  |  NDG & QGC  ; 
 HCD <=  NCD & TJD  |  HCD & ied  ; 
 HDD <=  GJD & TJD  |  HDD & ied  ; 
 hed <=  lkg  ; 
 HFD <=  qca  |  qee  ; 
 QJA <=  GGD & TJD  ; 
 OTC <=  GHD & TJD  ; 
 old <=  gld & TJD  |  gcd & tjd  |  GLD & tjd  ; 
 OSD <=  GHH & TJD  ; 
 OJD <= QJA ; 
 OTG <= JOC ; 
 OUE <= JOC ; 
 nad <= ged ; 
 ncd <= gcd ; 
 ndd <= jma ; 
 LFD <=  TIB & GQL  |  LED  ; 
 ndg <=  jmd & jme & JNA  |  nia & jna  ; 
 owk <= gqk ; 
 owl <= gql ; 
 LND <=  TID & nee  |  LMD  ; 
 LDD <= LCD ; 
 LED <= LDD ; 
 LGD <= LFD ; 
 LHD <= LGD ; 
 LID <= LHD ; 
 LJD <= LID ; 
 LKD <= LJD ; 
 LLD <= LKD ; 
 LOD <= LND ; 
 LPD <= LOD ; 
 PNA <=  BAD & TCU  |  PNA & tcu  ; 
 PNB <=  BAD & TCU  |  PNA & tcu  ; 
 PNC <=  BAD & TCU  |  PNA & tcu  ; 
 PID <=  bcd & bcc & TCU  |  PID & tcu  ; 
 PIE <=  bcd & bcc & TCU  |  PID & tcu  ; 
 PEF <=  bbf & bbe & TCM  |  PEF & tcm  ; 
 PAD <=  bbh & bbg & TCM  |  PAD & tcm  ; 
 PAE <=  bbh & bbg & TCM  |  PAD & tcm  ; 
 PAF <=  bbh & bbg & TCM  |  PAD & tcm  ; 
 PAG <=  bch & bcg & TCM  |  PAG & tcm  ; 
 PAH <=  bch & bcg & TCM  |  PAG & tcm  ; 
 cqe <=  bde & TCE  |  cqe & tce  ; 
 cqm <=  bae & TCE  |  cqm & tce  ; 
 ECE <=  DCK & TEM  |  ECE & tem  ; 
 ECM <=  DCM & TEM  |  ECM & tem  ; 
 ede <=  dfm & TEM  |  DDA & TEM  |  ede & tem  ; 
 EDM <=  DBT & TEM  |  ZZO & TEM  |  EDM & tem  ; 
 EBE <=  DDM & TEM  |  EBE & tem  ; 
 EBM <=  DFE & TEM  |  EBM & tem  ; 
 EAE <=  DAU & dek & dde & ddd & TEE  |  DCE & dde & ddd & TEE  |  DCW & ddd & TEE  |  DCU & def & TEE  |  EAE & tee  ; 
 EAM <=  DBU & dfd & dam & dbe & TEE  |  DEE & dam & dbe & TEE  |  ZZO & dbe & TEE  |  DCV & dem & TEE  |  EAM & tee  ; 
 qea <=  jaf & TCE  |  qea & tce  |  QCD  ; 
 qeb <=  jaf & TCE  |  qea & tce  |  QCD  ; 
 qec <=  jaf & TCE  |  qea & tce  |  QCD  ; 
 EEE <=  DGE & TEE  |  EEE & tee  ; 
 EEM <=  DGM & TEE  |  EEM & tee  ; 
 EQE <=  CQE & TEE  |  EQE & tee  ; 
 EQM <=  CQM & TEE  |  EQM & tee  ; 
 GLE <=  FAE & EAP & THE  |  GLE & the  ; 
 AAE <=  IAE & JAH  |  AAE & jah  ; 
 AAM <=  IAM & JAH  |  AAM & jah  ; 
 ABE <=  IBE & JAG  |  ABE & jag  ; 
 ABM <=  IBM & JAG  |  ABM & jag  ; 
 ACE <=  ICE & JAC  |  ACE & jac  ; 
 ACM <=  ICM & JAC  |  ACM & jac  ; 
 ADE <=  IDE & JAD  |  ADE & jad  ; 
 ADM <=  IDM & JAD  |  ADM & jad  ; 
 RAE <=  JAE & jbe  |  QDA & JBE  |  JBA & tce  ; 
 RAM <=  JAE & jbe  |  QDA & JBE  |  JBA & tce  ; 
 RAU <=  JAE & jbe  |  QDA & JBE  |  JBA & tce  ; 
 gqe <=  eqe & THK  |  gqe & thk  ; 
 gqm <=  eqm & THK  |  gqm & thk  ; 
 odf <=  MBE  |  MBF  |  MBG  |  MBH  |  QGB  ; 
 WDA <=  MBE  |  MBF  |  MBG  |  MBH  |  QGB  ; 
 WBA <=  MAE & JWE  |  MAF & JWE  |  MAG & JWE  |  MAH & JWE  ; 
 WBB <=  MAE & JWE  |  MAF & JWE  |  MAG & JWE  |  MAH & JWE  ; 
 GAE <=  FAE & TGA  |  FBE & TGB  |  FCE & TGC  |  GAE & the  ; 
 GDE <=  FDY & TGQ  |  GDE & tgq  ; 
 GEE <=  FDH & TGQ  |  GEE & tgq  ; 
 GHE <=  FDB & TGS  |  GHE & tgs  ; 
 GIE <=  ECM & TGS  |  GIE & tgs  ; 
 GBE <=  FAE & TGD  |  FBE & TGE  |  FCE & TGF  |  GBE & the  ; 
 GFE <=  FDT & TGR  |  GFE & tgr  ; 
 GGE <=  FDE & TGR  |  GGE & tgr  ; 
 GJE <=  FDV & TGT  |  GJE & tgt  ; 
 GKE <=  EBI & TGT  |  GKE & tgt  ; 
 GCE <=  FAE & TGG  |  FBE & TGH  |  FCE & TGI  |  GCE & the  ; 
 LCE <=  LBG  ; 
 LFE <=  LEE  ; 
 LME <=  TIC & ZZI  |  LLE  ; 
 LNE <=  TID & ZZI  |  LME  ; 
 NKE <= JGB & GQG ; 
 NKF <= JGB & GQH ; 
 NKG <= JGB & GQI ; 
 NKH <= JGB & ZZI ; 
 qae <=  jkd & qma  |  JKB & qmb  |  JKA & qmc  ; 
 qbe <=  jld & qma  |  JLB & qmb  |  JLA & qmc  ; 
 oae <= eqe ; 
 obe <= eqe ; 
 oce <= eqe ; 
 OWM <= GQM ; 
 KFE <=  JKF & TIE  ; 
 LQE <=  JLF & TJM  |  LPE  ; 
 LRE <=  LQE & TJM  ; 
 oam <= eqm ; 
 obm <= eqm ; 
 ocm <= eqm ; 
 OFE <= LSE ; 
 KIE <=  NKL & TIF  |  KHE  ; 
 KJE <=  NKP & TIF  |  KIE  ; 
 KLE <=  KKE  ; 
 LSE <=  LRE  ; 
 KGE <= KFE ; 
 KHE <= KGE ; 
 KKE <= KJE ; 
 OEE <= KLE ; 
 HAE <=  TII & JCE  |  HAE & qae  ; 
 HBE <=  TIJ & JCE  |  HBE & qae  ; 
 OVB <=  GKE & TJM  ; 
 OHE <=  NDE & TJM  |  NDH & QGC  ; 
 HCE <=  NCE & TJE  |  HCE & iee  ; 
 HDE <=  KCG & TJE  ; 
 hee <=  lng  ; 
 HFE <=  qee  |  jaf  ; 
 oja <=  tje  |  ggb  |  jnb  ; 
 ojb <=  tje  |  ggb  ; 
 ole <=  gle & TJE  |  gce & tje  |  GLE & tje  ; 
 OMA <=  gih & TJE  |  ggc & tje  ; 
 nce <= gce ; 
 nde <= jmb ; 
 ndh <=  JMD & JNA  |  nib & jna  ; 
 LDE <= LCE ; 
 LEE <= LDE ; 
 LGE <= LFE ; 
 LHE <= LGE ; 
 LIE <= LHE ; 
 LJE <= LIE ; 
 LKE <= LJE ; 
 LLE <= LKE ; 
 LOE <= LNE ; 
 LPE <= LOE ; 
 owu <= ram ; 
 PND <=  BAD & TCV  |  PND & tcv  ; 
 PNE <=  BAD & TCV  |  PND & tcv  ; 
 PNF <=  BAD & TCV  |  PND & tcv  ; 
 PJD <=  bcd & BBC & TCV  |  PJD & tcv  ; 
 PJE <=  bcd & BBC & TCV  |  PJD & tcv  ; 
 PJF <=  bcd & BBC & TCV  |  PJD & tcv  ; 
 PFF <=  bbf & BBE & TCN  |  PFF & tcn  ; 
 PFG <=  bbf & BBE & TCN  |  PFF & tcn  ; 
 PFH <=  bbf & BBE & TCN  |  PFF & tcn  ; 
 PBD <=  bbh & BBG & TCN  |  PBD & tcn  ; 
 PBE <=  bbh & BBG & TCN  |  PBD & tcn  ; 
 PBF <=  bbh & BBG & TCN  |  PBD & tcn  ; 
 PBG <=  bch & BCG & TCN  |  PBG & tcn  ; 
 PBH <=  bch & BCG & TCN  |  PBG & tcn  ; 
 cqf <=  bdf & TCF  |  cqf & tcf  ; 
 cqn <=  baf & TCF  |  cqn & tcf  ; 
 ECF <=  DCF & TEN  |  ZZO & TEN  |  ECF & ten  ; 
 ecn <=  dan & TEN  |  DFE & TEN  |  ecn & ten  ; 
 EDF <=  DCN & TEN  |  EDF & ten  ; 
 EDN <=  DFF & TEN  |  EDN & ten  ; 
 EBF <=  DDF & TEN  |  EBF & ten  ; 
 EBN <=  DBN & TEN  |  EBN & ten  ; 
 EAF <=  daf & dav & dbp & ZZI & TEF  |  ZZO & dbp & ZZI & TEF  |  ZZO & ZZI & TEF  |  ZZO & TEF  |  EAF & tef  ; 
 EAN <=  DAN & ZZI & ZZI & ZZI & TEF  |  DDN & ZZI & ZZI & TEF  |  DBV & ZZI & TEF  |  DBF & TEF  |  EAN & tef  ; 
 qed <=  jaf & TCF  |  qea & tcf  |  QCD  ; 
 qee <=  jaf & TCF  |  qea & tcf  |  QCD  ; 
 EEF <=  DFN & TEF  |  EEF & tef  ; 
 EEN <=  DAN & TEF  |  EEN & tef  ; 
 EQF <=  CQF & TEF  |  EQF & tef  ; 
 EQN <=  CQN & TEF  |  EQN & tef  ; 
 GLF <=  FAF & EAP & THF  |  GLF & thf  ; 
 EEG <=  DEN & TEF  |  EEG & tef  ; 
 AAF <=  IAF & JAH  |  AAF & jah  ; 
 AAN <=  IAN & JAH  |  AAN & jah  ; 
 ABF <=  IBF & JAG  |  ABF & jag  ; 
 ABN <=  IBN & JAG  |  ABN & jag  ; 
 ACF <=  ICF & JAC  |  ACF & jac  ; 
 ACN <=  ICN & JAC  |  ACN & jac  ; 
 ADF <=  IDF & JAD  |  ADF & jad  ; 
 ADN <=  IDN & JAD  |  ADN & jad  ; 
 RAF <=  JBA & TCF  |  QDB & JBE  |  JBB & tcf  ; 
 RAN <=  JBA & TCF  |  QDB & JBE  |  JBB & tcf  ; 
 RAV <=  JBA & TCF  |  QDB & JBE  |  JBB & tcf  ; 
 gqf <=  eqf & THK  |  gqf & thk  ; 
 gqn <=  eqn & THK  |  gqn & thk  ; 
 odg <=  MBE  |  MBF  |  MBG  |  MBH  |  QGB  ; 
 WDB <=  MBE  |  MBF  |  MBG  |  MBH  |  QGB  ; 
 WBC <=  MAE & JWF  |  MAF & JWF  |  MAG & JWF  |  MAH & JWF  ; 
 WBD <=  MAE & JWF  |  MAF & JWF  |  MAG & JWF  |  MAH & JWF  ; 
 GAF <=  FAF & TGA  |  FBF & TGB  |  FCF & TGC  |  GAF & thf  ; 
 GDF <=  FDC & TGQ  |  GDF & tgq  ; 
 GEF <=  FDI & TGQ  |  GEF & tgq  ; 
 GHF <=  FDA & TGS  |  GHF & tgs  ; 
 GIF <=  FDX & TGS  |  GIF & tgs  ; 
 GBF <=  FAF & TGD  |  FBF & TGE  |  FCF & TGF  |  GBF & thf  ; 
 GFF <=  FDU & TGR  |  GFF & tgr  ; 
 GGF <=  EBF & TGR  |  GGF & tgr  ; 
 GJF <=  FDW & TGT  |  GJF & tgt  ; 
 GKF <=  EDL & TGT  |  GKF & tgt  ; 
 GCF <=  FAF & TGG  |  FBF & TGH  |  FCF & TGI  |  GCF & thf  ; 
 LCF <=  TIA & ZZI  ; 
 LFF <=  TIB & ZZI  |  LEF  ; 
 LMF <=  TIC & ZZI  |  LLF  ; 
 NKI <= JGC & GQG ; 
 NKJ <= JGC & GQH ; 
 NKK <= JGC & GQI ; 
 NKL <= JGC & ZZI ; 
 qaf <=  jkd & qma  |  JKB & qmb  |  jka & qmc  ; 
 qbf <=  jld & qma  |  JLB & qmb  |  jla & qmc  ; 
 KBF <= KAF ; 
 KCF <= KBF ; 
 KDF <= KCF ; 
 KEF <= KDF ; 
 oaf <= eqf ; 
 obf <= eqf ; 
 ocf <= eqf ; 
 OWN <= GQN ; 
 KAF <=  NKD & TIE  ; 
 KFF <=  JKE & TIE  |  KEF  ; 
 LQF <=  JLG & TJN  |  LPF  ; 
 LRF <=  LQF & TJN  ; 
 oan <= eqn ; 
 obn <= eqn ; 
 ocn <= eqn ; 
 OFF <= LSF ; 
 KIF <=  JKG & TIF  |  KHF  ; 
 KJF <=  KIF & TIF  ; 
 KLF <=  JKI & TJN  |  KKF  ; 
 LSF <=  LRF & TJN  ; 
 KGF <= KFF ; 
 KHF <= KGF ; 
 KKF <= KJF ; 
 OEF <= KLF ; 
 HAF <=  TII & JCF  |  HAF & qaf  ; 
 HBF <=  TIJ & JCF  |  HBF & qaf  ; 
 OVC <=  GKF & TJN  ; 
 OHF <=  NDF & TJN  |  NDI & QGC  ; 
 HCF <=  NCF & TJF  |  HCF & ief  ; 
 HDF <=  KFG & TJF  ; 
 hef <=  lpg & nld  |  lpg & tjf  ; 
 HFF <=  qee & nld  ; 
 QIA <=  GJF & TJF  ; 
 QIB <=  GJG & TJF  ; 
 olf <=  glf & TJF  |  gcf & tjf  |  GLF & tjf  ; 
 OMB <=  gih & TJF  |  ggc & tjf  ; 
 QIC <= QIB ; 
 QID <= QIC ; 
 qie <= qcd ; 
 onb <= gif ; 
 OWS <= QEE ; 
 ncf <= gcf ; 
 ndf <= jmc ; 
 ndi <=  jmf & ZZI & JNA  |  nic & jna  ; 
 LNF <=  TID & nee  |  LMF  ; 
 LDF <= LCF ; 
 LEF <= LDF ; 
 LGF <= LFF ; 
 LIF <= LHF ; 
 LJF <= LIF ; 
 LKF <= LJF ; 
 LLF <= LKF ; 
 LOF <= LNF ; 
 LPF <= LOF ; 
 owv <= ran ; 
 PMA <=  BBB & TCW  |  PMA & tcw  ; 
 PMB <=  BBB & TCW  |  PMA & tcw  ; 
 PMC <=  BBB & TCW  |  PMA & tcw  ; 
 PKD <=  BCD & bcc & TCW  |  PKD & tcw  ; 
 PKE <=  BCD & bcc & TCW  |  PKD & tcw  ; 
 PKF <=  BCD & bcc & TCW  |  PKD & tcw  ; 
 PGF <=  BBF & bbe & TCO  |  PGF & tco  ; 
 PGG <=  BBF & bbe & TCO  |  PGF & tco  ; 
 PCD <=  BBH & bbg & TCO  |  PCD & tco  ; 
 PCE <=  BBH & bbg & TCO  |  PCD & tco  ; 
 PCF <=  BBH & bbg & TCO  |  PCD & tco  ; 
 PCG <=  BCH & bcg & TCO  |  PCG & tco  ; 
 cqg <=  bdg & TCG  |  cqg & tcg  ; 
 cqo <=  bag & TCG  |  cqo & tcg  ; 
 ECG <=  DBG & TEO  |  ECG & teo  ; 
 ECO <=  DBM & TEO  |  ECO & teo  ; 
 EDG <=  DDO & TEO  |  EDG & teo  ; 
 EDO <=  DFG & TEO  |  EDO & teo  ; 
 EBG <=  DDG & TEO  |  EBG & teo  ; 
 EAG <=  DAW & dag & ZZI & ZZI & TEG  |  ZZO & ZZI & ZZI & TEG  |  ZZO & ZZI & TEG  |  ZZO & TEG  |  EAG & teg  ; 
 EQG <=  CQG & TEG  |  EQG & teg  ; 
 EQO <=  CQO & TEG  |  EQO & teg  ; 
 GLG <=  FAG & EAP & THG  |  GLG & thg  ; 
 AAG <=  IAG & JAH  |  AAG & jah  ; 
 AAO <=  IAO & JAH  |  AAO & jah  ; 
 ABG <=  IBG & JAG  |  ABG & jag  ; 
 ABO <=  IBO & JAG  |  ABO & jag  ; 
 ACG <=  ICG & JAC  |  ACG & jac  ; 
 ACO <=  ICO & JAC  |  ACO & jac  ; 
 ADG <=  IDG & JAD  |  ADG & jad  ; 
 ADO <=  IDO & JAD  |  ADO & jad  ; 
 RAG <=  JBB & TCG  |  QDC & JBE  |  JBC & tcg  ; 
 RAO <=  JBB & TCG  |  QDC & JBE  |  JBC & tcg  ; 
 RAW <=  JBB & TCG  |  QDC & JBE  |  JBC & tcg  ; 
 QCD <=  QCD & qca  |  IKB  ; 
 QCE <=  QCD & qca  |  IKB  ; 
 gqg <=  eqg & THL  |  gqg & thl  ; 
 gqo <=  eqo & THL  |  gqo & thl  ; 
 odh <=  MBE  |  MBF  |  MBG  |  MBH  |  QGB  ; 
 WDC <=  MBE  |  MBF  |  MBG  |  MBH  |  QGB  ; 
 WBE <=  MAE & JWG  |  MAF & JWG  |  MAG & JWG  |  MAH & JWG  ; 
 WBF <=  MAE & JWG  |  MAF & JWG  |  MAG & JWG  |  MAH & JWG  ; 
 nei <= gfi ; 
 nku <= jgd ; 
 GAG <=  FAG & TGA  |  FBG & TGB  |  FCG & TGC  |  GAG & thg  ; 
 GDG <=  EBG & TGQ  |  GDG & tgq  ; 
 GEG <=  EDC & TGQ  |  GEG & tgq  ; 
 GHG <=  ECO & TGS  |  GHG & tgs  ; 
 GIG <=  EEJ & TGS  |  GIG & tgs  ; 
 GBG <=  FAG & TGD  |  FBG & TGE  |  FCG & TGF  |  GBG & thg  ; 
 GFI <=  FDZ & TGR  |  GFI & tgr  ; 
 GGG <=  FDQ & TGR  |  GGG & tgr  ; 
 GJG <=  EBM & TGT  |  GJG & tgt  ; 
 GKG <=  EED & TGT  |  GKG & tgt  ; 
 GCG <=  FAG & TGG  |  FBG & TGH  |  FCG & TGI  |  GCG & thg  ; 
 LCG <=  TIA & ZZI  |  LBG  ; 
 LFG <=  TIB & ZZI  |  LEG  ; 
 LMG <=  TIC & ZZI  |  LLG  ; 
 LNG <=  TID & ZZI  |  LMG  ; 
 NKM <= JGD & GQG ; 
 NKN <= JGD & GQH ; 
 NKO <= JGD & GQI ; 
 NKP <= JGD & ZZI ; 
 qag <=  jkd & qma  |  jkb & qmb  |  JKA & qmc  ; 
 qbg <=  jld & qma  |  jlb & qmb  |  JLA & qmc  ; 
 KBG <= KAG ; 
 KCG <= KBG ; 
 KDG <= KCG ; 
 KEG <= KDG ; 
 oag <= eqg ; 
 obg <= eqg ; 
 ocg <= eqg ; 
 OWO <= GQO ; 
 KAG <=  NKD & TIE  ; 
 KFG <=  NKH & TIE  |  KEG  ; 
 LQG <=  NLD & TJO  |  LPG  ; 
 oao <= eqo ; 
 obo <= eqo ; 
 oco <= eqo ; 
 KIG <=  NKL & TIF  |  KHG  ; 
 KJG <=  NKP & TIF  |  KIG  ; 
 KGG <= KFG ; 
 KHG <= KGG ; 
 HAG <=  TII & JCG  |  HAG & qag  ; 
 HBG <=  TIJ & JCG  |  HBG & qag  ; 
 OVD <=  GKG & TJO  ; 
 OHG <=  GGH & TJO  ; 
 HCG <=  NCG & TJG  |  HCG & ieg  ; 
 HDG <=  KGG & TJG  ; 
 HFG <=  GIG & TJG  |  IKC  |  qka & HFG  ; 
 ojc <=  tjg  |  ghg  ; 
 owr <=  tjg  ; 
 olg <=  glg & TJG  |  gcg & tjg  |  GLG & tjg  ; 
 ORD <=  GIH & TJG  ; 
 NAG <=  GEG & yyy  ; 
 nab <=  GEG & yyy  |  geb  ; 
 qka <= ikc ; 
 qkb <= ila ; 
 ncg <= gcg ; 
 OTE <= JOA ; 
 OUC <= JOA ; 
 OVE <= JOA ; 
 OPB <= JOA ; 
 OQB <= JOA ; 
 ORB <= JOA ; 
 OSB <= JOA ; 
 LHF <=  TIG  |  LGF  ; 
 LHG <=  TIG  |  LGG  ; 
 lbg <= hea ; 
 LDG <= LCG ; 
 LEG <= LDG ; 
 LGG <= LFG ; 
 LIG <= LHG ; 
 LJG <= LIG ; 
 LKG <= LJG ; 
 LLG <= LKG ; 
 LOG <= LNG ; 
 LPG <= LOG ; 
 oww <= rao ; 
 PMD <=  BBB & TCX  |  PMD & tcx  ; 
 PME <=  BBB & TCX  |  PMD & tcx  ; 
 PMF <=  BBB & TCX  |  PMD & tcx  ; 
 PLD <=  BCD & BBC & TCX  |  PLD & tcx  ; 
 PLE <=  BCD & BBC & TCX  |  PLD & tcx  ; 
 PLF <=  BCD & BBC & TCX  |  PLD & tcx  ; 
 PHF <=  BBF & BBE & TCP  |  PHF & tcp  ; 
 PHG <=  BBF & BBE & TCP  |  PHF & tcp  ; 
 PHH <=  BBF & BBE & TCP  |  PHF & tcp  ; 
 PDD <=  BBH & BBG & TCP  |  PDD & tcp  ; 
 PDE <=  BBH & BBG & TCP  |  PDD & tcp  ; 
 PDF <=  BBH & BBG & TCP  |  PDD & tcp  ; 
 PDG <=  BCH & BCG & TCP  |  PDG & tcp  ; 
 PDH <=  BCH & BCG & TCP  |  PDG & tcp  ; 
 cqh <=  bdh & TCH  |  cqh & tch  ; 
 cqp <=  bah & TCH  |  cqp & tch  ; 
 EDH <=  DBP & TEP  |  EDH & tep  ; 
 EDP <=  DDP & TEP  |  EDP & tep  ; 
 EAH <=  DAW & dah & dci & ZZI & TEH  |  DAP & dci & ZZI & TEH  |  DEM & ZZI & TEH  |  DBH & dci & TEH  |  EAH & teh  ; 
 EAP <=  DAT & ZZI & ZZI & ZZI & TEH  |  DDH & ZZI & ZZI & TEH  |  ZZO & ZZI & TEH  |  ZZO & TEH  |  EAP & teh  ; 
 EQH <=  CQH & TEH  |  EQH & teh  ; 
 EQP <=  CQP & TEH  |  EQP & teh  ; 
 GLH <=  FAH & EAP & THH  |  GLH & thh  ; 
 AAH <=  IAH & JAH  |  AAH & jah  ; 
 AAP <=  IAP & JAH  |  AAP & jah  ; 
 ABH <=  IBH & JAG  |  ABH & jag  ; 
 ABP <=  IBP & JAG  |  ABP & jag  ; 
 ACH <=  ICH & JAC  |  ACH & jac  ; 
 ACP <=  ICP & JAC  |  ACP & jac  ; 
 ADH <=  IDH & JAD  |  ADH & jad  ; 
 ADP <=  IDP & JAD  |  ADP & jad  ; 
 RAH <=  JBC & TCH  |  QDD & JBE  |  JBD & tch  ; 
 RAP <=  JBC & TCH  |  QDD & JBE  |  JBD & tch  ; 
 RAX <=  JBC & TCH  |  QDD & JBE  |  JBD & tch  ; 
 QCA <=  QCA & jae & ikb  |  IKA  ; 
 QCB <=  QCA & jae & ikb  |  IKA  ; 
 QCC <=  QCA & jae & ikb  |  IKA  ; 
 gqh <=  eqh & THL  |  gqh & thl  ; 
 gqp <=  eqp & THL  |  gqp & thl  ; 
 odi <=  MBE  |  MBF  |  MBG  |  MBH  |  QGB  ; 
 odj <=  MBE  |  MBF  |  MBG  |  MBH  |  QGB  ; 
 WBG <=  MAE & JWH  |  MAF & JWH  |  MAG & JWH  |  MAH & JWH  ; 
 WBH <=  MAE & JWH  |  MAF & JWH  |  MAG & JWH  |  MAH & JWH  ; 
 GAH <=  FAH & TGA  |  FBH & TGB  |  FCH & TGC  |  GAH & thh  ; 
 GDH <=  FDD & TGQ  |  GDH & tgq  ; 
 GHH <=  EEL & TGS  |  GHH & tgs  ; 
 GIH <=  EDH & TGS  |  GIH & tgs  ; 
 GBH <=  FAH & TGD  |  FBH & TGE  |  FCH & TGF  |  GBH & thh  ; 
 GGH <=  FDP & TGR  |  GGH & tgr  ; 
 GJH <=  EDP & TGT  |  GJH & tgt  ; 
 GCH <=  FAH & TGG  |  FBH & TGH  |  FCH & TGI  |  GCH & thh  ; 
 NKQ <= JGE & GQG ; 
 NKR <= JGE & GQH ; 
 NKS <= JGE & GQI ; 
 NKT <= JGE & ZZI ; 
 qah <=  jkd & qma  |  jkb & qmb  |  jka & qmc  ; 
 qbh <=  jld & qma  |  jlb & qmb  |  jla & qmc  ; 
 QMA <= IKQ ; 
 QMB <= IKQ ; 
 QMC <= IKQ ; 
 QMD <= IKQ ; 
 oah <= eqh ; 
 obh <= eqh ; 
 och <= eqh ; 
 oap <= eqp ; 
 obp <= eqp ; 
 ocp <= eqp ; 
 qda <=  IGB  |  IGA  ; 
 qdb <=  IGB  |  iga  ; 
 qdc <=  igb  |  IGA  ; 
 qdd <=  igb  |  iga  ; 
 oka <= jae ; 
 HAH <=  TII & JCH  |  HAH & qah  ; 
 HBH <=  TIJ & JCH  |  HBH & qah  ; 
 QLA <=  GHG & TJP  ; 
 QLB <=  QLA & TJP  ; 
 QLC <= QLB ; 
 HCH <=  NCH & TJH  |  HCH & ieh  ; 
 HDH <=  NKU & TJH  |  KIG & ieh  ; 
 HFH <=  GHG & TJP  |  QLA  |  QLB  |  QGA  |  QLC  ; 
 QGA <=  qfa & qga & THM  |  GJE & TJH  |  JFD  ; 
 QGB <=  qfa & qga & THM  |  GJE & TJH  |  JFD  ; 
 olh <=  glh & TJH  |  gch & tjh  |  GLH & tjh  ; 
 OXC <=  GJH & TJH  |  ZZO & tjh  |  ZZO & tjh  ; 
 OIA <= THM ; 
 OIB <= THM ; 
 owp <= gqp ; 
 OWQ <= THM ; 
 nee <= jgi ; 
 nch <= gch ; 
 OTF <= JOB ; 
 OUD <= JOB ; 
 OVF <= JOB ; 
 owx <= rap ; 
 OPC <= JOB ; 
 OQC <= JOB ; 
 ORC <= JOB ; 
 OSC <= JOB ; 
 end 
endmodule;
