module me( IZZ,
 IAB, 
 IAC, 
 IAD, 
 IAE, 
 IAF, 
 IAG, 
 IAH, 
 IAI, 
 IAJ, 
 IAK, 
 IAL, 
 IAM, 
 IAN, 
 IAO, 
 IAP, 
 IAQ, 
 IAR, 
 IAS, 
 IAT, 
 IAU, 
 IAV, 
 IAW, 
 IAX, 
 IAY, 
 IAZ, 
 IBA, 
 IBB, 
 IBC, 
 IBD, 
 IBE, 
 IBF, 
 IBG, 
 IBH, 
 IBI, 
 IBJ, 
 IBK, 
 IBL, 
 IBM, 
 IBN, 
 IBO, 
 IBP, 
 IBQ, 
 IBR, 
 IBS, 
 IBT, 
 IBU, 
 IBV, 
 IBW, 
 IBX, 
 IBY, 
 IBZ, 
 ICB, 
 ICC, 
 ICD, 
 ICE, 
 ICF, 
 ICG, 
 ICH, 
 ICI, 
 ICK, 
 ICL, 
 ICM, 
 ICN, 
 ICO, 
 ICP, 
 ICQ, 
 ICS, 
 ICT, 
 ICU, 
 ICV, 
 ICW, 
 ICX, 
 ICY, 
 ICZ, 
 IDA, 
 IDB, 
 IDC, 
 IDD, 
 IDE, 
 IDF, 
 IDG, 
 IDH, 
 IDI, 
 IDJ, 
 IDK, 
 IDL, 
 IDM, 
 IDN, 
 IDO, 
 IDP, 
 IDQ, 
 IDR, 
 IDS, 
 IDT, 
 IDU, 
 IDV, 
 IDW, 
 IDX, 
 IDY, 
 IDZ, 
 IEF, 
 IEG, 
 IEH, 
 IEI, 
 IEO, 
 IEP, 
 IEQ, 
 IFFF , 
 IFO, 
 IGA, 
 IGB, 
 IGC, 
 IGD, 
 IGE, 
 IGF, 
 IGG, 
 IGH, 
 IGI, 
 IGJ, 
 IGK, 
 IGL, 
 IGM, 
 IGN, 
 IGO, 
 IGP, 
 IHA, 
 IHB, 
 IHC, 
 IHD, 
 IHE, 
 IHF, 
 IHG, 
 IHH, 
 IHI, 
 IHJ, 
 IHK, 
 IHL, 
 IHM, 
 IHN, 
 IHO, 
 IHP, 
 IUA, 
 IUB, 
 IVA, 
 IVB, 
 IVC, 
 IVD, 
 IVE, 
 IVF, 
 OAA, 
 OAB, 
 OAC, 
 OAD, 
 OAE, 
 OAF, 
 OAG, 
 OAH, 
 OAI, 
 OAJ, 
 OAK, 
 OAL, 
 OAM, 
 OAN, 
 OAO, 
 OAP, 
 OAQ, 
 OAR, 
 OAS, 
 OAT, 
 OAU, 
 OAV, 
 OAW, 
 OAX, 
 OBA, 
 OBB, 
 OBC, 
 OBD, 
 OBE, 
 OBF, 
 OBG, 
 OBH, 
 OBI, 
 OBJ, 
 OBK, 
 OBL, 
 OBM, 
 OBN, 
 OBO, 
 OBP, 
 OBQ, 
 OBR, 
 OBS, 
 OBT, 
 OBU, 
 OBV, 
 OBW, 
 OBX, 
 OCA, 
 OCB, 
 OCC, 
 OCD, 
 OCE, 
 OCF, 
 OCG, 
 OCH, 
 OCI, 
 OCJ, 
 OCK, 
 OCL, 
 OCM, 
 OCN, 
 OCO, 
 OCP, 
 ODA, 
 ODB, 
 ODC, 
 OEA, 
 OEB, 
 OEC, 
 OFA, 
 OFB, 
 OFC, 
 OGA, 
 OGB, 
 OGC, 
 OHA, 
 OHB, 
 OHC, 
 OIA, 
 OIB, 
 OIC, 
 OID, 
 OJA, 
 OJB, 
 OJC, 
 OJD, 
 OJE, 
 OJF, 
 OKA, 
 OLA, 
 OMA, 
 OMB, 
 OMC, 
OMD ); 
    
 input IZZ; 
 input IAB; 
 input IAC; 
 input IAD; 
 input IAE; 
 input IAF; 
 input IAG; 
 input IAH; 
 input IAI; 
 input IAJ; 
 input IAK; 
 input IAL; 
 input IAM; 
 input IAN; 
 input IAO; 
 input IAP; 
 input IAQ; 
 input IAR; 
 input IAS; 
 input IAT; 
 input IAU; 
 input IAV; 
 input IAW; 
 input IAX; 
 input IAY; 
 input IAZ; 
 input IBA; 
 input IBB; 
 input IBC; 
 input IBD; 
 input IBE; 
 input IBF; 
 input IBG; 
 input IBH; 
 input IBI; 
 input IBJ; 
 input IBK; 
 input IBL; 
 input IBM; 
 input IBN; 
 input IBO; 
 input IBP; 
 input IBQ; 
 input IBR; 
 input IBS; 
 input IBT; 
 input IBU; 
 input IBV; 
 input IBW; 
 input IBX; 
 input IBY; 
 input IBZ; 
 input ICB; 
 input ICC; 
 input ICD; 
 input ICE; 
 input ICF; 
 input ICG; 
 input ICH; 
 input ICI; 
 input ICK; 
 input ICL; 
 input ICM; 
 input ICN; 
 input ICO; 
 input ICP; 
 input ICQ; 
 input ICS; 
 input ICT; 
 input ICU; 
 input ICV; 
 input ICW; 
 input ICX; 
 input ICY; 
 input ICZ; 
 input IDA; 
 input IDB; 
 input IDC; 
 input IDD; 
 input IDE; 
 input IDF; 
 input IDG; 
 input IDH; 
 input IDI; 
 input IDJ; 
 input IDK; 
 input IDL; 
 input IDM; 
 input IDN; 
 input IDO; 
 input IDP; 
 input IDQ; 
 input IDR; 
 input IDS; 
 input IDT; 
 input IDU; 
 input IDV; 
 input IDW; 
 input IDX; 
 input IDY; 
 input IDZ; 
 input IEF; 
 input IEG; 
 input IEH; 
 input IEI; 
 input IEO; 
 input IEP; 
 input IEQ; 
 input IFFF ; 
 input IFO; 
 input IGA; 
 input IGB; 
 input IGC; 
 input IGD; 
 input IGE; 
 input IGF; 
 input IGG; 
 input IGH; 
 input IGI; 
 input IGJ; 
 input IGK; 
 input IGL; 
 input IGM; 
 input IGN; 
 input IGO; 
 input IGP; 
 input IHA; 
 input IHB; 
 input IHC; 
 input IHD; 
 input IHE; 
 input IHF; 
 input IHG; 
 input IHH; 
 input IHI; 
 input IHJ; 
 input IHK; 
 input IHL; 
 input IHM; 
 input IHN; 
 input IHO; 
 input IHP; 
 input IUA; 
 input IUB; 
 input IVA; 
 input IVB; 
 input IVC; 
 input IVD; 
 input IVE; 
 input IVF; 
 output OAA; 
 output OAB; 
 output OAC; 
 output OAD; 
 output OAE; 
 output OAF; 
 output OAG; 
 output OAH; 
 output OAI; 
 output OAJ; 
 output OAK; 
 output OAL; 
 output OAM; 
 output OAN; 
 output OAO; 
 output OAP; 
 output OAQ; 
 output OAR; 
 output OAS; 
 output OAT; 
 output OAU; 
 output OAV; 
 output OAW; 
 output OAX; 
 output OBA; 
 output OBB; 
 output OBC; 
 output OBD; 
 output OBE; 
 output OBF; 
 output OBG; 
 output OBH; 
 output OBI; 
 output OBJ; 
 output OBK; 
 output OBL; 
 output OBM; 
 output OBN; 
 output OBO; 
 output OBP; 
 output OBQ; 
 output OBR; 
 output OBS; 
 output OBT; 
 output OBU; 
 output OBV; 
 output OBW; 
 output OBX; 
 output OCA; 
 output OCB; 
 output OCC; 
 output OCD; 
 output OCE; 
 output OCF; 
 output OCG; 
 output OCH; 
 output OCI; 
 output OCJ; 
 output OCK; 
 output OCL; 
 output OCM; 
 output OCN; 
 output OCO; 
 output OCP; 
 output ODA; 
 output ODB; 
 output ODC; 
 output OEA; 
 output OEB; 
 output OEC; 
 output OFA; 
 output OFB; 
 output OFC; 
 output OGA; 
 output OGB; 
 output OGC; 
 output OHA; 
 output OHB; 
 output OHC; 
 output OIA; 
 output OIB; 
 output OIC; 
 output OID; 
 output OJA; 
 output OJB; 
 output OJC; 
 output OJD; 
 output OJE; 
 output OJF; 
 output OKA; 
 output OLA; 
 output OMA; 
 output OMB; 
 output OMC; 
 output OMD; 
  
  
reg  AAA ;
reg  AAB ;
reg  AAC ;
reg  AAD ;
reg  AAE ;
reg  AAF ;
reg  AAG ;
reg  AAH ;
reg  AAI ;
reg  AAJ ;
reg  AAK ;
reg  AAL ;
reg  AAM ;
reg  AAN ;
reg  AAO ;
reg  AAP ;
reg  ABB ;
reg  ABC ;
reg  ABD ;
reg  ABE ;
reg  ABF ;
reg  ABG ;
reg  ABH ;
reg  ABI ;
reg  ABJ ;
reg  ABK ;
reg  ABL ;
reg  ABM ;
reg  ABN ;
reg  ABO ;
reg  ABP ;
reg  ACA ;
reg  ACB ;
reg  ACC ;
reg  ACD ;
reg  ACE ;
reg  ACF ;
reg  ACG ;
reg  ACH ;
reg  ACI ;
reg  ACJ ;
reg  ACK ;
reg  ACL ;
reg  ACM ;
reg  ACN ;
reg  ACO ;
reg  ACP ;
reg  ADA ;
reg  ADB ;
reg  ADC ;
reg  ADD ;
reg  ADE ;
reg  ADF ;
reg  ADG ;
reg  ADH ;
reg  ADI ;
reg  ADJ ;
reg  ADK ;
reg  ADL ;
reg  ADM ;
reg  ADN ;
reg  ADO ;
reg  ADP ;
reg  AEA ;
reg  AEB ;
reg  AEC ;
reg  AED ;
reg  AEE ;
reg  AEF ;
reg  AEG ;
reg  AEH ;
reg  AEI ;
reg  AEJ ;
reg  AEK ;
reg  AEL ;
reg  AEM ;
reg  AEN ;
reg  AEO ;
reg  AEP ;
reg  AFA ;
reg  AFB ;
reg  AFC ;
reg  AFD ;
reg  AFE ;
reg  AFF ;
reg  AFG ;
reg  AFH ;
reg  AFI ;
reg  AFJ ;
reg  AFK ;
reg  AFL ;
reg  AFM ;
reg  AFN ;
reg  AFO ;
reg  AFP ;
reg  AGA ;
reg  AGB ;
reg  AGC ;
reg  AGD ;
reg  AGE ;
reg  AGF ;
reg  AGG ;
reg  AGH ;
reg  AGI ;
reg  AGJ ;
reg  AGK ;
reg  AGL ;
reg  AGM ;
reg  AGN ;
reg  AGO ;
reg  AGP ;
reg  AHA ;
reg  AHB ;
reg  AHC ;
reg  AHD ;
reg  AHE ;
reg  AHF ;
reg  AHG ;
reg  AHH ;
reg  AHI ;
reg  AHJ ;
reg  AHK ;
reg  AHL ;
reg  AHM ;
reg  AHN ;
reg  AHO ;
reg  AHP ;
reg  AIA ;
reg  AIB ;
reg  AIC ;
reg  AID ;
reg  AIE ;
reg  AIF ;
reg  AIG ;
reg  AIH ;
reg  AII ;
reg  AIJ ;
reg  AIK ;
reg  AIL ;
reg  AIM ;
reg  AIN ;
reg  AIO ;
reg  AIP ;
reg  AJA ;
reg  AJB ;
reg  AJC ;
reg  AJD ;
reg  AJE ;
reg  AJF ;
reg  AJG ;
reg  AJH ;
reg  AJI ;
reg  AJJ ;
reg  AJK ;
reg  AJL ;
reg  AJM ;
reg  AJN ;
reg  AJO ;
reg  AJP ;
reg  AKA ;
reg  AKB ;
reg  AKC ;
reg  AKD ;
reg  AKE ;
reg  AKF ;
reg  AKG ;
reg  AKH ;
reg  AKI ;
reg  AKJ ;
reg  AKK ;
reg  AKL ;
reg  AKM ;
reg  AKN ;
reg  AKO ;
reg  AKP ;
reg  ALA ;
reg  ALB ;
reg  ALC ;
reg  ALD ;
reg  ALE ;
reg  ALF ;
reg  ALG ;
reg  ALH ;
reg  ALI ;
reg  ALJ ;
reg  ALK ;
reg  ALL ;
reg  ALM ;
reg  ALN ;
reg  ALO ;
reg  ALP ;
reg  AMA ;
reg  AMB ;
reg  AMC ;
reg  AMD ;
reg  AME ;
reg  AMF ;
reg  AMG ;
reg  AMH ;
reg  AMI ;
reg  AMJ ;
reg  AMK ;
reg  AML ;
reg  AMM ;
reg  AMN ;
reg  AMO ;
reg  AMP ;
reg  ANA ;
reg  ANB ;
reg  ANC ;
reg  ANDD  ;
reg  ANE ;
reg  ANF ;
reg  ANG ;
reg  ANH ;
reg  ANI ;
reg  ANJ ;
reg  ANK ;
reg  ANL ;
reg  ANM ;
reg  ANN ;
reg  ANO ;
reg  ANP ;
reg  AOA ;
reg  AOB ;
reg  AOC ;
reg  AOD ;
reg  AOE ;
reg  AOF ;
reg  AOG ;
reg  AOH ;
reg  AOI ;
reg  AOJ ;
reg  AOK ;
reg  AOL ;
reg  AOM ;
reg  AON ;
reg  AOO ;
reg  AOP ;
reg  BAA ;
reg  bab ;
reg  bac ;
reg  BAD ;
reg  BAE ;
reg  BAF ;
reg  BAG ;
reg  BAH ;
reg  BAI ;
reg  BAJ ;
reg  BAK ;
reg  BAL ;
reg  BAM ;
reg  BAN ;
reg  BAO ;
reg  BAP ;
reg  BAQ ;
reg  BAR ;
reg  BAS ;
reg  BAT ;
reg  BAU ;
reg  BAV ;
reg  BAW ;
reg  BAX ;
reg  BAY ;
reg  BAZ ;
reg  BBA ;
reg  BBB ;
reg  BBC ;
reg  BBD ;
reg  BBE ;
reg  BBF ;
reg  BBG ;
reg  BBH ;
reg  BBI ;
reg  BBJ ;
reg  BBK ;
reg  BBL ;
reg  BBM ;
reg  BBN ;
reg  BBO ;
reg  BBP ;
reg  BBQ ;
reg  BBR ;
reg  BBS ;
reg  BBT ;
reg  BBU ;
reg  BBV ;
reg  BBW ;
reg  BBX ;
reg  BBY ;
reg  BBZ ;
reg  BCB ;
reg  BCC ;
reg  BCD ;
reg  BCE ;
reg  BCF ;
reg  bcg ;
reg  bch ;
reg  bci ;
reg  bcj ;
reg  BCK ;
reg  BCL ;
reg  BCM ;
reg  BCN ;
reg  BCO ;
reg  bcp ;
reg  bcq ;
reg  bcr ;
reg  BCS ;
reg  BCT ;
reg  BCU ;
reg  BCV ;
reg  BCW ;
reg  BCX ;
reg  BCY ;
reg  BCZ ;
reg  BDA ;
reg  BDB ;
reg  BDC ;
reg  BDD ;
reg  BDE ;
reg  BDF ;
reg  BDG ;
reg  BDH ;
reg  BDI ;
reg  BDJ ;
reg  BDK ;
reg  BDL ;
reg  BDM ;
reg  BDN ;
reg  BDO ;
reg  BDP ;
reg  BDQ ;
reg  BDR ;
reg  BDS ;
reg  BDT ;
reg  BDU ;
reg  BDV ;
reg  BDW ;
reg  BDX ;
reg  BDY ;
reg  BDZ ;
reg  bea ;
reg  beb ;
reg  bec ;
reg  bed ;
reg  bee ;
reg  bef ;
reg  beg ;
reg  beh ;
reg  bei ;
reg  bej ;
reg  bek ;
reg  bel ;
reg  bem ;
reg  ben ;
reg  beo ;
reg  bep ;
reg  BFA ;
reg  BFB ;
reg  BFC ;
reg  BFD ;
reg  BFE ;
reg  BFF ;
reg  BFG ;
reg  BFH ;
reg  BFI ;
reg  BFJ ;
reg  BFK ;
reg  BFL ;
reg  BFM ;
reg  BFN ;
reg  BFO ;
reg  BFP ;
reg  BGA ;
reg  BGB ;
reg  BGC ;
reg  BGD ;
reg  BGE ;
reg  BGF ;
reg  BGG ;
reg  BGH ;
reg  BGI ;
reg  BGJ ;
reg  BGK ;
reg  BGL ;
reg  BGM ;
reg  BGN ;
reg  BGO ;
reg  BGP ;
reg  BHA ;
reg  BHB ;
reg  BHC ;
reg  BHD ;
reg  BHE ;
reg  BHF ;
reg  BHG ;
reg  BHH ;
reg  BHI ;
reg  BHJ ;
reg  BHK ;
reg  BHL ;
reg  BHM ;
reg  BHN ;
reg  BHO ;
reg  BHP ;
reg  FAB ;
reg  FAC ;
reg  FAD ;
reg  FAE ;
reg  FBB ;
reg  FBC ;
reg  FBD ;
reg  FBE ;
reg  fbf ;
reg  fbg ;
reg  fbh ;
reg  FCB ;
reg  FCC ;
reg  FCD ;
reg  FCE ;
reg  fcf ;
reg  fcg ;
reg  fch ;
reg  FDB ;
reg  FDC ;
reg  fdf ;
reg  fdg ;
reg  FEA ;
reg  FEB ;
reg  FEC ;
reg  FED ;
reg  FFA ;
reg  FFB ;
reg  FFC ;
reg  FFD ;
reg  FFE ;
reg  FGA ;
reg  FGB ;
reg  FGC ;
reg  FGD ;
reg  FGE ;
reg  FHA ;
reg  FHB ;
reg  FHC ;
reg  FIA ;
reg  GAA ;
reg  GAB ;
reg  GAC ;
reg  GAD ;
reg  GAE ;
reg  GBB ;
reg  GBC ;
reg  GBD ;
reg  GBE ;
reg  gbf ;
reg  gbg ;
reg  gbh ;
reg  GCB ;
reg  GCC ;
reg  GCD ;
reg  GCE ;
reg  gcf ;
reg  gcg ;
reg  gch ;
reg  GDB ;
reg  GDC ;
reg  GDD ;
reg  GDE ;
reg  gdf ;
reg  gdg ;
reg  gdh ;
reg  GEB ;
reg  GEC ;
reg  GED ;
reg  GEE ;
reg  gef ;
reg  geg ;
reg  geh ;
reg  GFB ;
reg  GFC ;
reg  GFD ;
reg  GFE ;
reg  gff ;
reg  gfg ;
reg  gfh ;
reg  GGB ;
reg  GGC ;
reg  GGD ;
reg  GGE ;
reg  ggf ;
reg  ggg ;
reg  ggh ;
reg  GHB ;
reg  GHC ;
reg  GHD ;
reg  GHE ;
reg  ghf ;
reg  ghg ;
reg  ghh ;
reg  gib ;
reg  GIC ;
reg  GID ;
reg  GIE ;
reg  gif ;
reg  gig ;
reg  gih ;
reg  GJB ;
reg  GJC ;
reg  GJD ;
reg  GJE ;
reg  gjf ;
reg  gjg ;
reg  gjh ;
reg  GKB ;
reg  GKC ;
reg  GKD ;
reg  GKE ;
reg  gkf ;
reg  gkg ;
reg  gkh ;
reg  GLB ;
reg  GLC ;
reg  GLD ;
reg  GLE ;
reg  glf ;
reg  glg ;
reg  glh ;
reg  GMB ;
reg  gmf ;
reg  HAA ;
reg  HAB ;
reg  HAC ;
reg  HAD ;
reg  HBA ;
reg  HBB ;
reg  HBC ;
reg  HBD ;
reg  HBE ;
reg  HCA ;
reg  HCB ;
reg  HCC ;
reg  HCD ;
reg  hce ;
reg  HDA ;
reg  HDB ;
reg  HDC ;
reg  HDD ;
reg  HDE ;
reg  HEA ;
reg  HEB ;
reg  HEC ;
reg  HED ;
reg  hee ;
reg  HFA ;
reg  HFB ;
reg  HFC ;
reg  HFD ;
reg  hfe ;
reg  hff ;
reg  HGA ;
reg  HGB ;
reg  HGC ;
reg  HGD ;
reg  hge ;
reg  hgf ;
reg  HHA ;
reg  HHB ;
reg  HHC ;
reg  HHD ;
reg  hhe ;
reg  hhf ;
reg  HIA ;
reg  HIB ;
reg  HIC ;
reg  HID ;
reg  hie ;
reg  HJA ;
reg  HJB ;
reg  HJC ;
reg  HJD ;
reg  hje ;
reg  hjf ;
reg  HKA ;
reg  HKB ;
reg  HKC ;
reg  HKD ;
reg  hke ;
reg  hkf ;
reg  HLA ;
reg  HLB ;
reg  HLC ;
reg  HLD ;
reg  hle ;
reg  hlf ;
reg  HMA ;
reg  JEA ;
reg  JED ;
reg  LAA ;
reg  LAB ;
reg  LAC ;
reg  LAD ;
reg  LBA ;
reg  LBB ;
reg  LBC ;
reg  LBD ;
reg  LBE ;
reg  LBF ;
reg  LBG ;
reg  LBH ;
reg  LCA ;
reg  LCB ;
reg  LCC ;
reg  LCD ;
reg  LCE ;
reg  LCF ;
reg  LCG ;
reg  LCH ;
reg  LDA ;
reg  LDB ;
reg  LDC ;
reg  LDD ;
reg  LDE ;
reg  LDF ;
reg  LDG ;
reg  LDH ;
reg  LEA ;
reg  LEB ;
reg  LEC ;
reg  LED ;
reg  LEE ;
reg  LEF ;
reg  LEG ;
reg  LEH ;
reg  LFA ;
reg  LFB ;
reg  LFC ;
reg  LFD ;
reg  LFE ;
reg  LFF ;
reg  LFG ;
reg  LFH ;
reg  LGA ;
reg  LGB ;
reg  LGC ;
reg  LGD ;
reg  LGE ;
reg  LGF ;
reg  LGG ;
reg  LGH ;
reg  LHA ;
reg  LHB ;
reg  LHC ;
reg  LHD ;
reg  LHE ;
reg  LHF ;
reg  LHG ;
reg  LHH ;
reg  LIA ;
reg  LIB ;
reg  LIC ;
reg  LID ;
reg  LIE ;
reg  LIF ;
reg  LIG ;
reg  LIH ;
reg  LJA ;
reg  LJB ;
reg  LJC ;
reg  LJD ;
reg  LJE ;
reg  LJF ;
reg  LJG ;
reg  LJH ;
reg  LKA ;
reg  LKB ;
reg  LKC ;
reg  LKD ;
reg  LKE ;
reg  LKF ;
reg  LKG ;
reg  LKH ;
reg  LLA ;
reg  LLB ;
reg  LLC ;
reg  LLD ;
reg  LLE ;
reg  LLF ;
reg  LLG ;
reg  LLH ;
reg  LMA ;
reg  LME ;
reg  OAA ;
reg  OAB ;
reg  OAC ;
reg  OAD ;
reg  OAE ;
reg  OAF ;
reg  OAG ;
reg  OAH ;
reg  OAI ;
reg  OAJ ;
reg  OAK ;
reg  OAL ;
reg  OAM ;
reg  OAN ;
reg  OAO ;
reg  OAP ;
reg  OAQ ;
reg  OAR ;
reg  OAS ;
reg  OAT ;
reg  OAU ;
reg  OAV ;
reg  OAW ;
reg  OAX ;
reg  OBA ;
reg  OBB ;
reg  OBC ;
reg  OBD ;
reg  OBE ;
reg  OBF ;
reg  OBG ;
reg  OBH ;
reg  OBI ;
reg  OBJ ;
reg  OBK ;
reg  OBL ;
reg  OBM ;
reg  OBN ;
reg  OBO ;
reg  OBP ;
reg  OBQ ;
reg  OBR ;
reg  OBS ;
reg  OBT ;
reg  OBU ;
reg  OBV ;
reg  OBW ;
reg  OBX ;
reg  OCA ;
reg  OCB ;
reg  OCC ;
reg  OCD ;
reg  OCE ;
reg  OCF ;
reg  OCG ;
reg  OCH ;
reg  OCI ;
reg  OCJ ;
reg  OCK ;
reg  OCL ;
reg  OCM ;
reg  OCN ;
reg  OCO ;
reg  OCP ;
reg  ODA ;
reg  ODB ;
reg  ODC ;
reg  OEA ;
reg  OEB ;
reg  OEC ;
reg  OFA ;
reg  OFB ;
reg  OFC ;
reg  OGA ;
reg  OGB ;
reg  OGC ;
reg  OHA ;
reg  OHB ;
reg  OHC ;
reg  OIA ;
reg  OIB ;
reg  OIC ;
reg  OID ;
reg  OJA ;
reg  OJB ;
reg  OJC ;
reg  OJD ;
reg  OJE ;
reg  OJF ;
reg  OKA ;
reg  OLA ;
reg  OMA ;
reg  OMB ;
reg  OMC ;
reg  OMD ;
reg  pab ;
reg  pac ;
reg  pad ;
reg  pae ;
reg  paf ;
reg  pag ;
reg  pah ;
reg  pai ;
reg  PAJ ;
reg  PAK ;
reg  PAL ;
reg  PAM ;
reg  PBA ;
reg  pca ;
reg  PDB ;
reg  PDC ;
reg  PDD ;
reg  PDE ;
reg  PDF ;
reg  pdg ;
reg  pdh ;
reg  pdi ;
reg  pdj ;
reg  pdk ;
reg  pdl ;
reg  PDM ;
reg  PDN ;
reg  PDO ;
reg  qaa ;
reg  qab ;
reg  qac ;
reg  qad ;
reg  qae ;
reg  qaf ;
reg  qag ;
reg  qah ;
reg  qai ;
reg  qaj ;
reg  qba ;
reg  qbb ;
reg  qbc ;
reg  qbd ;
reg  qbe ;
reg  qbf ;
reg  qbg ;
reg  qbh ;
reg  qbi ;
reg  qbj ;
reg  qbk ;
reg  qbl ;
reg  qbm ;
reg  qca ;
reg  qcb ;
reg  qcc ;
reg  QCD ;
reg  qce ;
reg  qcf ;
reg  qcg ;
reg  qch ;
reg  qci ;
reg  qcj ;
reg  qck ;
reg  qda ;
reg  qdb ;
reg  qdc ;
reg  qdd ;
reg  qde ;
reg  qdf ;
reg  qdg ;
reg  qdh ;
reg  qdi ;
reg  qdj ;
reg  qdk ;
reg  qdl ;
reg  qdm ;
reg  qdn ;
reg  qdo ;
reg  qea ;
reg  qeb ;
reg  qec ;
reg  qed ;
reg  qee ;
reg  qef ;
reg  qeg ;
reg  qeh ;
reg  qei ;
reg  qej ;
reg  qek ;
reg  qel ;
reg  qem ;
reg  qfa ;
reg  qfb ;
reg  qfc ;
reg  qfd ;
reg  qfe ;
reg  qff ;
reg  qfg ;
reg  qfh ;
reg  qfi ;
reg  qfj ;
reg  qfk ;
reg  qga ;
reg  qgb ;
reg  qgc ;
reg  qgd ;
reg  qge ;
reg  qgf ;
reg  qgg ;
reg  qgh ;
reg  qgi ;
reg  qgj ;
reg  qha ;
reg  qhb ;
reg  qhc ;
reg  qhd ;
reg  qhe ;
reg  qhf ;
reg  qhg ;
reg  QIA ;
reg  QJA ;
reg  QJB ;
reg  QJC ;
reg  QJD ;
reg  QJE ;
reg  QJF ;
reg  QJG ;
reg  QJH ;
reg  QJI ;
reg  QJJ ;
reg  QJK ;
reg  QJL ;
reg  QJM ;
reg  QJN ;
reg  QJO ;
reg  QJP ;
reg  QJQ ;
reg  QJR ;
reg  QJS ;
reg  QKA ;
reg  QKB ;
reg  QKC ;
reg  QKD ;
reg  QKE ;
reg  QKF ;
reg  QKL ;
reg  QKM ;
reg  QKN ;
reg  QKO ;
reg  QKP ;
reg  QKQ ;
reg  QKR ;
reg  qks ;
reg  QKT ;
reg  QKU ;
reg  QKV ;
reg  QKW ;
reg  QKX ;
reg  QKY ;
reg  QLA ;
reg  QLB ;
reg  QLC ;
reg  QLD ;
reg  QLE ;
reg  QLF ;
reg  QLG ;
reg  QLH ;
reg  QLI ;
reg  QLJ ;
reg  QLK ;
reg  QLL ;
reg  QLM ;
reg  QLN ;
reg  QLO ;
reg  QLP ;
reg  QLQ ;
reg  QLR ;
reg  QLS ;
reg  QLT ;
reg  QLU ;
reg  QLV ;
reg  qma ;
reg  QMB ;
reg  QMC ;
reg  QMD ;
reg  qme ;
reg  QMF ;
reg  QMG ;
reg  QMH ;
reg  QMI ;
reg  QMJ ;
reg  qmk ;
reg  qml ;
reg  qmm ;
reg  qmn ;
reg  qmo ;
reg  QNA ;
reg  QNE ;
reg  QNF ;
reg  QNH ;
reg  QNI ;
reg  QNJ ;
reg  QNK ;
reg  qnl ;
reg  qnm ;
reg  QNO ;
reg  QOA ;
reg  QOB ;
reg  qoc ;
reg  QOD ;
reg  QOE ;
reg  QOF ;
reg  QOG ;
reg  QOH ;
reg  QOI ;
reg  QOJ ;
reg  QOL ;
reg  QPA ;
reg  QPB ;
reg  QPC ;
reg  QPD ;
reg  QQA ;
reg  QQB ;
reg  QRA ;
reg  QRB ;
reg  QRC ;
reg  QRD ;
reg  QRE ;
reg  QRF ;
reg  QRG ;
reg  QRH ;
reg  QRI ;
reg  QRJ ;
reg  QRK ;
reg  TAA ;
reg  TAB ;
reg  TBA ;
reg  TBB ;
reg  TCA ;
reg  TCB ;
reg  TDA ;
reg  TDB ;
reg  TEA ;
reg  TEB ;
reg  TFA ;
reg  TFB ;
reg  TGA ;
reg  TGB ;
reg  THA ;
reg  THB ;
reg  TIA ;
reg  TIB ;
reg  TKA ;
reg  TKB ;
reg  TKC ;
reg  TKD ;
reg  TKE ;
reg  TKF ;
reg  TKG ;
reg  TKH ;
reg  tki ;
reg  tkj ;
reg  tkk ;
reg  tkl ;
reg  tkm ;
reg  tkn ;
reg  tko ;
reg  tkp ;
reg  TKQ ;
reg  TKR ;
reg  TKS ;
reg  TKT ;
reg  tku ;
reg  tkv ;
reg  tkw ;
reg  tkx ;
reg  TLA ;
reg  TLB ;
reg  TLC ;
reg  TLD ;
reg  TLE ;
reg  TLF ;
reg  TLG ;
reg  TLH ;
reg  TLI ;
reg  TLJ ;
reg  TLK ;
reg  TLL ;
reg  TLM ;
reg  TLN ;
reg  TLO ;
reg  TLP ;
reg  tna ;
reg  tnb ;
reg  tnc ;
reg  tnd ;
reg  tne ;
reg  tnf ;
wire  aaa ;
wire  aab ;
wire  aac ;
wire  aad ;
wire  aae ;
wire  aaf ;
wire  aag ;
wire  aah ;
wire  aai ;
wire  aaj ;
wire  aak ;
wire  aal ;
wire  aam ;
wire  aan ;
wire  aao ;
wire  aap ;
wire  abb ;
wire  abc ;
wire  abd ;
wire  abe ;
wire  abf ;
wire  abg ;
wire  abh ;
wire  abi ;
wire  abj ;
wire  abk ;
wire  abl ;
wire  abm ;
wire  abn ;
wire  abo ;
wire  abp ;
wire  aca ;
wire  acb ;
wire  acc ;
wire  acd ;
wire  ace ;
wire  acf ;
wire  acg ;
wire  ach ;
wire  aci ;
wire  acj ;
wire  ack ;
wire  acl ;
wire  acm ;
wire  acn ;
wire  aco ;
wire  acp ;
wire  ada ;
wire  adb ;
wire  adc ;
wire  add ;
wire  ade ;
wire  adf ;
wire  adg ;
wire  adh ;
wire  adi ;
wire  adj ;
wire  adk ;
wire  adl ;
wire  adm ;
wire  adn ;
wire  ado ;
wire  adp ;
wire  aea ;
wire  aeb ;
wire  aec ;
wire  aed ;
wire  aee ;
wire  aef ;
wire  aeg ;
wire  aeh ;
wire  aei ;
wire  aej ;
wire  aek ;
wire  ael ;
wire  aem ;
wire  aen ;
wire  aeo ;
wire  aep ;
wire  afa ;
wire  afb ;
wire  afc ;
wire  afd ;
wire  afe ;
wire  aff ;
wire  afg ;
wire  afh ;
wire  afi ;
wire  afj ;
wire  afk ;
wire  afl ;
wire  afm ;
wire  afn ;
wire  afo ;
wire  afp ;
wire  aga ;
wire  agb ;
wire  agc ;
wire  agd ;
wire  age ;
wire  agf ;
wire  agg ;
wire  agh ;
wire  agi ;
wire  agj ;
wire  agk ;
wire  agl ;
wire  agm ;
wire  agn ;
wire  ago ;
wire  agp ;
wire  aha ;
wire  ahb ;
wire  ahc ;
wire  ahd ;
wire  ahe ;
wire  ahf ;
wire  ahg ;
wire  ahh ;
wire  ahi ;
wire  ahj ;
wire  ahk ;
wire  ahl ;
wire  ahm ;
wire  ahn ;
wire  aho ;
wire  ahp ;
wire  aia ;
wire  aib ;
wire  aic ;
wire  aid ;
wire  aie ;
wire  aif ;
wire  aig ;
wire  aih ;
wire  aii ;
wire  aij ;
wire  aik ;
wire  ail ;
wire  aim ;
wire  ain ;
wire  aio ;
wire  aip ;
wire  aja ;
wire  ajb ;
wire  ajc ;
wire  ajd ;
wire  aje ;
wire  ajf ;
wire  ajg ;
wire  ajh ;
wire  aji ;
wire  ajj ;
wire  ajk ;
wire  ajl ;
wire  ajm ;
wire  ajn ;
wire  ajo ;
wire  ajp ;
wire  aka ;
wire  akb ;
wire  akc ;
wire  akd ;
wire  ake ;
wire  akf ;
wire  akg ;
wire  akh ;
wire  aki ;
wire  akj ;
wire  akk ;
wire  akl ;
wire  akm ;
wire  akn ;
wire  ako ;
wire  akp ;
wire  ala ;
wire  alb ;
wire  alc ;
wire  ald ;
wire  ale ;
wire  alf ;
wire  alg ;
wire  alh ;
wire  ali ;
wire  alj ;
wire  alk ;
wire  all ;
wire  alm ;
wire  aln ;
wire  alo ;
wire  alp ;
wire  ama ;
wire  amb ;
wire  amc ;
wire  amd ;
wire  ame ;
wire  amf ;
wire  amg ;
wire  amh ;
wire  ami ;
wire  amj ;
wire  amk ;
wire  aml ;
wire  amm ;
wire  amn ;
wire  amo ;
wire  amp ;
wire  ana ;
wire  anb ;
wire  anc ;
wire  andd  ;
wire  ane ;
wire  anf ;
wire  ang ;
wire  anh ;
wire  ani ;
wire  anj ;
wire  ank ;
wire  anl ;
wire  anm ;
wire  ann ;
wire  ano ;
wire  anp ;
wire  aoa ;
wire  aob ;
wire  aoc ;
wire  aod ;
wire  aoe ;
wire  aof ;
wire  aog ;
wire  aoh ;
wire  aoi ;
wire  aoj ;
wire  aok ;
wire  aol ;
wire  aom ;
wire  aon ;
wire  aoo ;
wire  aop ;
wire  baa ;
wire  BAB ;
wire  BAC ;
wire  bad ;
wire  bae ;
wire  baf ;
wire  bag ;
wire  bah ;
wire  bai ;
wire  baj ;
wire  bak ;
wire  bal ;
wire  bam ;
wire  ban ;
wire  bao ;
wire  bap ;
wire  baq ;
wire  bar ;
wire  bas ;
wire  bat ;
wire  bau ;
wire  bav ;
wire  baw ;
wire  bax ;
wire  bay ;
wire  baz ;
wire  bba ;
wire  bbb ;
wire  bbc ;
wire  bbd ;
wire  bbe ;
wire  bbf ;
wire  bbg ;
wire  bbh ;
wire  bbi ;
wire  bbj ;
wire  bbk ;
wire  bbl ;
wire  bbm ;
wire  bbn ;
wire  bbo ;
wire  bbp ;
wire  bbq ;
wire  bbr ;
wire  bbs ;
wire  bbt ;
wire  bbu ;
wire  bbv ;
wire  bbw ;
wire  bbx ;
wire  bby ;
wire  bbz ;
wire  bcb ;
wire  bcc ;
wire  bcd ;
wire  bce ;
wire  bcf ;
wire  BCG ;
wire  BCH ;
wire  BCI ;
wire  BCJ ;
wire  bck ;
wire  bcl ;
wire  bcm ;
wire  bcn ;
wire  bco ;
wire  BCP ;
wire  BCQ ;
wire  BCR ;
wire  bcs ;
wire  bct ;
wire  bcu ;
wire  bcv ;
wire  bcw ;
wire  bcx ;
wire  bcy ;
wire  bcz ;
wire  bda ;
wire  bdb ;
wire  bdc ;
wire  bdd ;
wire  bde ;
wire  bdf ;
wire  bdg ;
wire  bdh ;
wire  bdi ;
wire  bdj ;
wire  bdk ;
wire  bdl ;
wire  bdm ;
wire  bdn ;
wire  bdo ;
wire  bdp ;
wire  bdq ;
wire  bdr ;
wire  bds ;
wire  bdt ;
wire  bdu ;
wire  bdv ;
wire  bdw ;
wire  bdx ;
wire  bdy ;
wire  bdz ;
wire  BEA ;
wire  BEB ;
wire  BEC ;
wire  BED ;
wire  BEE ;
wire  BEF ;
wire  BEG ;
wire  BEH ;
wire  BEI ;
wire  BEJ ;
wire  BEK ;
wire  BEL ;
wire  BEM ;
wire  BEN ;
wire  BEO ;
wire  BEP ;
wire  bfa ;
wire  bfb ;
wire  bfc ;
wire  bfd ;
wire  bfe ;
wire  bff ;
wire  bfg ;
wire  bfh ;
wire  bfi ;
wire  bfj ;
wire  bfk ;
wire  bfl ;
wire  bfm ;
wire  bfn ;
wire  bfo ;
wire  bfp ;
wire  bga ;
wire  bgb ;
wire  bgc ;
wire  bgd ;
wire  bge ;
wire  bgf ;
wire  bgg ;
wire  bgh ;
wire  bgi ;
wire  bgj ;
wire  bgk ;
wire  bgl ;
wire  bgm ;
wire  bgn ;
wire  bgo ;
wire  bgp ;
wire  bha ;
wire  bhb ;
wire  bhc ;
wire  bhd ;
wire  bhe ;
wire  bhf ;
wire  bhg ;
wire  bhh ;
wire  bhi ;
wire  bhj ;
wire  bhk ;
wire  bhl ;
wire  bhm ;
wire  bhn ;
wire  bho ;
wire  bhp ;
wire  caa ;
wire  CAA ;
wire  cab ;
wire  CAB ;
wire  cac ;
wire  CAC ;
wire  cad ;
wire  CAD ;
wire  cba ;
wire  CBA ;
wire  cbb ;
wire  CBB ;
wire  cbc ;
wire  CBC ;
wire  cbd ;
wire  CBD ;
wire  cca ;
wire  CCA ;
wire  ccb ;
wire  CCB ;
wire  ccc ;
wire  CCC ;
wire  ccd ;
wire  CCD ;
wire  cda ;
wire  CDA ;
wire  cdb ;
wire  CDB ;
wire  cdc ;
wire  CDC ;
wire  cdd ;
wire  CDD ;
wire  cea ;
wire  CEA ;
wire  ceb ;
wire  CEB ;
wire  cec ;
wire  CEC ;
wire  ced ;
wire  CED ;
wire  cfa ;
wire  CFA ;
wire  cfb ;
wire  CFB ;
wire  cfc ;
wire  CFC ;
wire  cfd ;
wire  CFD ;
wire  cga ;
wire  CGA ;
wire  cgb ;
wire  CGB ;
wire  cgc ;
wire  CGC ;
wire  cgd ;
wire  CGD ;
wire  cha ;
wire  CHA ;
wire  chb ;
wire  CHB ;
wire  chc ;
wire  CHC ;
wire  chd ;
wire  CHD ;
wire  cia ;
wire  CIA ;
wire  cib ;
wire  CIB ;
wire  cic ;
wire  CIC ;
wire  cid ;
wire  CID ;
wire  cja ;
wire  CJA ;
wire  cjb ;
wire  CJB ;
wire  cjc ;
wire  CJC ;
wire  cjd ;
wire  CJD ;
wire  cka ;
wire  CKA ;
wire  ckb ;
wire  CKB ;
wire  ckc ;
wire  CKC ;
wire  ckd ;
wire  CKD ;
wire  cla ;
wire  CLA ;
wire  clb ;
wire  CLB ;
wire  clc ;
wire  CLC ;
wire  cld ;
wire  CLD ;
wire  cma ;
wire  CMA ;
wire  cna ;
wire  CNA ;
wire  daa ;
wire  DAA ;
wire  dab ;
wire  DAB ;
wire  dac ;
wire  DAC ;
wire  dad ;
wire  DAD ;
wire  dba ;
wire  DBA ;
wire  dbb ;
wire  DBB ;
wire  dbc ;
wire  DBC ;
wire  dbd ;
wire  DBD ;
wire  dca ;
wire  DCA ;
wire  dcb ;
wire  DCB ;
wire  dcc ;
wire  DCC ;
wire  dcd ;
wire  DCD ;
wire  dda ;
wire  DDA ;
wire  ddb ;
wire  DDB ;
wire  ddc ;
wire  DDC ;
wire  ddd ;
wire  DDD ;
wire  dea ;
wire  DEA ;
wire  deb ;
wire  DEB ;
wire  dec ;
wire  DEC ;
wire  ded ;
wire  DED ;
wire  dfa ;
wire  DFA ;
wire  dfb ;
wire  DFB ;
wire  dfc ;
wire  DFC ;
wire  dfd ;
wire  DFD ;
wire  dga ;
wire  DGA ;
wire  dgb ;
wire  DGB ;
wire  dgc ;
wire  DGC ;
wire  dgd ;
wire  DGD ;
wire  dha ;
wire  DHA ;
wire  dhb ;
wire  DHB ;
wire  dhc ;
wire  DHC ;
wire  dhd ;
wire  DHD ;
wire  dia ;
wire  DIA ;
wire  dib ;
wire  DIB ;
wire  dic ;
wire  DIC ;
wire  did ;
wire  DID ;
wire  dja ;
wire  DJA ;
wire  djb ;
wire  DJB ;
wire  djc ;
wire  DJC ;
wire  djd ;
wire  DJD ;
wire  dka ;
wire  DKA ;
wire  dkb ;
wire  DKB ;
wire  dkc ;
wire  DKC ;
wire  dkd ;
wire  DKD ;
wire  dla ;
wire  DLA ;
wire  dlb ;
wire  DLB ;
wire  dlc ;
wire  DLC ;
wire  dld ;
wire  DLD ;
wire  dma ;
wire  DMA ;
wire  eaa ;
wire  EAA ;
wire  eab ;
wire  EAB ;
wire  eac ;
wire  EAC ;
wire  ead ;
wire  EAD ;
wire  eae ;
wire  EAE ;
wire  eaf ;
wire  EAF ;
wire  eag ;
wire  EAG ;
wire  eah ;
wire  EAH ;
wire  eai ;
wire  EAI ;
wire  eaj ;
wire  EAJ ;
wire  eak ;
wire  EAK ;
wire  eal ;
wire  EAL ;
wire  eam ;
wire  EAM ;
wire  ean ;
wire  EAN ;
wire  eao ;
wire  EAO ;
wire  eba ;
wire  EBA ;
wire  ebb ;
wire  EBB ;
wire  ebc ;
wire  EBC ;
wire  ebd ;
wire  EBD ;
wire  ebe ;
wire  EBE ;
wire  ebf ;
wire  EBF ;
wire  ebg ;
wire  EBG ;
wire  ebh ;
wire  EBH ;
wire  ebi ;
wire  EBI ;
wire  ebj ;
wire  EBJ ;
wire  ebk ;
wire  EBK ;
wire  ebl ;
wire  EBL ;
wire  ebm ;
wire  EBM ;
wire  ebn ;
wire  EBN ;
wire  ebo ;
wire  EBO ;
wire  ecb ;
wire  ECB ;
wire  ecc ;
wire  ECC ;
wire  ecd ;
wire  ECD ;
wire  edb ;
wire  EDB ;
wire  edc ;
wire  EDC ;
wire  edd ;
wire  EDD ;
wire  ede ;
wire  EDE ;
wire  edf ;
wire  EDF ;
wire  edg ;
wire  EDG ;
wire  eeb ;
wire  EEB ;
wire  eec ;
wire  EEC ;
wire  eed ;
wire  EED ;
wire  eee ;
wire  EEE ;
wire  eef ;
wire  EEF ;
wire  eeg ;
wire  EEG ;
wire  efb ;
wire  EFB ;
wire  efc ;
wire  EFC ;
wire  efe ;
wire  EFE ;
wire  eff ;
wire  EFF ;
wire  egb ;
wire  EGB ;
wire  egc ;
wire  EGC ;
wire  egd ;
wire  EGD ;
wire  fab ;
wire  fac ;
wire  fad ;
wire  fae ;
wire  fbb ;
wire  fbc ;
wire  fbd ;
wire  fbe ;
wire  FBF ;
wire  FBG ;
wire  FBH ;
wire  fcb ;
wire  fcc ;
wire  fcd ;
wire  fce ;
wire  FCF ;
wire  FCG ;
wire  FCH ;
wire  fdb ;
wire  fdc ;
wire  FDF ;
wire  FDG ;
wire  fea ;
wire  feb ;
wire  fec ;
wire  fed ;
wire  ffa ;
wire  ffb ;
wire  ffc ;
wire  ffd ;
wire  ffe ;
wire  fga ;
wire  fgb ;
wire  fgc ;
wire  fgd ;
wire  fge ;
wire  fha ;
wire  fhb ;
wire  fhc ;
wire  fia ;
wire  gaa ;
wire  gab ;
wire  gac ;
wire  gad ;
wire  gae ;
wire  gbb ;
wire  gbc ;
wire  gbd ;
wire  gbe ;
wire  GBF ;
wire  GBG ;
wire  GBH ;
wire  gcb ;
wire  gcc ;
wire  gcd ;
wire  gce ;
wire  GCF ;
wire  GCG ;
wire  GCH ;
wire  gdb ;
wire  gdc ;
wire  gdd ;
wire  gde ;
wire  GDF ;
wire  GDG ;
wire  GDH ;
wire  geb ;
wire  gec ;
wire  ged ;
wire  gee ;
wire  GEF ;
wire  GEG ;
wire  GEH ;
wire  gfb ;
wire  gfc ;
wire  gfd ;
wire  gfe ;
wire  GFF ;
wire  GFG ;
wire  GFH ;
wire  ggb ;
wire  ggc ;
wire  ggd ;
wire  gge ;
wire  GGF ;
wire  GGG ;
wire  GGH ;
wire  ghb ;
wire  ghc ;
wire  ghd ;
wire  ghe ;
wire  GHF ;
wire  GHG ;
wire  GHH ;
wire  GIB ;
wire  gic ;
wire  gid ;
wire  gie ;
wire  GIF ;
wire  GIG ;
wire  GIH ;
wire  gjb ;
wire  gjc ;
wire  gjd ;
wire  gje ;
wire  GJF ;
wire  GJG ;
wire  GJH ;
wire  gkb ;
wire  gkc ;
wire  gkd ;
wire  gke ;
wire  GKF ;
wire  GKG ;
wire  GKH ;
wire  glb ;
wire  glc ;
wire  gld ;
wire  gle ;
wire  GLF ;
wire  GLG ;
wire  GLH ;
wire  gmb ;
wire  GMF ;
wire  haa ;
wire  hab ;
wire  hac ;
wire  had ;
wire  hba ;
wire  hbb ;
wire  hbc ;
wire  hbd ;
wire  hbe ;
wire  hca ;
wire  hcb ;
wire  hcc ;
wire  hcd ;
wire  HCE ;
wire  hda ;
wire  hdb ;
wire  hdc ;
wire  hdd ;
wire  hde ;
wire  hea ;
wire  heb ;
wire  hec ;
wire  hed ;
wire  HEE ;
wire  hfa ;
wire  hfb ;
wire  hfc ;
wire  hfd ;
wire  HFE ;
wire  HFF ;
wire  hga ;
wire  hgb ;
wire  hgc ;
wire  hgd ;
wire  HGE ;
wire  HGF ;
wire  hha ;
wire  hhb ;
wire  hhc ;
wire  hhd ;
wire  HHE ;
wire  HHF ;
wire  hia ;
wire  hib ;
wire  hic ;
wire  hid ;
wire  HIE ;
wire  hja ;
wire  hjb ;
wire  hjc ;
wire  hjd ;
wire  HJE ;
wire  HJF ;
wire  hka ;
wire  hkb ;
wire  hkc ;
wire  hkd ;
wire  HKE ;
wire  HKF ;
wire  hla ;
wire  hlb ;
wire  hlc ;
wire  hld ;
wire  HLE ;
wire  HLF ;
wire  hma ;
wire  iab ;
wire  iac ;
wire  iad ;
wire  iae ;
wire  iaf ;
wire  iag ;
wire  iah ;
wire  iai ;
wire  iaj ;
wire  iak ;
wire  ial ;
wire  iam ;
wire  ian ;
wire  iao ;
wire  iap ;
wire  iaq ;
wire  iar ;
wire  ias ;
wire  iat ;
wire  iau ;
wire  iav ;
wire  iaw ;
wire  iax ;
wire  iay ;
wire  iaz ;
wire  iba ;
wire  ibb ;
wire  ibc ;
wire  ibd ;
wire  ibe ;
wire  ibf ;
wire  ibg ;
wire  ibh ;
wire  ibi ;
wire  ibj ;
wire  ibk ;
wire  ibl ;
wire  ibm ;
wire  ibn ;
wire  ibo ;
wire  ibp ;
wire  ibq ;
wire  ibr ;
wire  ibs ;
wire  ibt ;
wire  ibu ;
wire  ibv ;
wire  ibw ;
wire  ibx ;
wire  iby ;
wire  ibz ;
wire  icb ;
wire  icc ;
wire  icd ;
wire  ice ;
wire  icf ;
wire  icg ;
wire  ich ;
wire  ici ;
wire  ick ;
wire  icl ;
wire  icm ;
wire  icn ;
wire  ico ;
wire  icp ;
wire  icq ;
wire  ics ;
wire  ict ;
wire  icu ;
wire  icv ;
wire  icw ;
wire  icx ;
wire  icy ;
wire  icz ;
wire  ida ;
wire  idb ;
wire  idc ;
wire  idd ;
wire  ide ;
wire  idf ;
wire  idg ;
wire  idh ;
wire  idi ;
wire  idj ;
wire  idk ;
wire  idl ;
wire  idm ;
wire  idn ;
wire  ido ;
wire  idp ;
wire  idq ;
wire  idr ;
wire  ids ;
wire  idt ;
wire  idu ;
wire  idv ;
wire  idw ;
wire  idx ;
wire  idy ;
wire  idz ;
wire  ief ;
wire  ieg ;
wire  ieh ;
wire  iei ;
wire  ieo ;
wire  iep ;
wire  ieq ;
wire  ifff  ;
wire  ifo ;
wire  iga ;
wire  igb ;
wire  igc ;
wire  igd ;
wire  ige ;
wire  igf ;
wire  igg ;
wire  igh ;
wire  igi ;
wire  igj ;
wire  igk ;
wire  igl ;
wire  igm ;
wire  ign ;
wire  igo ;
wire  igp ;
wire  iha ;
wire  ihb ;
wire  ihc ;
wire  ihd ;
wire  ihe ;
wire  ihf ;
wire  ihg ;
wire  ihh ;
wire  ihi ;
wire  ihj ;
wire  ihk ;
wire  ihl ;
wire  ihm ;
wire  ihn ;
wire  iho ;
wire  ihp ;
wire  iua ;
wire  iub ;
wire  iva ;
wire  ivb ;
wire  ivc ;
wire  ivd ;
wire  ive ;
wire  ivf ;
wire  jaa ;
wire  JAA ;
wire  jab ;
wire  JAB ;
wire  jba ;
wire  JBA ;
wire  jbb ;
wire  JBB ;
wire  jbc ;
wire  JBC ;
wire  jca ;
wire  JCA ;
wire  jcb ;
wire  JCB ;
wire  jcc ;
wire  JCC ;
wire  jcd ;
wire  JCD ;
wire  jdc ;
wire  JDC ;
wire  jdd ;
wire  JDD ;
wire  jde ;
wire  JDE ;
wire  jdf ;
wire  JDF ;
wire  jdg ;
wire  JDG ;
wire  jdi ;
wire  JDI ;
wire  jdj ;
wire  JDJ ;
wire  jdk ;
wire  JDK ;
wire  jdl ;
wire  JDL ;
wire  jdm ;
wire  JDM ;
wire  jdo ;
wire  JDO ;
wire  jea ;
wire  jeb ;
wire  JEB ;
wire  jec ;
wire  JEC ;
wire  jed ;
wire  jee ;
wire  JEE ;
wire  jfa ;
wire  JFA ;
wire  jga ;
wire  JGA ;
wire  jgb ;
wire  JGB ;
wire  jgd ;
wire  JGD ;
wire  jge ;
wire  JGE ;
wire  kaa ;
wire  KAA ;
wire  kab ;
wire  KAB ;
wire  kac ;
wire  KAC ;
wire  kad ;
wire  KAD ;
wire  kbb ;
wire  KBB ;
wire  kbc ;
wire  KBC ;
wire  kbd ;
wire  KBD ;
wire  kbf ;
wire  KBF ;
wire  kbg ;
wire  KBG ;
wire  kbh ;
wire  KBH ;
wire  kcb ;
wire  KCB ;
wire  kcc ;
wire  KCC ;
wire  kcd ;
wire  KCD ;
wire  kcf ;
wire  KCF ;
wire  kcg ;
wire  KCG ;
wire  kch ;
wire  KCH ;
wire  kdb ;
wire  KDB ;
wire  kdc ;
wire  KDC ;
wire  kdd ;
wire  KDD ;
wire  kdf ;
wire  KDF ;
wire  kdg ;
wire  KDG ;
wire  kdh ;
wire  KDH ;
wire  keb ;
wire  KEB ;
wire  kec ;
wire  KEC ;
wire  ked ;
wire  KED ;
wire  kef ;
wire  KEF ;
wire  keg ;
wire  KEG ;
wire  keh ;
wire  KEH ;
wire  kfb ;
wire  KFB ;
wire  kfc ;
wire  KFC ;
wire  kfd ;
wire  KFD ;
wire  kff ;
wire  KFF ;
wire  kfg ;
wire  KFG ;
wire  kfh ;
wire  KFH ;
wire  kgb ;
wire  KGB ;
wire  kgc ;
wire  KGC ;
wire  kgd ;
wire  KGD ;
wire  kgf ;
wire  KGF ;
wire  kgg ;
wire  KGG ;
wire  kgh ;
wire  KGH ;
wire  khb ;
wire  KHB ;
wire  khc ;
wire  KHC ;
wire  khd ;
wire  KHD ;
wire  khf ;
wire  KHF ;
wire  khg ;
wire  KHG ;
wire  khh ;
wire  KHH ;
wire  kib ;
wire  KIB ;
wire  kic ;
wire  KIC ;
wire  kid ;
wire  KID ;
wire  kif ;
wire  KIF ;
wire  kig ;
wire  KIG ;
wire  kih ;
wire  KIH ;
wire  kjb ;
wire  KJB ;
wire  kjc ;
wire  KJC ;
wire  kjd ;
wire  KJD ;
wire  kjf ;
wire  KJF ;
wire  kjg ;
wire  KJG ;
wire  kjh ;
wire  KJH ;
wire  kkb ;
wire  KKB ;
wire  kkc ;
wire  KKC ;
wire  kkd ;
wire  KKD ;
wire  kkf ;
wire  KKF ;
wire  kkg ;
wire  KKG ;
wire  kkh ;
wire  KKH ;
wire  klb ;
wire  KLB ;
wire  klc ;
wire  KLC ;
wire  kld ;
wire  KLD ;
wire  klf ;
wire  KLF ;
wire  klg ;
wire  KLG ;
wire  klh ;
wire  KLH ;
wire  kma ;
wire  KMA ;
wire  kmb ;
wire  KMB ;
wire  kna ;
wire  KNA ;
wire  knb ;
wire  KNB ;
wire  koa ;
wire  KOA ;
wire  kob ;
wire  KOB ;
wire  kpa ;
wire  KPA ;
wire  kpb ;
wire  KPB ;
wire  kqa ;
wire  KQA ;
wire  kqb ;
wire  KQB ;
wire  laa ;
wire  lab ;
wire  lac ;
wire  lad ;
wire  lba ;
wire  lbb ;
wire  lbc ;
wire  lbd ;
wire  lbe ;
wire  lbf ;
wire  lbg ;
wire  lbh ;
wire  lca ;
wire  lcb ;
wire  lcc ;
wire  lcd ;
wire  lce ;
wire  lcf ;
wire  lcg ;
wire  lch ;
wire  lda ;
wire  ldb ;
wire  ldc ;
wire  ldd ;
wire  lde ;
wire  ldf ;
wire  ldg ;
wire  ldh ;
wire  lea ;
wire  leb ;
wire  lec ;
wire  led ;
wire  lee ;
wire  lef ;
wire  leg ;
wire  leh ;
wire  lfa ;
wire  lfb ;
wire  lfc ;
wire  lfd ;
wire  lfe ;
wire  lff ;
wire  lfg ;
wire  lfh ;
wire  lga ;
wire  lgb ;
wire  lgc ;
wire  lgd ;
wire  lge ;
wire  lgf ;
wire  lgg ;
wire  lgh ;
wire  lha ;
wire  lhb ;
wire  lhc ;
wire  lhd ;
wire  lhe ;
wire  lhf ;
wire  lhg ;
wire  lhh ;
wire  lia ;
wire  lib ;
wire  lic ;
wire  lid ;
wire  lie ;
wire  lif ;
wire  lig ;
wire  lih ;
wire  lja ;
wire  ljb ;
wire  ljc ;
wire  ljd ;
wire  lje ;
wire  ljf ;
wire  ljg ;
wire  ljh ;
wire  lka ;
wire  lkb ;
wire  lkc ;
wire  lkd ;
wire  lke ;
wire  lkf ;
wire  lkg ;
wire  lkh ;
wire  lla ;
wire  llb ;
wire  llc ;
wire  lld ;
wire  lle ;
wire  llf ;
wire  llg ;
wire  llh ;
wire  lma ;
wire  lme ;
wire  mae ;
wire  MAE ;
wire  maf ;
wire  MAF ;
wire  mag ;
wire  MAG ;
wire  mah ;
wire  MAH ;
wire  mai ;
wire  MAI ;
wire  maj ;
wire  MAJ ;
wire  mak ;
wire  MAK ;
wire  mal ;
wire  MAL ;
wire  mam ;
wire  MAM ;
wire  man ;
wire  MAN ;
wire  mao ;
wire  MAO ;
wire  map ;
wire  MAP ;
wire  maq ;
wire  MAQ ;
wire  mar ;
wire  MAR ;
wire  mas ;
wire  MAS ;
wire  mat ;
wire  MAT ;
wire  mau ;
wire  MAU ;
wire  mav ;
wire  MAV ;
wire  maw ;
wire  MAW ;
wire  max ;
wire  MAX ;
wire  mba ;
wire  MBA ;
wire  mbb ;
wire  MBB ;
wire  mbc ;
wire  MBC ;
wire  mbd ;
wire  MBD ;
wire  mbe ;
wire  MBE ;
wire  mbf ;
wire  MBF ;
wire  mbg ;
wire  MBG ;
wire  mbh ;
wire  MBH ;
wire  mbi ;
wire  MBI ;
wire  mbj ;
wire  MBJ ;
wire  mbk ;
wire  MBK ;
wire  mbl ;
wire  MBL ;
wire  mbm ;
wire  MBM ;
wire  mbn ;
wire  MBN ;
wire  mbo ;
wire  MBO ;
wire  mbp ;
wire  MBP ;
wire  mbq ;
wire  MBQ ;
wire  mbr ;
wire  MBR ;
wire  mbs ;
wire  MBS ;
wire  mbt ;
wire  MBT ;
wire  mbu ;
wire  MBU ;
wire  mbv ;
wire  MBV ;
wire  mbw ;
wire  MBW ;
wire  mbx ;
wire  MBX ;
wire  mby ;
wire  MBY ;
wire  nbb ;
wire  NBB ;
wire  nbc ;
wire  NBC ;
wire  ncb ;
wire  NCB ;
wire  ncc ;
wire  NCC ;
wire  ndb ;
wire  NDB ;
wire  ndc ;
wire  NDC ;
wire  neb ;
wire  NEB ;
wire  nec ;
wire  NEC ;
wire  oaa ;
wire  oab ;
wire  oac ;
wire  oad ;
wire  oae ;
wire  oaf ;
wire  oag ;
wire  oah ;
wire  oai ;
wire  oaj ;
wire  oak ;
wire  oal ;
wire  oam ;
wire  oan ;
wire  oao ;
wire  oap ;
wire  oaq ;
wire  oar ;
wire  oas ;
wire  oat ;
wire  oau ;
wire  oav ;
wire  oaw ;
wire  oax ;
wire  oba ;
wire  obb ;
wire  obc ;
wire  obd ;
wire  obe ;
wire  obf ;
wire  obg ;
wire  obh ;
wire  obi ;
wire  obj ;
wire  obk ;
wire  obl ;
wire  obm ;
wire  obn ;
wire  obo ;
wire  obp ;
wire  obq ;
wire  obr ;
wire  obs ;
wire  obt ;
wire  obu ;
wire  obv ;
wire  obw ;
wire  obx ;
wire  oca ;
wire  ocb ;
wire  occ ;
wire  ocd ;
wire  oce ;
wire  ocf ;
wire  ocg ;
wire  och ;
wire  oci ;
wire  ocj ;
wire  ock ;
wire  ocl ;
wire  ocm ;
wire  ocn ;
wire  oco ;
wire  ocp ;
wire  oda ;
wire  odb ;
wire  odc ;
wire  oea ;
wire  oeb ;
wire  oec ;
wire  ofa ;
wire  ofb ;
wire  ofc ;
wire  oga ;
wire  ogb ;
wire  ogc ;
wire  oha ;
wire  ohb ;
wire  ohc ;
wire  oia ;
wire  oib ;
wire  oic ;
wire  oid ;
wire  oja ;
wire  ojb ;
wire  ojc ;
wire  ojd ;
wire  oje ;
wire  ojf ;
wire  oka ;
wire  ola ;
wire  oma ;
wire  omb ;
wire  omc ;
wire  omd ;
wire  PAB ;
wire  PAC ;
wire  PAD ;
wire  PAE ;
wire  PAF ;
wire  PAG ;
wire  PAH ;
wire  PAI ;
wire  paj ;
wire  pak ;
wire  pal ;
wire  pam ;
wire  pba ;
wire  PCA ;
wire  pdb ;
wire  pdc ;
wire  pdd ;
wire  pde ;
wire  pdf ;
wire  PDG ;
wire  PDH ;
wire  PDI ;
wire  PDJ ;
wire  PDK ;
wire  PDL ;
wire  pdm ;
wire  pdn ;
wire  pdo ;
wire  QAA ;
wire  QAB ;
wire  QAC ;
wire  QAD ;
wire  QAE ;
wire  QAF ;
wire  QAG ;
wire  QAH ;
wire  QAI ;
wire  QAJ ;
wire  QBA ;
wire  QBB ;
wire  QBC ;
wire  QBD ;
wire  QBE ;
wire  QBF ;
wire  QBG ;
wire  QBH ;
wire  QBI ;
wire  QBJ ;
wire  QBK ;
wire  QBL ;
wire  QBM ;
wire  QCA ;
wire  QCB ;
wire  QCC ;
wire  qcd ;
wire  QCE ;
wire  QCF ;
wire  QCG ;
wire  QCH ;
wire  QCI ;
wire  QCJ ;
wire  QCK ;
wire  QDA ;
wire  QDB ;
wire  QDC ;
wire  QDD ;
wire  QDE ;
wire  QDF ;
wire  QDG ;
wire  QDH ;
wire  QDI ;
wire  QDJ ;
wire  QDK ;
wire  QDL ;
wire  QDM ;
wire  QDN ;
wire  QDO ;
wire  QEA ;
wire  QEB ;
wire  QEC ;
wire  QED ;
wire  QEE ;
wire  QEF ;
wire  QEG ;
wire  QEH ;
wire  QEI ;
wire  QEJ ;
wire  QEK ;
wire  QEL ;
wire  QEM ;
wire  QFA ;
wire  QFB ;
wire  QFC ;
wire  QFD ;
wire  QFE ;
wire  QFF ;
wire  QFG ;
wire  QFH ;
wire  QFI ;
wire  QFJ ;
wire  QFK ;
wire  QGA ;
wire  QGB ;
wire  QGC ;
wire  QGD ;
wire  QGE ;
wire  QGF ;
wire  QGG ;
wire  QGH ;
wire  QGI ;
wire  QGJ ;
wire  QHA ;
wire  QHB ;
wire  QHC ;
wire  QHD ;
wire  QHE ;
wire  QHF ;
wire  QHG ;
wire  qia ;
wire  qja ;
wire  qjb ;
wire  qjc ;
wire  qjd ;
wire  qje ;
wire  qjf ;
wire  qjg ;
wire  qjh ;
wire  qji ;
wire  qjj ;
wire  qjk ;
wire  qjl ;
wire  qjm ;
wire  qjn ;
wire  qjo ;
wire  qjp ;
wire  qjq ;
wire  qjr ;
wire  qjs ;
wire  qka ;
wire  qkb ;
wire  qkc ;
wire  qkd ;
wire  qke ;
wire  qkf ;
wire  qkl ;
wire  qkm ;
wire  qkn ;
wire  qko ;
wire  qkp ;
wire  qkq ;
wire  qkr ;
wire  QKS ;
wire  qkt ;
wire  qku ;
wire  qkv ;
wire  qkw ;
wire  qkx ;
wire  qky ;
wire  qla ;
wire  qlb ;
wire  qlc ;
wire  qld ;
wire  qle ;
wire  qlf ;
wire  qlg ;
wire  qlh ;
wire  qli ;
wire  qlj ;
wire  qlk ;
wire  qll ;
wire  qlm ;
wire  qln ;
wire  qlo ;
wire  qlp ;
wire  qlq ;
wire  qlr ;
wire  qls ;
wire  qlt ;
wire  qlu ;
wire  qlv ;
wire  QMA ;
wire  qmb ;
wire  qmc ;
wire  qmd ;
wire  QME ;
wire  qmf ;
wire  qmg ;
wire  qmh ;
wire  qmi ;
wire  qmj ;
wire  QMK ;
wire  QML ;
wire  QMM ;
wire  QMN ;
wire  QMO ;
wire  qna ;
wire  qne ;
wire  qnf ;
wire  qnh ;
wire  qni ;
wire  qnj ;
wire  qnk ;
wire  QNL ;
wire  QNM ;
wire  qno ;
wire  qoa ;
wire  qob ;
wire  QOC ;
wire  qod ;
wire  qoe ;
wire  qof ;
wire  qog ;
wire  qoh ;
wire  qoi ;
wire  qoj ;
wire  qol ;
wire  qpa ;
wire  qpb ;
wire  qpc ;
wire  qpd ;
wire  qqa ;
wire  qqb ;
wire  qra ;
wire  qrb ;
wire  qrc ;
wire  qrd ;
wire  qre ;
wire  qrf ;
wire  qrg ;
wire  qrh ;
wire  qri ;
wire  qrj ;
wire  qrk ;
wire  taa ;
wire  tab ;
wire  tba ;
wire  tbb ;
wire  tca ;
wire  tcb ;
wire  tda ;
wire  tdb ;
wire  tea ;
wire  teb ;
wire  tfa ;
wire  tfb ;
wire  tga ;
wire  tgb ;
wire  tha ;
wire  thb ;
wire  tia ;
wire  tib ;
wire  tka ;
wire  tkb ;
wire  tkc ;
wire  tkd ;
wire  tke ;
wire  tkf ;
wire  tkg ;
wire  tkh ;
wire  TKI ;
wire  TKJ ;
wire  TKK ;
wire  TKL ;
wire  TKM ;
wire  TKN ;
wire  TKO ;
wire  TKP ;
wire  tkq ;
wire  tkr ;
wire  tks ;
wire  tkt ;
wire  TKU ;
wire  TKV ;
wire  TKW ;
wire  TKX ;
wire  tla ;
wire  tlb ;
wire  tlc ;
wire  tld ;
wire  tle ;
wire  tlf ;
wire  tlg ;
wire  tlh ;
wire  tli ;
wire  tlj ;
wire  tlk ;
wire  tll ;
wire  tlm ;
wire  tln ;
wire  tlo ;
wire  tlp ;
wire  TNA ;
wire  TNB ;
wire  TNC ;
wire  TND ;
wire  TNE ;
wire  TNF ;
wire  toa ;
wire  TOA ;
wire  tob ;
wire  TOB ;
wire  toc ;
wire  TOC ;
wire  tod ;
wire  TOD ;
wire  toe ;
wire  TOE ;
wire  tof ;
wire  TOF ;
wire  tog ;
wire  TOG ;
wire  toh ;
wire  TOH ;
wire  toi ;
wire  TOI ;
wire  toj ;
wire  TOJ ;
wire  tok ;
wire  TOK ;
wire  tol ;
wire  TOL ;
wire  tom ;
wire  TOM ;
wire  ton ;
wire  TON ;
wire  too ;
wire  TOO ;
wire  ZZI ;
wire  ZZO ;
assign ZZI = 1'b1;
assign ZZO = 1'b0;
assign fea = ~FEA;  //complement 
assign EAA =  AEA & AFA  ; 
assign eaa = ~EAA;  //complement 
assign eba =  aea & afa  ; 
assign EBA = ~eba;  //complement 
assign aea = ~AEA;  //complement 
assign aeb = ~AEB;  //complement 
assign aca = ~ACA;  //complement 
assign acb = ~ACB;  //complement 
assign qnf = ~QNF;  //complement 
assign EAB =  AEB & AFB  ; 
assign eab = ~EAB;  //complement 
assign ebb =  aeb & afb  ; 
assign EBB = ~ebb;  //complement 
assign afa = ~AFA;  //complement 
assign afb = ~AFB;  //complement 
assign ada = ~ADA;  //complement 
assign adb = ~ADB;  //complement 
assign fad = ~FAD;  //complement 
assign fac = ~FAC;  //complement 
assign JBA =  aca & acb & acc & acd & ace & acf  ; 
assign jba = ~JBA;  //complement  
assign JCA =  ada & adb  ; 
assign jca = ~JCA;  //complement 
assign QMA = ~qma;  //complement 
assign ECB =  FEB & fab  |  feb & FAB  ; 
assign ecb = ~ECB;  //complement 
assign qne = ~QNE;  //complement 
assign qka = ~QKA;  //complement 
assign qjb = ~QJB;  //complement 
assign qjc = ~QJC;  //complement 
assign qje = ~QJE;  //complement 
assign qjf = ~QJF;  //complement 
assign aha = ~AHA;  //complement 
assign ahb = ~AHB;  //complement 
assign aga = ~AGA;  //complement 
assign agb = ~AGB;  //complement 
assign qkb = ~QKB;  //complement 
assign qjj = ~QJJ;  //complement 
assign JDD =  ahc & ahb & aha  ; 
assign jdd = ~JDD;  //complement 
assign pdb = ~PDB;  //complement 
assign QBB = ~qbb;  //complement 
assign feb = ~FEB;  //complement 
assign qjd = ~QJD;  //complement 
assign aka = ~AKA;  //complement 
assign akb = ~AKB;  //complement 
assign fab = ~FAB;  //complement 
assign JDC =  ahb & aha  ; 
assign jdc = ~JDC;  //complement 
assign aia = ~AIA;  //complement 
assign aib = ~AIB;  //complement 
assign aja = ~AJA;  //complement 
assign ajb = ~AJB;  //complement 
assign ala = ~ALA;  //complement 
assign alb = ~ALB;  //complement 
assign ama = ~AMA;  //complement 
assign amb = ~AMB;  //complement 
assign ana = ~ANA;  //complement 
assign anb = ~ANB;  //complement 
assign aoa = ~AOA;  //complement 
assign aob = ~AOB;  //complement 
assign bfa = ~BFA;  //complement 
assign bfb = ~BFB;  //complement 
assign bha = ~BHA;  //complement 
assign bhb = ~BHB;  //complement 
assign BEA = ~bea;  //complement 
assign BEB = ~beb;  //complement 
assign bga = ~BGA;  //complement 
assign bgb = ~BGB;  //complement 
assign tla = ~TLA;  //complement 
assign tlb = ~TLB;  //complement 
assign tlc = ~TLC;  //complement 
assign tld = ~TLD;  //complement 
assign QBA = ~qba;  //complement 
assign QDA = ~qda;  //complement 
assign qmb = ~QMB;  //complement 
assign qmd = ~QMD;  //complement 
assign qmc = ~QMC;  //complement 
assign haa = ~HAA;  //complement 
assign kdd =  gdd & hdd  |  GDD & HDD  ; 
assign KDD = ~kdd;  //complement 
assign kdh =  gdh & hdd  |  GDH & HDD  ; 
assign KDH = ~kdh;  //complement 
assign ldd = ~LDD;  //complement 
assign ldh = ~LDH;  //complement 
assign GCH = ~gch;  //complement 
assign QAA = ~qaa;  //complement 
assign QCA = ~qca;  //complement 
assign QFA = ~qfa;  //complement 
assign QEA = ~qea;  //complement 
assign qja = ~QJA;  //complement 
assign odc = ~ODC;  //complement 
assign oda = ~ODA;  //complement 
assign odb = ~ODB;  //complement 
assign hea = ~HEA;  //complement 
assign khd =  ghd & hhd  |  GHD & HHD  ; 
assign KHD = ~khd;  //complement 
assign khh =  ghh & hhd  |  GHH & HHD  ; 
assign KHH = ~khh;  //complement 
assign jfa =  qaa & qba & qca & qda  ; 
assign JFA = ~jfa;  //complement  
assign jga =  qaa & qia  ; 
assign JGA = ~jga;  //complement 
assign lea = ~LEA;  //complement 
assign lee = ~LEE;  //complement 
assign lhd = ~LHD;  //complement 
assign lhh = ~LHH;  //complement 
assign GGH = ~ggh;  //complement 
assign oea = ~OEA;  //complement 
assign oeb = ~OEB;  //complement 
assign oec = ~OEC;  //complement 
assign bbz = ~BBZ;  //complement 
assign pam = ~PAM;  //complement 
assign hia = ~HIA;  //complement 
assign kld =  gld & hld  |  GLD & HLD  ; 
assign KLD = ~kld;  //complement 
assign klh =  glh & hld  |  GLH & HLD  ; 
assign KLH = ~klh;  //complement 
assign lia = ~LIA;  //complement 
assign lie = ~LIE;  //complement 
assign lld = ~LLD;  //complement 
assign llh = ~LLH;  //complement 
assign GKH = ~gkh;  //complement 
assign lma = ~LMA;  //complement 
assign lme = ~LME;  //complement 
assign hma = ~HMA;  //complement 
assign aaa = ~AAA;  //complement 
assign aab = ~AAB;  //complement 
assign abb = ~ABB;  //complement 
assign BAC = ~bac;  //complement 
assign bcc = ~BCC;  //complement 
assign GBF = ~gbf;  //complement 
assign GBG = ~gbg;  //complement 
assign GBH = ~gbh;  //complement 
assign CAA =  BAD & BCD & tka  |  BAE & BCE & TKA  ; 
assign caa = ~CAA;  //complement 
assign daa =  bad & bcd & tka  |  bae & bce & TKA  ; 
assign DAA = ~daa;  //complement 
assign bad = ~BAD;  //complement 
assign bae = ~BAE;  //complement 
assign bcd = ~BCD;  //complement 
assign bce = ~BCE;  //complement 
assign hdd = ~HDD;  //complement 
assign CDD =  BAS & BCS & tka  |  BAT & BCT & TKA  ; 
assign cdd = ~CDD;  //complement 
assign ddd =  bas & bcs & tka  |  bat & bct & TKA  ; 
assign DDD = ~ddd;  //complement 
assign oaa = ~OAA;  //complement 
assign oab = ~OAB;  //complement 
assign GFF = ~gff;  //complement 
assign GFG = ~gfg;  //complement 
assign GFH = ~gfh;  //complement 
assign CEA =  BAT & BCT & tkq  |  BAU & BCU & TKQ  ; 
assign cea = ~CEA;  //complement 
assign dea =  bat & bct & tkq  |  bau & bcu & TKQ  ; 
assign DEA = ~dea;  //complement 
assign bat = ~BAT;  //complement 
assign bau = ~BAU;  //complement 
assign bct = ~BCT;  //complement 
assign bcu = ~BCU;  //complement 
assign MAQ =  LEA & pae  |  LEE & PAE  ; 
assign maq = ~MAQ;  //complement 
assign MAR =  LEB & pae  |  LEF & PAE  ; 
assign mar = ~MAR;  //complement 
assign hhd = ~HHD;  //complement 
assign CHD =  BBI & BDI & tki  |  BBJ & BDJ & TKI  ; 
assign chd = ~CHD;  //complement 
assign dhd =  bbi & bdi & tki  |  bbj & bdj & TKI  ; 
assign DHD = ~dhd;  //complement 
assign oaq = ~OAQ;  //complement 
assign oar = ~OAR;  //complement 
assign GJF = ~gjf;  //complement 
assign GJG = ~gjg;  //complement 
assign GJH = ~gjh;  //complement 
assign CIA =  BBJ & BDJ & tku  |  BBK & BDK & TKU  ; 
assign cia = ~CIA;  //complement 
assign dia =  bbj & bdj & tku  |  bbk & bdk & TKU  ; 
assign DIA = ~dia;  //complement 
assign bbj = ~BBJ;  //complement 
assign bbk = ~BBK;  //complement 
assign bdj = ~BDJ;  //complement 
assign bdk = ~BDK;  //complement 
assign MBI =  LIA & pai  |  LIE & PAI  ; 
assign mbi = ~MBI;  //complement 
assign MBJ =  LIB & pai  |  LIF & PAI  ; 
assign mbj = ~MBJ;  //complement 
assign hld = ~HLD;  //complement 
assign CLD =  BBY & BDY & tki  |  BBZ & BDZ & TKI  ; 
assign cld = ~CLD;  //complement 
assign dld =  bby & bdy & tki  |  bbz & bdz & TKI  ; 
assign DLD = ~dld;  //complement 
assign obi = ~OBI;  //complement 
assign obj = ~OBJ;  //complement 
assign MBY =  LMA & pam  |  LME & PAM  ; 
assign mby = ~MBY;  //complement 
assign GMF = ~gmf;  //complement 
assign gmb = ~GMB;  //complement 
assign CMA =  BBZ & BDZ & tki  ; 
assign cma = ~CMA;  //complement 
assign dma =  bbz & bdz & tki  |  TKI  ; 
assign DMA = ~dma;  //complement 
assign bdz = ~BDZ;  //complement 
assign fec = ~FEC;  //complement 
assign EAC =  AEC & AFC  ; 
assign eac = ~EAC;  //complement 
assign ebc =  aec & afc  ; 
assign EBC = ~ebc;  //complement 
assign aec = ~AEC;  //complement 
assign aed = ~AED;  //complement 
assign acc = ~ACC;  //complement 
assign acd = ~ACD;  //complement 
assign fed = ~FED;  //complement 
assign EAD =  AED & AFD  ; 
assign ead = ~EAD;  //complement 
assign ebd =  aed & afd  ; 
assign EBD = ~ebd;  //complement 
assign afc = ~AFC;  //complement 
assign afd = ~AFD;  //complement 
assign adc = ~ADC;  //complement 
assign add = ~ADD;  //complement 
assign fae = ~FAE;  //complement 
assign JCB =  adc & add & ade & adf & adg  ; 
assign jcb = ~JCB;  //complement  
assign jgb =  qka & qkb & qkc & qkd  ; 
assign JGB = ~jgb;  //complement 
assign jgd =  qka & qkc  ; 
assign JGD = ~jgd;  //complement 
assign jge =  qka & qkd  ; 
assign JGE = ~jge;  //complement 
assign ECC =  FEC & fac  |  fec & FAC  ; 
assign ecc = ~ECC;  //complement 
assign ECD =  FED & fad  |  fed & FAD  ; 
assign ecd = ~ECD;  //complement 
assign EGB =  FAE  ; 
assign egb = ~EGB;  //complement 
assign QDB = ~qdb;  //complement 
assign QBC = ~qbc;  //complement 
assign QDC = ~qdc;  //complement 
assign ahc = ~AHC;  //complement 
assign ahd = ~AHD;  //complement 
assign agc = ~AGC;  //complement 
assign agd = ~AGD;  //complement 
assign qkc = ~QKC;  //complement 
assign oga = ~OGA;  //complement 
assign ogb = ~OGB;  //complement 
assign ogc = ~OGC;  //complement 
assign JDF =  aha & ahb & ahc & ahd & ahe  ; 
assign jdf = ~JDF;  //complement  
assign JDE =  aha & ahb & ahc & ahd  ; 
assign jde = ~JDE;  //complement 
assign pdc = ~PDC;  //complement 
assign pdd = ~PDD;  //complement 
assign qkd = ~QKD;  //complement 
assign QAB = ~qab;  //complement 
assign QEB = ~qeb;  //complement 
assign QFB = ~qfb;  //complement 
assign QCB = ~qcb;  //complement 
assign akc = ~AKC;  //complement 
assign akd = ~AKD;  //complement 
assign QAC = ~qac;  //complement 
assign QEC = ~qec;  //complement 
assign QFC = ~qfc;  //complement 
assign QCC = ~qcc;  //complement 
assign aic = ~AIC;  //complement 
assign aid = ~AID;  //complement 
assign ajc = ~AJC;  //complement 
assign ajd = ~AJD;  //complement 
assign alc = ~ALC;  //complement 
assign ald = ~ALD;  //complement 
assign amc = ~AMC;  //complement 
assign amd = ~AMD;  //complement 
assign anc = ~ANC;  //complement 
assign andd  = ~ANDD ;  //complement 
assign aoc = ~AOC;  //complement 
assign aod = ~AOD;  //complement 
assign bfc = ~BFC;  //complement 
assign bfd = ~BFD;  //complement 
assign bhc = ~BHC;  //complement 
assign bhd = ~BHD;  //complement 
assign BEC = ~bec;  //complement 
assign BED = ~bed;  //complement 
assign bgc = ~BGC;  //complement 
assign bgd = ~BGD;  //complement 
assign kaa =  gaa & haa  |  GAA & HAA  ; 
assign KAA = ~kaa;  //complement 
assign kab =  gab & hab  |  GAB & HAB  ; 
assign KAB = ~kab;  //complement 
assign qpa = ~QPA;  //complement 
assign oma = ~OMA;  //complement 
assign hab = ~HAB;  //complement 
assign kdc =  gdc & hdc  |  GDC & HDC  ; 
assign KDC = ~kdc;  //complement 
assign kdg =  gdg & hdc  |  GDG & HDC  ; 
assign KDG = ~kdg;  //complement 
assign ldc = ~LDC;  //complement 
assign ldg = ~LDG;  //complement 
assign laa = ~LAA;  //complement 
assign lab = ~LAB;  //complement 
assign GCF = ~gcf;  //complement 
assign GCG = ~gcg;  //complement 
assign keb =  geb & heb  |  GEB & HEB  ; 
assign KEB = ~keb;  //complement 
assign kef =  gef & heb  |  GEF & HEB  ; 
assign KEF = ~kef;  //complement 
assign ndb =  hee  |  hff  ; 
assign NDB = ~ndb;  //complement 
assign PAI = ~pai;  //complement 
assign heb = ~HEB;  //complement 
assign khc =  ghc & hhc  |  GHC & HHC  ; 
assign KHC = ~khc;  //complement 
assign khg =  ghg & hhc  |  GHG & HHC  ; 
assign KHG = ~khg;  //complement 
assign neb =  hie  |  hjf  ; 
assign NEB = ~neb;  //complement 
assign leb = ~LEB;  //complement 
assign lef = ~LEF;  //complement 
assign lhc = ~LHC;  //complement 
assign lhg = ~LHG;  //complement 
assign GGF = ~ggf;  //complement 
assign GGG = ~ggg;  //complement 
assign kib =  gib & hib  |  GIB & HIB  ; 
assign KIB = ~kib;  //complement 
assign kif =  gif & hib  |  GIF & HIB  ; 
assign KIF = ~kif;  //complement 
assign pal = ~PAL;  //complement 
assign hib = ~HIB;  //complement 
assign klc =  glc & hlc  |  GLC & HLC  ; 
assign KLC = ~klc;  //complement 
assign klg =  glg & hlc  |  GLG & HLC  ; 
assign KLG = ~klg;  //complement 
assign lib = ~LIB;  //complement 
assign lif = ~LIF;  //complement 
assign llc = ~LLC;  //complement 
assign llg = ~LLG;  //complement 
assign GKF = ~gkf;  //complement 
assign GKG = ~gkg;  //complement 
assign aac = ~AAC;  //complement 
assign aad = ~AAD;  //complement 
assign abc = ~ABC;  //complement 
assign abd = ~ABD;  //complement 
assign BAB = ~bab;  //complement 
assign bcb = ~BCB;  //complement 
assign gbb = ~GBB;  //complement 
assign gbc = ~GBC;  //complement 
assign gbd = ~GBD;  //complement 
assign CAB =  BAE & BCE & tkb  |  BAF & BCF & TKB  ; 
assign cab = ~CAB;  //complement 
assign dab =  bae & bce & tkb  |  baf & bcf & TKB  ; 
assign DAB = ~dab;  //complement 
assign oao = ~OAO;  //complement 
assign oap = ~OAP;  //complement 
assign MAO =  LDC & pad  |  LDG & PAD  ; 
assign mao = ~MAO;  //complement 
assign MAP =  LDD & pad  |  LDH & PAD  ; 
assign map = ~MAP;  //complement 
assign hdc = ~HDC;  //complement 
assign CDC =  BAR & BCR & tkb  |  BAS & BCS & TKB  ; 
assign cdc = ~CDC;  //complement 
assign ddc =  bar & bcr & tkb  |  bas & bcs & TKB  ; 
assign DDC = ~ddc;  //complement 
assign bar = ~BAR;  //complement 
assign bas = ~BAS;  //complement 
assign bcs = ~BCS;  //complement 
assign gfb = ~GFB;  //complement 
assign gfc = ~GFC;  //complement 
assign gfd = ~GFD;  //complement 
assign CEB =  BAU & BCU & tkr  |  BAV & BCV & TKR  ; 
assign ceb = ~CEB;  //complement 
assign deb =  bau & bcu & tkr  |  bav & bcv & TKR  ; 
assign DEB = ~deb;  //complement 
assign obg = ~OBG;  //complement 
assign obh = ~OBH;  //complement 
assign MBG =  LHC & pah  |  LHG & PAH  ; 
assign mbg = ~MBG;  //complement 
assign MBH =  LHD & pah  |  LHH & PAH  ; 
assign mbh = ~MBH;  //complement 
assign hhc = ~HHC;  //complement 
assign CHC =  BBH & BDH & tkj  |  BBI & BDI & TKJ  ; 
assign chc = ~CHC;  //complement 
assign dhc =  bbh & bdh & tkj  |  bbi & bdi & TKJ  ; 
assign DHC = ~dhc;  //complement 
assign bbh = ~BBH;  //complement 
assign bbi = ~BBI;  //complement 
assign bdh = ~BDH;  //complement 
assign bdi = ~BDI;  //complement 
assign gjb = ~GJB;  //complement 
assign gjc = ~GJC;  //complement 
assign gjd = ~GJD;  //complement 
assign CIB =  BBK & BDK & tkv  |  BBL & BDL & TKV  ; 
assign cib = ~CIB;  //complement 
assign dib =  bbk & bdk & tkv  |  bbl & bdl & TKV  ; 
assign DIB = ~dib;  //complement 
assign obw = ~OBW;  //complement 
assign obx = ~OBX;  //complement 
assign MBW =  LLC & pal  |  LLG & PAL  ; 
assign mbw = ~MBW;  //complement 
assign MBX =  LLD & pal  |  LLH & PAL  ; 
assign mbx = ~MBX;  //complement 
assign hlc = ~HLC;  //complement 
assign CLC =  BBX & BDX & tkj  |  BBY & BDY & TKJ  ; 
assign clc = ~CLC;  //complement 
assign dlc =  bbx & bdx & tkj  |  bby & bdy & TKJ  ; 
assign DLC = ~dlc;  //complement 
assign bbx = ~BBX;  //complement 
assign bby = ~BBY;  //complement 
assign bdx = ~BDX;  //complement 
assign bdy = ~BDY;  //complement 
assign oca = ~OCA;  //complement 
assign ocb = ~OCB;  //complement 
assign occ = ~OCC;  //complement 
assign ocd = ~OCD;  //complement 
assign qia = ~QIA;  //complement 
assign QGA = ~qga;  //complement 
assign ffa = ~FFA;  //complement 
assign EAE =  AEE & AFE  ; 
assign eae = ~EAE;  //complement 
assign ebe =  aee & afe  ; 
assign EBE = ~ebe;  //complement 
assign aee = ~AEE;  //complement 
assign aef = ~AEF;  //complement 
assign ace = ~ACE;  //complement 
assign acf = ~ACF;  //complement 
assign fbe = ~FBE;  //complement 
assign EAF =  AEF & AFF  ; 
assign eaf = ~EAF;  //complement 
assign ebf =  aef & aff  ; 
assign EBF = ~ebf;  //complement 
assign afe = ~AFE;  //complement 
assign aff = ~AFF;  //complement 
assign ade = ~ADE;  //complement 
assign adf = ~ADF;  //complement 
assign fbd = ~FBD;  //complement 
assign fbc = ~FBC;  //complement 
assign QBD = ~qbd;  //complement 
assign QDD = ~qdd;  //complement 
assign qrb = ~QRB;  //complement 
assign qre = ~QRE;  //complement 
assign qra = ~QRA;  //complement 
assign EDB =  FFB & fbb  |  ffb & FBB  ; 
assign edb = ~EDB;  //complement 
assign EDE =  FFB & fbf  |  ffb & FBF  ; 
assign ede = ~EDE;  //complement 
assign EDC =  FFC & fbc  |  ffc & FBC  ; 
assign edc = ~EDC;  //complement 
assign EDF =  FFC & fbg  |  ffc & FBG  ; 
assign edf = ~EDF;  //complement 
assign qrc = ~QRC;  //complement 
assign qrf = ~QRF;  //complement 
assign qrh = ~QRH;  //complement 
assign qrj = ~QRJ;  //complement 
assign qjh = ~QJH;  //complement 
assign qji = ~QJI;  //complement 
assign ahe = ~AHE;  //complement 
assign ahf = ~AHF;  //complement 
assign age = ~AGE;  //complement 
assign agf = ~AGF;  //complement 
assign qrd = ~QRD;  //complement 
assign qrg = ~QRG;  //complement 
assign qri = ~QRI;  //complement 
assign qrk = ~QRK;  //complement 
assign qjg = ~QJG;  //complement 
assign JDG =  aha & ahb & ahc & ahd & ahe & ahf  ; 
assign jdg = ~JDG;  //complement  
assign pde = ~PDE;  //complement 
assign pdf = ~PDF;  //complement 
assign qqb = ~QQB;  //complement 
assign qke = ~QKE;  //complement 
assign oka = ~OKA;  //complement 
assign ake = ~AKE;  //complement 
assign akf = ~AKF;  //complement 
assign QAD = ~qad;  //complement 
assign QED = ~qed;  //complement 
assign QFD = ~qfd;  //complement 
assign qcd = ~QCD;  //complement 
assign QHC = ~qhc;  //complement 
assign QHE = ~qhe;  //complement 
assign QHG = ~qhg;  //complement 
assign aie = ~AIE;  //complement 
assign aif = ~AIF;  //complement 
assign aje = ~AJE;  //complement 
assign ajf = ~AJF;  //complement 
assign ale = ~ALE;  //complement 
assign alf = ~ALF;  //complement 
assign ame = ~AME;  //complement 
assign amf = ~AMF;  //complement 
assign ane = ~ANE;  //complement 
assign anf = ~ANF;  //complement 
assign aoe = ~AOE;  //complement 
assign aof = ~AOF;  //complement 
assign bfe = ~BFE;  //complement 
assign bff = ~BFF;  //complement 
assign bhe = ~BHE;  //complement 
assign bhf = ~BHF;  //complement 
assign ffb = ~FFB;  //complement 
assign BEE = ~bee;  //complement 
assign BEF = ~bef;  //complement 
assign bge = ~BGE;  //complement 
assign bgf = ~BGF;  //complement 
assign tle = ~TLE;  //complement 
assign tlf = ~TLF;  //complement 
assign tlg = ~TLG;  //complement 
assign tlh = ~TLH;  //complement 
assign kac =  gac & hac  |  GAC & HAC  ; 
assign KAC = ~kac;  //complement 
assign kad =  gad & had  |  GAD & HAD  ; 
assign KAD = ~kad;  //complement 
assign PAE = ~pae;  //complement 
assign PAD = ~pad;  //complement 
assign gaa = ~GAA;  //complement 
assign gab = ~GAB;  //complement 
assign kdb =  gdb & hdb  |  GDB & HDB  ; 
assign KDB = ~kdb;  //complement 
assign kdf =  gdf & hdb  |  GDF & HDB  ; 
assign KDF = ~kdf;  //complement 
assign fbb = ~FBB;  //complement 
assign ldb = ~LDB;  //complement 
assign ldf = ~LDF;  //complement 
assign lac = ~LAC;  //complement 
assign lad = ~LAD;  //complement 
assign gcb = ~GCB;  //complement 
assign gcc = ~GCC;  //complement 
assign kec =  gec & hec  |  GEC & HEC  ; 
assign KEC = ~kec;  //complement 
assign keg =  geg & hec  |  GEG & HEC  ; 
assign KEG = ~keg;  //complement 
assign ndc =  hee  |  hff  |  hgf  ; 
assign NDC = ~ndc;  //complement 
assign PAF = ~paf;  //complement 
assign HEE = ~hee;  //complement 
assign khb =  ghb & hhb  |  GHB & HHB  ; 
assign KHB = ~khb;  //complement 
assign khf =  ghf & hhb  |  GHF & HHB  ; 
assign KHF = ~khf;  //complement 
assign nec =  hie  |  hjf  |  hkf  ; 
assign NEC = ~nec;  //complement 
assign lec = ~LEC;  //complement 
assign leg = ~LEG;  //complement 
assign lhb = ~LHB;  //complement 
assign lhf = ~LHF;  //complement 
assign ggb = ~GGB;  //complement 
assign ggc = ~GGC;  //complement 
assign kic =  gic & hic  |  GIC & HIC  ; 
assign KIC = ~kic;  //complement 
assign kig =  gig & hic  |  GIG & HIC  ; 
assign KIG = ~kig;  //complement 
assign paj = ~PAJ;  //complement 
assign HIE = ~hie;  //complement 
assign klb =  glb & hlb  |  GLB & HLB  ; 
assign KLB = ~klb;  //complement 
assign klf =  glf & hlb  |  GLF & HLB  ; 
assign KLF = ~klf;  //complement 
assign QMO = ~qmo;  //complement 
assign lic = ~LIC;  //complement 
assign lig = ~LIG;  //complement 
assign llb = ~LLB;  //complement 
assign llf = ~LLF;  //complement 
assign gkb = ~GKB;  //complement 
assign gkc = ~GKC;  //complement 
assign QHB = ~qhb;  //complement 
assign QHD = ~qhd;  //complement 
assign QHF = ~qhf;  //complement 
assign qqa = ~QQA;  //complement 
assign aae = ~AAE;  //complement 
assign aaf = ~AAF;  //complement 
assign abe = ~ABE;  //complement 
assign abf = ~ABF;  //complement 
assign CNA =  BAA & BCB & BCC  |  BAB & BCC  |  BAC  ; 
assign cna = ~CNA;  //complement 
assign baa = ~BAA;  //complement 
assign oac = ~OAC;  //complement 
assign oad = ~OAD;  //complement 
assign hac = ~HAC;  //complement 
assign gbe = ~GBE;  //complement 
assign CAC =  BAF & BCF & tkc  |  BAG & BCG & TKC  ; 
assign cac = ~CAC;  //complement 
assign dac =  baf & bcf & tkc  |  bag & bcg & TKC  ; 
assign DAC = ~dac;  //complement 
assign baf = ~BAF;  //complement 
assign BCG = ~bcg;  //complement 
assign bcf = ~BCF;  //complement 
assign hdb = ~HDB;  //complement 
assign CDB =  BAQ & BCQ & tkc  |  BAR & BCR & TKC  ; 
assign cdb = ~CDB;  //complement 
assign ddb =  baq & bcq & tkc  |  bar & bcr & TKC  ; 
assign DDB = ~ddb;  //complement 
assign baq = ~BAQ;  //complement 
assign BCR = ~bcr;  //complement 
assign hec = ~HEC;  //complement 
assign gfe = ~GFE;  //complement 
assign CEC =  BAV & BCV & tkc  |  BAW & BCW & TKC  ; 
assign cec = ~CEC;  //complement 
assign dec =  bav & bcv & tkc  |  baw & bcw & TKC  ; 
assign DEC = ~dec;  //complement 
assign bav = ~BAV;  //complement 
assign baw = ~BAW;  //complement 
assign bcv = ~BCV;  //complement 
assign bcw = ~BCW;  //complement 
assign MAS =  LEC & pae  |  LEG & PAE  ; 
assign mas = ~MAS;  //complement 
assign MAT =  LED & pae  |  LEH & PAE  ; 
assign mat = ~MAT;  //complement 
assign hhb = ~HHB;  //complement 
assign CHB =  BBG & BDG & tkk  |  BBH & BDH & TKK  ; 
assign chb = ~CHB;  //complement 
assign dhb =  bbg & bdg & tkk  |  bbh & bdh & TKK  ; 
assign DHB = ~dhb;  //complement 
assign oas = ~OAS;  //complement 
assign oat = ~OAT;  //complement 
assign hic = ~HIC;  //complement 
assign gje = ~GJE;  //complement 
assign CIC =  BBL & BDL & tkk  |  BBM & BDM & TKK  ; 
assign cic = ~CIC;  //complement 
assign dic =  bbl & bdl & tkk  |  bbm & bdm & TKK  ; 
assign DIC = ~dic;  //complement 
assign bbl = ~BBL;  //complement 
assign bbm = ~BBM;  //complement 
assign bdl = ~BDL;  //complement 
assign bdm = ~BDM;  //complement 
assign MBK =  LIC & pai  |  LIG & PAI  ; 
assign mbk = ~MBK;  //complement 
assign MBL =  LID & pai  |  LIH & PAI  ; 
assign mbl = ~MBL;  //complement 
assign hlb = ~HLB;  //complement 
assign CLB =  BBW & BDW & tkk  |  BBX & BDX & TKK  ; 
assign clb = ~CLB;  //complement 
assign dlb =  bbw & bdw & tkk  |  bbx & bdx & TKK  ; 
assign DLB = ~dlb;  //complement 
assign obk = ~OBK;  //complement 
assign obl = ~OBL;  //complement 
assign ffd = ~FFD;  //complement 
assign qpc = ~QPC;  //complement 
assign omc = ~OMC;  //complement 
assign QHA = ~qha;  //complement 
assign ffc = ~FFC;  //complement 
assign EAG =  AEG & AFG  ; 
assign eag = ~EAG;  //complement 
assign ebg =  aeg & afg  ; 
assign EBG = ~ebg;  //complement 
assign aeg = ~AEG;  //complement 
assign aeh = ~AEH;  //complement 
assign acg = ~ACG;  //complement 
assign ach = ~ACH;  //complement 
assign ffe = ~FFE;  //complement 
assign EAH =  AEH & AFH  ; 
assign eah = ~EAH;  //complement 
assign ebh =  aeh & afh  ; 
assign EBH = ~ebh;  //complement 
assign afg = ~AFG;  //complement 
assign afh = ~AFH;  //complement 
assign adg = ~ADG;  //complement 
assign adh = ~ADH;  //complement 
assign FBH = ~fbh;  //complement 
assign FBF = ~fbf;  //complement 
assign FBG = ~fbg;  //complement 
assign JBB =  acg & ach & aci & acj & ack & acl  ; 
assign jbb = ~JBB;  //complement  
assign tba = ~TBA;  //complement 
assign tbb = ~TBB;  //complement 
assign tca = ~TCA;  //complement 
assign tcb = ~TCB;  //complement 
assign EDD =  FFD & fbd  |  ffd & FBD  ; 
assign edd = ~EDD;  //complement 
assign EDG =  FFD & fbh  |  ffd & FBH  ; 
assign edg = ~EDG;  //complement 
assign EGC =  FAE & FFE  |  FBE  ; 
assign egc = ~EGC;  //complement 
assign QBE = ~qbe;  //complement 
assign QDE = ~qde;  //complement 
assign QBF = ~qbf;  //complement 
assign QDF = ~qdf;  //complement 
assign ahg = ~AHG;  //complement 
assign ahh = ~AHH;  //complement 
assign agg = ~AGG;  //complement 
assign agh = ~AGH;  //complement 
assign tga = ~TGA;  //complement 
assign tgb = ~TGB;  //complement 
assign ofa = ~OFA;  //complement 
assign ofb = ~OFB;  //complement 
assign ofc = ~OFC;  //complement 
assign JDI =  ahg & ahh  ; 
assign jdi = ~JDI;  //complement  
assign JDJ =  ahg & ahh & ahi  ; 
assign jdj = ~JDJ;  //complement 
assign PDG = ~pdg;  //complement 
assign PDH = ~pdh;  //complement 
assign qjs = ~QJS;  //complement 
assign akg = ~AKG;  //complement 
assign akh = ~AKH;  //complement 
assign QAF = ~qaf;  //complement 
assign QEF = ~qef;  //complement 
assign QFF = ~qff;  //complement 
assign QCF = ~qcf;  //complement 
assign QAE = ~qae;  //complement 
assign QEE = ~qee;  //complement 
assign QFE = ~qfe;  //complement 
assign QCE = ~qce;  //complement 
assign aig = ~AIG;  //complement 
assign aih = ~AIH;  //complement 
assign ajg = ~AJG;  //complement 
assign ajh = ~AJH;  //complement 
assign alg = ~ALG;  //complement 
assign alh = ~ALH;  //complement 
assign amg = ~AMG;  //complement 
assign amh = ~AMH;  //complement 
assign ang = ~ANG;  //complement 
assign anh = ~ANH;  //complement 
assign aog = ~AOG;  //complement 
assign aoh = ~AOH;  //complement 
assign bfg = ~BFG;  //complement 
assign bfh = ~BFH;  //complement 
assign bhg = ~BHG;  //complement 
assign bhh = ~BHH;  //complement 
assign PAH = ~pah;  //complement 
assign BEG = ~beg;  //complement 
assign BEH = ~beh;  //complement 
assign bgg = ~BGG;  //complement 
assign bgh = ~BGH;  //complement 
assign PAB = ~pab;  //complement 
assign PAC = ~pac;  //complement 
assign gac = ~GAC;  //complement 
assign taa = ~TAA;  //complement 
assign tab = ~TAB;  //complement 
assign qjk = ~QJK;  //complement 
assign qjl = ~QJL;  //complement 
assign lda = ~LDA;  //complement 
assign lde = ~LDE;  //complement 
assign gcd = ~GCD;  //complement 
assign ked =  ged & hed  |  GED & HED  ; 
assign KED = ~ked;  //complement 
assign keh =  geh & hed  |  GEH & HED  ; 
assign KEH = ~keh;  //complement 
assign nbb =  gee & gfe & gfe  |  hfe & gfe  ; 
assign NBB = ~nbb;  //complement 
assign PAG = ~pag;  //complement 
assign gee = ~GEE;  //complement 
assign ncb =  gie & gje & gje  |  hje & gje  ; 
assign NCB = ~ncb;  //complement 
assign lha = ~LHA;  //complement 
assign lhe = ~LHE;  //complement 
assign led = ~LED;  //complement 
assign leh = ~LEH;  //complement 
assign ggd = ~GGD;  //complement 
assign kid =  gid & hid  |  GID & HID  ; 
assign KID = ~kid;  //complement 
assign kih =  gih & hid  |  GIH & HID  ; 
assign KIH = ~kih;  //complement 
assign pak = ~PAK;  //complement 
assign GIB = ~gib;  //complement 
assign gic = ~GIC;  //complement 
assign QNM = ~qnm;  //complement 
assign lla = ~LLA;  //complement 
assign lle = ~LLE;  //complement 
assign lid = ~LID;  //complement 
assign lih = ~LIH;  //complement 
assign gkd = ~GKD;  //complement 
assign aag = ~AAG;  //complement 
assign aah = ~AAH;  //complement 
assign abg = ~ABG;  //complement 
assign abh = ~ABH;  //complement 
assign tkq = ~TKQ;  //complement 
assign tkr = ~TKR;  //complement 
assign tka = ~TKA;  //complement 
assign tkb = ~TKB;  //complement 
assign had = ~HAD;  //complement 
assign hbe = ~HBE;  //complement 
assign CAD =  BAG & BCG & tkd  |  BAH & BCH & TKD  ; 
assign cad = ~CAD;  //complement 
assign dad =  bag & bcg & tkd  |  bah & bch & TKD  ; 
assign DAD = ~dad;  //complement 
assign bag = ~BAG;  //complement 
assign BCH = ~bch;  //complement 
assign MAM =  LDA & pad  |  LDE & PAD  ; 
assign mam = ~MAM;  //complement 
assign MAN =  LDB & pad  |  LDF & PAD  ; 
assign man = ~MAN;  //complement 
assign hda = ~HDA;  //complement 
assign CDA =  BAP & BCP & tkd  |  BAQ & BCQ & TKD  ; 
assign cda = ~CDA;  //complement 
assign dda =  bap & bcp & tkd  |  baq & bcq & TKD  ; 
assign DDA = ~dda;  //complement 
assign bap = ~BAP;  //complement 
assign BCQ = ~bcq;  //complement 
assign hed = ~HED;  //complement 
assign HFE = ~hfe;  //complement 
assign HFF = ~hff;  //complement 
assign CED =  BAW & BCW & tkd  |  BAX & BCX & TKD  ; 
assign ced = ~CED;  //complement 
assign ded =  baw & bcw & tkd  |  bax & bcx & TKD  ; 
assign DED = ~ded;  //complement 
assign oam = ~OAM;  //complement 
assign oan = ~OAN;  //complement 
assign MBE =  LHA & pah  |  LHE & PAH  ; 
assign mbe = ~MBE;  //complement 
assign MBF =  LHB & pah  |  LHF & PAH  ; 
assign mbf = ~MBF;  //complement 
assign hha = ~HHA;  //complement 
assign CHA =  BBF & BDF & tkl  |  BBG & BDG & TKL  ; 
assign cha = ~CHA;  //complement 
assign dha =  bbf & bdf & tkl  |  bbg & bdg & TKL  ; 
assign DHA = ~dha;  //complement 
assign bbf = ~BBF;  //complement 
assign bbg = ~BBG;  //complement 
assign bdf = ~BDF;  //complement 
assign bdg = ~BDG;  //complement 
assign hid = ~HID;  //complement 
assign HJE = ~hje;  //complement 
assign HJF = ~hjf;  //complement 
assign CID =  BBM & BDM & tkl  |  BBN & BDN & TKL  ; 
assign cid = ~CID;  //complement 
assign did =  bbm & bdm & tkl  |  bbn & bdn & TKL  ; 
assign DID = ~did;  //complement 
assign obe = ~OBE;  //complement 
assign obf = ~OBF;  //complement 
assign MBU =  LLA & pal  |  LLE & PAL  ; 
assign mbu = ~MBU;  //complement 
assign MBV =  LLB & pal  |  LLF & PAL  ; 
assign mbv = ~MBV;  //complement 
assign hla = ~HLA;  //complement 
assign CLA =  BBV & BDV & tkl  |  BBW & BDW & TKL  ; 
assign cla = ~CLA;  //complement 
assign dla =  bbv & bdv & tkl  |  bbw & bdw & TKL  ; 
assign DLA = ~dla;  //complement 
assign bbv = ~BBV;  //complement 
assign bbw = ~BBW;  //complement 
assign bdv = ~BDV;  //complement 
assign bdw = ~BDW;  //complement 
assign oce = ~OCE;  //complement 
assign ocf = ~OCF;  //complement 
assign ocg = ~OCG;  //complement 
assign och = ~OCH;  //complement 
assign TKI = ~tki;  //complement 
assign TKJ = ~tkj;  //complement 
assign TKU = ~tku;  //complement 
assign TKV = ~tkv;  //complement 
assign obu = ~OBU;  //complement 
assign obv = ~OBV;  //complement 
assign fga = ~FGA;  //complement 
assign EAI =  AEI & AFI  ; 
assign eai = ~EAI;  //complement 
assign ebi =  aei & afi  ; 
assign EBI = ~ebi;  //complement 
assign aei = ~AEI;  //complement 
assign aej = ~AEJ;  //complement 
assign aci = ~ACI;  //complement 
assign acj = ~ACJ;  //complement 
assign fce = ~FCE;  //complement 
assign EAJ =  AEJ & AFJ  ; 
assign eaj = ~EAJ;  //complement 
assign ebj =  aej & afj  ; 
assign EBJ = ~ebj;  //complement 
assign afi = ~AFI;  //complement 
assign afj = ~AFJ;  //complement 
assign adi = ~ADI;  //complement 
assign adj = ~ADJ;  //complement 
assign fcd = ~FCD;  //complement 
assign fcb = ~FCB;  //complement 
assign fcc = ~FCC;  //complement 
assign JCC =  adh & adi & adj & adk & adl  ; 
assign jcc = ~JCC;  //complement  
assign tea = ~TEA;  //complement 
assign teb = ~TEB;  //complement 
assign tda = ~TDA;  //complement 
assign tdb = ~TDB;  //complement 
assign EEB =  FGB & fcb  |  fgb & FCB  ; 
assign eeb = ~EEB;  //complement 
assign EEE =  FGB & fcf  |  fgb & FCF  ; 
assign eee = ~EEE;  //complement 
assign EEC =  FGC & fcc  |  fgc & FCC  ; 
assign eec = ~EEC;  //complement 
assign EEF =  FGC & fcg  |  fgc & FCG  ; 
assign eef = ~EEF;  //complement 
assign tfa = ~TFA;  //complement 
assign tfb = ~TFB;  //complement 
assign qlc = ~QLC;  //complement 
assign qle = ~QLE;  //complement 
assign qjn = ~QJN;  //complement 
assign qjo = ~QJO;  //complement 
assign qld = ~QLD;  //complement 
assign ahi = ~AHI;  //complement 
assign ahj = ~AHJ;  //complement 
assign agi = ~AGI;  //complement 
assign agj = ~AGJ;  //complement 
assign QBG = ~qbg;  //complement 
assign QDG = ~qdg;  //complement 
assign QBH = ~qbh;  //complement 
assign QDH = ~qdh;  //complement 
assign qjm = ~QJM;  //complement 
assign JDL =  ahg & ahh & ahi & ahj & ahk  ; 
assign jdl = ~JDL;  //complement  
assign JDK =  ahg & ahh & ahi & ahj  ; 
assign jdk = ~JDK;  //complement 
assign PDI = ~pdi;  //complement 
assign PDJ = ~pdj;  //complement 
assign qlb = ~QLB;  //complement 
assign ojd = ~OJD;  //complement 
assign oje = ~OJE;  //complement 
assign ojf = ~OJF;  //complement 
assign aki = ~AKI;  //complement 
assign akj = ~AKJ;  //complement 
assign QAH = ~qah;  //complement 
assign QEH = ~qeh;  //complement 
assign QFH = ~qfh;  //complement 
assign QCH = ~qch;  //complement 
assign QAG = ~qag;  //complement 
assign QEG = ~qeg;  //complement 
assign QFG = ~qfg;  //complement 
assign QCG = ~qcg;  //complement 
assign aii = ~AII;  //complement 
assign aij = ~AIJ;  //complement 
assign aji = ~AJI;  //complement 
assign ajj = ~AJJ;  //complement 
assign ali = ~ALI;  //complement 
assign alj = ~ALJ;  //complement 
assign ami = ~AMI;  //complement 
assign amj = ~AMJ;  //complement 
assign ani = ~ANI;  //complement 
assign anj = ~ANJ;  //complement 
assign aoi = ~AOI;  //complement 
assign aoj = ~AOJ;  //complement 
assign bfi = ~BFI;  //complement 
assign bfj = ~BFJ;  //complement 
assign bhi = ~BHI;  //complement 
assign bhj = ~BHJ;  //complement 
assign fgb = ~FGB;  //complement 
assign BEI = ~bei;  //complement 
assign BEJ = ~bej;  //complement 
assign bgi = ~BGI;  //complement 
assign bgj = ~BGJ;  //complement 
assign tli = ~TLI;  //complement 
assign tlj = ~TLJ;  //complement 
assign tlk = ~TLK;  //complement 
assign tll = ~TLL;  //complement 
assign qlf = ~QLF;  //complement 
assign lba = ~LBA;  //complement 
assign lbe = ~LBE;  //complement 
assign lcd = ~LCD;  //complement 
assign lch = ~LCH;  //complement 
assign gad = ~GAD;  //complement 
assign kcd =  gcd & hcd  |  GCD & HCD  ; 
assign KCD = ~kcd;  //complement 
assign kch =  gch & hcd  |  GCH & HCD  ; 
assign KCH = ~kch;  //complement 
assign KMA =  GAE & HBE & HCE & HDE  |  GBE & HCE & HDE  |  GCE & HDE  |  GDE  ; 
assign kma = ~KMA;  //complement 
assign gce = ~GCE;  //complement 
assign oia = ~OIA;  //complement 
assign oib = ~OIB;  //complement 
assign oic = ~OIC;  //complement 
assign oid = ~OID;  //complement 
assign KPA =  HEE & HFF & HGF & HHF  ; 
assign kpa = ~KPA;  //complement  
assign lfa = ~LFA;  //complement 
assign lfe = ~LFE;  //complement 
assign lgd = ~LGD;  //complement 
assign lgh = ~LGH;  //complement 
assign ged = ~GED;  //complement 
assign kgd =  ggd & hgd  |  GGD & HGD  ; 
assign KGD = ~kgd;  //complement 
assign kgh =  ggh & hgd  |  GGH & HGD  ; 
assign KGH = ~kgh;  //complement 
assign KQB =  HIE & HJF & HKF & HLF  ; 
assign kqb = ~KQB;  //complement  
assign KNA =  GEE & HFE & HGE & HHE  |  GFE & HGE & HHE  |  GGE & HHE  |  GHE  ; 
assign kna = ~KNA;  //complement 
assign gge = ~GGE;  //complement 
assign qnh = ~QNH;  //complement 
assign qni = ~QNI;  //complement 
assign KQA =  HIE & HJF & HKF & HLF  ; 
assign kqa = ~KQA;  //complement  
assign lja = ~LJA;  //complement 
assign lje = ~LJE;  //complement 
assign lkd = ~LKD;  //complement 
assign lkh = ~LKH;  //complement 
assign gid = ~GID;  //complement 
assign kkd =  gkd & hkd  |  GKD & HKD  ; 
assign KKD = ~kkd;  //complement 
assign kkh =  gkh & hkd  |  GKH & HKD  ; 
assign KKH = ~kkh;  //complement 
assign KOA =  GIE & HJE & HKE & HLE  |  GJE & HKE & HLE  |  GKE & HLE  |  GLE  ; 
assign koa = ~KOA;  //complement 
assign gke = ~GKE;  //complement 
assign QNL = ~qnl;  //complement 
assign aai = ~AAI;  //complement 
assign aaj = ~AAJ;  //complement 
assign abi = ~ABI;  //complement 
assign abj = ~ABJ;  //complement 
assign tkc = ~TKC;  //complement 
assign tkd = ~TKD;  //complement 
assign tke = ~TKE;  //complement 
assign tkf = ~TKF;  //complement 
assign oae = ~OAE;  //complement 
assign oaf = ~OAF;  //complement 
assign MAE =  LBA & pab  |  LBE & PAB  ; 
assign mae = ~MAE;  //complement 
assign MAF =  LBB & pab  |  LBF & PAB  ; 
assign maf = ~MAF;  //complement 
assign hba = ~HBA;  //complement 
assign CBA =  BAH & BCH & tke  |  BAI & BCI & TKE  ; 
assign cba = ~CBA;  //complement 
assign dba =  bah & bch & tke  |  bai & bci & TKE  ; 
assign DBA = ~dba;  //complement 
assign bah = ~BAH;  //complement 
assign BCI = ~bci;  //complement 
assign hcd = ~HCD;  //complement 
assign hde = ~HDE;  //complement 
assign CCD =  BAO & BCO & tke  |  BAP & BCP & TKE  ; 
assign ccd = ~CCD;  //complement 
assign dcd =  bao & bco & tke  |  bap & bcp & TKE  ; 
assign DCD = ~dcd;  //complement 
assign bao = ~BAO;  //complement 
assign BCP = ~bcp;  //complement 
assign MAU =  LFA & paf  |  LFE & PAF  ; 
assign mau = ~MAU;  //complement 
assign MAV =  LFB & paf  |  LFF & PAF  ; 
assign mav = ~MAV;  //complement 
assign hfa = ~HFA;  //complement 
assign CFA =  BAX & BCX & tke  |  BAY & BCY & TKE  ; 
assign cfa = ~CFA;  //complement 
assign dfa =  bax & bcx & tke  |  bay & bcy & TKE  ; 
assign DFA = ~dfa;  //complement 
assign bax = ~BAX;  //complement 
assign bay = ~BAY;  //complement 
assign bcx = ~BCX;  //complement 
assign bcy = ~BCY;  //complement 
assign hgd = ~HGD;  //complement 
assign HHE = ~hhe;  //complement 
assign HHF = ~hhf;  //complement 
assign CGD =  BBE & BDE & tkm  |  BBF & BDF & TKM  ; 
assign cgd = ~CGD;  //complement 
assign dgd =  bbe & bde & tkm  |  bbf & bdf & TKM  ; 
assign DGD = ~dgd;  //complement 
assign oau = ~OAU;  //complement 
assign oav = ~OAV;  //complement 
assign MBM =  LJA & paj  |  LJE & PAJ  ; 
assign mbm = ~MBM;  //complement 
assign MBN =  LJB & paj  |  LJF & PAJ  ; 
assign mbn = ~MBN;  //complement 
assign hja = ~HJA;  //complement 
assign CJA =  BBN & BDN & tkm  |  BBO & BDO & TKM  ; 
assign cja = ~CJA;  //complement 
assign dja =  bbn & bdn & tkm  |  bbo & bdo & TKM  ; 
assign DJA = ~dja;  //complement 
assign bbn = ~BBN;  //complement 
assign bbo = ~BBO;  //complement 
assign bdn = ~BDN;  //complement 
assign bdo = ~BDO;  //complement 
assign hkd = ~HKD;  //complement 
assign HLE = ~hle;  //complement 
assign HLF = ~hlf;  //complement 
assign CKD =  BBU & BDU & tkm  |  BBV & BDV & TKM  ; 
assign ckd = ~CKD;  //complement 
assign dkd =  bbu & bdu & tkm  |  bbv & bdv & TKM  ; 
assign DKD = ~dkd;  //complement 
assign obm = ~OBM;  //complement 
assign obn = ~OBN;  //complement 
assign fgd = ~FGD;  //complement 
assign TKK = ~tkk;  //complement 
assign TKL = ~tkl;  //complement 
assign TKM = ~tkm;  //complement 
assign TKN = ~tkn;  //complement 
assign fgc = ~FGC;  //complement 
assign EAK =  AEK & AFK  ; 
assign eak = ~EAK;  //complement 
assign ebk =  aek & afk  ; 
assign EBK = ~ebk;  //complement 
assign aek = ~AEK;  //complement 
assign ael = ~AEL;  //complement 
assign ack = ~ACK;  //complement 
assign acl = ~ACL;  //complement 
assign fge = ~FGE;  //complement 
assign EAL =  AEL & AFL  ; 
assign eal = ~EAL;  //complement 
assign ebl =  ael & afl  ; 
assign EBL = ~ebl;  //complement 
assign afk = ~AFK;  //complement 
assign afl = ~AFL;  //complement 
assign adk = ~ADK;  //complement 
assign adl = ~ADL;  //complement 
assign FCH = ~fch;  //complement 
assign FCF = ~fcf;  //complement 
assign FCG = ~fcg;  //complement 
assign QBI = ~qbi;  //complement 
assign QDI = ~qdi;  //complement 
assign QBJ = ~qbj;  //complement 
assign QDJ = ~qdj;  //complement 
assign qkf = ~QKF;  //complement 
assign EED =  FGD & fcd  |  fgd & FCD  ; 
assign eed = ~EED;  //complement 
assign EEG =  FGD & fch  |  fgd & FCH  ; 
assign eeg = ~EEG;  //complement 
assign EGD =  FAE & FFE & FGE  |  FBE & FGE  |  FCE  ; 
assign egd = ~EGD;  //complement 
assign QMK = ~qmk;  //complement 
assign qna = ~QNA;  //complement 
assign ahk = ~AHK;  //complement 
assign ahl = ~AHL;  //complement 
assign agk = ~AGK;  //complement 
assign agl = ~AGL;  //complement 
assign QML = ~qml;  //complement 
assign oha = ~OHA;  //complement 
assign ohb = ~OHB;  //complement 
assign ohc = ~OHC;  //complement 
assign JDM =  ahg & ahh & ahi & ahj & ahk & ahl  ; 
assign jdm = ~JDM;  //complement  
assign PDK = ~pdk;  //complement 
assign PDL = ~pdl;  //complement 
assign qla = ~QLA;  //complement 
assign qjr = ~QJR;  //complement 
assign ojc = ~OJC;  //complement 
assign akk = ~AKK;  //complement 
assign akl = ~AKL;  //complement 
assign QAJ = ~qaj;  //complement 
assign QEJ = ~qej;  //complement 
assign QFJ = ~qfj;  //complement 
assign QCJ = ~qcj;  //complement 
assign QAI = ~qai;  //complement 
assign QEI = ~qei;  //complement 
assign QFI = ~qfi;  //complement 
assign QCI = ~qci;  //complement 
assign aik = ~AIK;  //complement 
assign ail = ~AIL;  //complement 
assign ajk = ~AJK;  //complement 
assign ajl = ~AJL;  //complement 
assign alk = ~ALK;  //complement 
assign all = ~ALL;  //complement 
assign amk = ~AMK;  //complement 
assign aml = ~AML;  //complement 
assign ank = ~ANK;  //complement 
assign anl = ~ANL;  //complement 
assign aok = ~AOK;  //complement 
assign aol = ~AOL;  //complement 
assign bfk = ~BFK;  //complement 
assign bfl = ~BFL;  //complement 
assign bhk = ~BHK;  //complement 
assign bhl = ~BHL;  //complement 
assign BEK = ~bek;  //complement 
assign BEL = ~bel;  //complement 
assign bgk = ~BGK;  //complement 
assign bgl = ~BGL;  //complement 
assign kbb =  gbb & hbb  |  GBB & HBB  ; 
assign KBB = ~kbb;  //complement 
assign kbf =  gbf & hbb  |  GBF & HBB  ; 
assign KBF = ~kbf;  //complement 
assign lbb = ~LBB;  //complement 
assign lbf = ~LBF;  //complement 
assign lcc = ~LCC;  //complement 
assign lcg = ~LCG;  //complement 
assign gae = ~GAE;  //complement 
assign kcc =  gcc & hcc  |  GCC & HCC  ; 
assign KCC = ~kcc;  //complement 
assign kcg =  gcg & hcc  |  GCG & HCC  ; 
assign KCG = ~kcg;  //complement 
assign KMB =  GAE & HBE & HCE & HDE  |  GBE & HCE & HDE  |  GCE & HDE  |  GDE  ; 
assign kmb = ~KMB;  //complement 
assign HCE = ~hce;  //complement 
assign kfb =  gfb & hfb  |  GFB & HFB  ; 
assign KFB = ~kfb;  //complement 
assign kff =  gff & hfb  |  GFF & HFB  ; 
assign KFF = ~kff;  //complement 
assign KPB =  HEE & HFF & HGF & HHF  ; 
assign kpb = ~KPB;  //complement  
assign lfb = ~LFB;  //complement 
assign lff = ~LFF;  //complement 
assign lgc = ~LGC;  //complement 
assign lgg = ~LGG;  //complement 
assign geb = ~GEB;  //complement 
assign gec = ~GEC;  //complement 
assign kgc =  ggc & hgc  |  GGC & HGC  ; 
assign KGC = ~kgc;  //complement 
assign kgg =  ggg & hgc  |  GGG & HGC  ; 
assign KGG = ~kgg;  //complement 
assign QMM = ~qmm;  //complement 
assign tia = ~TIA;  //complement 
assign tib = ~TIB;  //complement 
assign KNB =  GEE & HFE & HGE & HHE  |  GFE & HGE & HHE  |  GGE & HHE  |  GHE  ; 
assign knb = ~KNB;  //complement 
assign HGE = ~hge;  //complement 
assign HGF = ~hgf;  //complement 
assign kjb =  gjb & hjb  |  GJB & HJB  ; 
assign KJB = ~kjb;  //complement 
assign kjf =  gjf & hjb  |  GJF & HJB  ; 
assign KJF = ~kjf;  //complement 
assign ljb = ~LJB;  //complement 
assign ljf = ~LJF;  //complement 
assign lkc = ~LKC;  //complement 
assign lkg = ~LKG;  //complement 
assign gie = ~GIE;  //complement 
assign kkc =  gkc & hkc  |  GKC & HKC  ; 
assign KKC = ~kkc;  //complement 
assign kkg =  gkg & hkc  |  GKG & HKC  ; 
assign KKG = ~kkg;  //complement 
assign KOB =  GIE & HJE & HKE & HLE  |  GJE & HKE & HLE  |  GKE & HLE  |  GLE  ; 
assign kob = ~KOB;  //complement 
assign HKE = ~hke;  //complement 
assign HKF = ~hkf;  //complement 
assign aak = ~AAK;  //complement 
assign aal = ~AAL;  //complement 
assign abk = ~ABK;  //complement 
assign abl = ~ABL;  //complement 
assign tks = ~TKS;  //complement 
assign tkt = ~TKT;  //complement 
assign tkg = ~TKG;  //complement 
assign tkh = ~TKH;  //complement 
assign oak = ~OAK;  //complement 
assign oal = ~OAL;  //complement 
assign MAK =  LCC & pac  |  LCG & PAC  ; 
assign mak = ~MAK;  //complement 
assign MAL =  LCD & pac  |  LCH & PAC  ; 
assign mal = ~MAL;  //complement 
assign hbb = ~HBB;  //complement 
assign CBB =  BAI & BCI & tkf  |  BAJ & BCJ & TKF  ; 
assign cbb = ~CBB;  //complement 
assign dbb =  bai & bci & tkf  |  baj & bcj & TKF  ; 
assign DBB = ~dbb;  //complement 
assign bai = ~BAI;  //complement 
assign BCJ = ~bcj;  //complement 
assign hcc = ~HCC;  //complement 
assign gde = ~GDE;  //complement 
assign CCC =  BAN & BCN & tkf  |  BAO & BCO & TKF  ; 
assign ccc = ~CCC;  //complement 
assign dcc =  ban & bcn & tkf  |  bao & bco & TKF  ; 
assign DCC = ~dcc;  //complement 
assign ban = ~BAN;  //complement 
assign bcn = ~BCN;  //complement 
assign bco = ~BCO;  //complement 
assign MBC =  LGC & pag  |  LGG & PAG  ; 
assign mbc = ~MBC;  //complement 
assign MBD =  LGD & pag  |  LGH & PAG  ; 
assign mbd = ~MBD;  //complement 
assign hfb = ~HFB;  //complement 
assign CFB =  BAY & BCY & tkf  |  BAZ & BCZ & TKF  ; 
assign cfb = ~CFB;  //complement 
assign dfb =  bay & bcy & tkf  |  baz & bcz & TKF  ; 
assign DFB = ~dfb;  //complement 
assign obc = ~OBC;  //complement 
assign obd = ~OBD;  //complement 
assign hgc = ~HGC;  //complement 
assign ghe = ~GHE;  //complement 
assign CGC =  BBD & BDD & tkn  |  BBE & BDE & TKN  ; 
assign cgc = ~CGC;  //complement 
assign dgc =  bbd & bdd & tkn  |  bbe & bde & TKN  ; 
assign DGC = ~dgc;  //complement 
assign bbd = ~BBD;  //complement 
assign bbe = ~BBE;  //complement 
assign bdd = ~BDD;  //complement 
assign bde = ~BDE;  //complement 
assign MBS =  LKC & pak  |  LKG & PAK  ; 
assign mbs = ~MBS;  //complement 
assign MBT =  LKD & pak  |  LKH & PAK  ; 
assign mbt = ~MBT;  //complement 
assign hjb = ~HJB;  //complement 
assign CJB =  BBO & BDO & tkn  |  BBP & BDP & TKN  ; 
assign cjb = ~CJB;  //complement 
assign djb =  bbo & bdo & tkn  |  bbp & bdp & TKN  ; 
assign DJB = ~djb;  //complement 
assign obs = ~OBS;  //complement 
assign obt = ~OBT;  //complement 
assign hkc = ~HKC;  //complement 
assign gle = ~GLE;  //complement 
assign CKC =  BBT & BDT & tkn  |  BBU & BDU & TKN  ; 
assign ckc = ~CKC;  //complement 
assign dkc =  bbt & bdt & tkn  |  bbu & bdu & TKN  ; 
assign DKC = ~dkc;  //complement 
assign bbt = ~BBT;  //complement 
assign bbu = ~BBU;  //complement 
assign bdt = ~BDT;  //complement 
assign bdu = ~BDU;  //complement 
assign oci = ~OCI;  //complement 
assign ocj = ~OCJ;  //complement 
assign ock = ~OCK;  //complement 
assign ocl = ~OCL;  //complement 
assign TKO = ~tko;  //complement 
assign TKP = ~tkp;  //complement 
assign TKW = ~tkw;  //complement 
assign TKX = ~tkx;  //complement 
assign fhb = ~FHB;  //complement 
assign fha = ~FHA;  //complement 
assign EAM =  AEM & AFM  ; 
assign eam = ~EAM;  //complement 
assign ebm =  aem & afm  ; 
assign EBM = ~ebm;  //complement 
assign aem = ~AEM;  //complement 
assign aen = ~AEN;  //complement 
assign qlq = ~QLQ;  //complement 
assign qlu = ~QLU;  //complement 
assign acm = ~ACM;  //complement 
assign acn = ~ACN;  //complement 
assign qmi = ~QMI;  //complement 
assign qoh = ~QOH;  //complement 
assign EAN =  AEN & AFN  ; 
assign ean = ~EAN;  //complement 
assign ebn =  aen & afn  ; 
assign EBN = ~ebn;  //complement 
assign afm = ~AFM;  //complement 
assign afn = ~AFN;  //complement 
assign adm = ~ADM;  //complement 
assign adn = ~ADN;  //complement 
assign FDF = ~fdf;  //complement 
assign FDG = ~fdg;  //complement 
assign fdb = ~FDB;  //complement 
assign fdc = ~FDC;  //complement 
assign JCD =  adm & adn & ADO  ; 
assign jcd = ~JCD;  //complement 
assign JAB =  ADM & ado  ; 
assign jab = ~JAB;  //complement 
assign JBC =  acm & acn & ADO  ; 
assign jbc = ~JBC;  //complement 
assign JAA =  ACN & aco  ; 
assign jaa = ~JAA;  //complement 
assign EFB =  FHB & fdb  |  fhb & FDB  ; 
assign efb = ~EFB;  //complement 
assign EFE =  FHB & fdf  |  fhb & FDF  ; 
assign efe = ~EFE;  //complement 
assign qkn = ~QKN;  //complement 
assign qkq = ~QKQ;  //complement 
assign qoi = ~QOI;  //complement 
assign QMN = ~qmn;  //complement 
assign QBK = ~qbk;  //complement 
assign QDK = ~qdk;  //complement 
assign QBL = ~qbl;  //complement 
assign QDL = ~qdl;  //complement 
assign qkm = ~QKM;  //complement 
assign qkp = ~QKP;  //complement 
assign qko = ~QKO;  //complement 
assign qkr = ~QKR;  //complement 
assign ahm = ~AHM;  //complement 
assign ahn = ~AHN;  //complement 
assign agm = ~AGM;  //complement 
assign agn = ~AGN;  //complement 
assign qkl = ~QKL;  //complement 
assign qpb = ~QPB;  //complement 
assign omb = ~OMB;  //complement 
assign JDO =  ahm & ahn  ; 
assign jdo = ~JDO;  //complement  
assign pdm = ~PDM;  //complement 
assign TNA = ~tna;  //complement 
assign TNB = ~tnb;  //complement 
assign TNC = ~tnc;  //complement 
assign qjq = ~QJQ;  //complement 
assign ojb = ~OJB;  //complement 
assign akm = ~AKM;  //complement 
assign akn = ~AKN;  //complement 
assign JEC =  aio & qne & QLR & QLD  ; 
assign jec = ~JEC;  //complement  
assign JEB =  ain & AIO & qne & qlv  ; 
assign jeb = ~JEB;  //complement 
assign QCK = ~qck;  //complement 
assign QEK = ~qek;  //complement 
assign QFK = ~qfk;  //complement 
assign QEL = ~qel;  //complement 
assign aim = ~AIM;  //complement 
assign ain = ~AIN;  //complement 
assign ajm = ~AJM;  //complement 
assign ajn = ~AJN;  //complement 
assign alm = ~ALM;  //complement 
assign aln = ~ALN;  //complement 
assign amn = ~AMN;  //complement 
assign amm = ~AMM;  //complement 
assign anm = ~ANM;  //complement 
assign ann = ~ANN;  //complement 
assign aom = ~AOM;  //complement 
assign aon = ~AON;  //complement 
assign bfm = ~BFM;  //complement 
assign bfn = ~BFN;  //complement 
assign bhm = ~BHM;  //complement 
assign bhn = ~BHN;  //complement 
assign qlv = ~QLV;  //complement 
assign qlr = ~QLR;  //complement 
assign BEM = ~bem;  //complement 
assign BEN = ~ben;  //complement 
assign bgm = ~BGM;  //complement 
assign bgn = ~BGN;  //complement 
assign tlm = ~TLM;  //complement 
assign tln = ~TLN;  //complement 
assign tlo = ~TLO;  //complement 
assign tlp = ~TLP;  //complement 
assign kbc =  gbc & hbc  |  GBC & HBC  ; 
assign KBC = ~kbc;  //complement 
assign kbg =  gbg & hbc  |  GBG & HBC  ; 
assign KBG = ~kbg;  //complement 
assign lbc = ~LBC;  //complement 
assign lbg = ~LBG;  //complement 
assign lcb = ~LCB;  //complement 
assign lcf = ~LCF;  //complement 
assign TOA =  PBA  |  PCA  ; 
assign toa = ~TOA;  //complement 
assign TOC =  PBA  |  PCA  ; 
assign toc = ~TOC;  //complement 
assign kcb =  gcb & hcb  |  GCB & HCB  ; 
assign KCB = ~kcb;  //complement 
assign kcf =  gcf & hcb  |  GCF & HCB  ; 
assign KCF = ~kcf;  //complement 
assign pba = ~PBA;  //complement 
assign hcb = ~HCB;  //complement 
assign kfc =  gfc & hfc  |  GFC & HFC  ; 
assign KFC = ~kfc;  //complement 
assign kfg =  gfg & hfc  |  GFG & HFC  ; 
assign KFG = ~kfg;  //complement 
assign nbc =  ZZI & gee & gfe & gge  |  hfe & gfe & gge  |  hge & gge  ; 
assign NBC = ~nbc;  //complement 
assign lfc = ~LFC;  //complement 
assign lfg = ~LFG;  //complement 
assign lgb = ~LGB;  //complement 
assign lgf = ~LGF;  //complement 
assign GEF = ~gef;  //complement 
assign GEG = ~geg;  //complement 
assign kgb =  ggb & hgb  |  GGB & HGB  ; 
assign KGB = ~kgb;  //complement 
assign kgf =  ggf & hgb  |  GGF & HGB  ; 
assign KGF = ~kgf;  //complement 
assign ncc =  ZZI & gie & gje & gke  |  hje & gje & gke  |  hke & gke  ; 
assign NCC = ~ncc;  //complement 
assign toi =  pba & pca  ; 
assign TOI = ~toi;  //complement 
assign toj =  pba & pca  ; 
assign TOJ = ~toj;  //complement 
assign tog =  pba & pca  ; 
assign TOG = ~tog;  //complement 
assign hgb = ~HGB;  //complement 
assign kjc =  gjc & hjc  |  GJC & HJC  ; 
assign KJC = ~kjc;  //complement 
assign kjg =  gjg & hjc  |  GJG & HJC  ; 
assign KJG = ~kjg;  //complement 
assign toh =  pba & pca  ; 
assign TOH = ~toh;  //complement 
assign tom =  pba & pca  ; 
assign TOM = ~tom;  //complement 
assign toe =  pba & pca  ; 
assign TOE = ~toe;  //complement 
assign ljc = ~LJC;  //complement 
assign ljg = ~LJG;  //complement 
assign lkb = ~LKB;  //complement 
assign lkf = ~LKF;  //complement 
assign GIF = ~gif;  //complement 
assign GIG = ~gig;  //complement 
assign kkb =  gkb & hkb  |  GKB & HKB  ; 
assign KKB = ~kkb;  //complement 
assign kkf =  gkf & hkb  |  GKF & HKB  ; 
assign KKF = ~kkf;  //complement 
assign hkb = ~HKB;  //complement 
assign aam = ~AAM;  //complement 
assign aan = ~AAN;  //complement 
assign abm = ~ABM;  //complement 
assign abn = ~ABN;  //complement 
assign MAG =  LBC & pab  |  LBG & PAB  ; 
assign mag = ~MAG;  //complement 
assign MAH =  LBD & pab  |  LBH & PAB  ; 
assign mah = ~MAH;  //complement 
assign hbc = ~HBC;  //complement 
assign CBC =  BAJ & BCJ & tkg  |  BAK & BCK & TKG  ; 
assign cbc = ~CBC;  //complement 
assign dbc =  baj & bcj & tkg  |  bak & bck & TKG  ; 
assign DBC = ~dbc;  //complement 
assign baj = ~BAJ;  //complement 
assign bak = ~BAK;  //complement 
assign bck = ~BCK;  //complement 
assign gdb = ~GDB;  //complement 
assign gdc = ~GDC;  //complement 
assign gdd = ~GDD;  //complement 
assign CCB =  BAM & BCM & tkt  |  BAN & BCN & TKT  ; 
assign ccb = ~CCB;  //complement 
assign dcb =  bam & bcm & tkt  |  ban & bcn & TKT  ; 
assign DCB = ~dcb;  //complement 
assign oag = ~OAG;  //complement 
assign oah = ~OAH;  //complement 
assign MAW =  LFC & paf  |  LFG & PAF  ; 
assign maw = ~MAW;  //complement 
assign MAX =  LFD & paf  |  LFH & PAF  ; 
assign max = ~MAX;  //complement 
assign hfc = ~HFC;  //complement 
assign CFC =  BAZ & BCZ & tkg  |  BBA & BDA & TKG  ; 
assign cfc = ~CFC;  //complement 
assign dfc =  baz & bcz & tkg  |  bba & bda & TKG  ; 
assign DFC = ~dfc;  //complement 
assign baz = ~BAZ;  //complement 
assign bba = ~BBA;  //complement 
assign bcz = ~BCZ;  //complement 
assign bda = ~BDA;  //complement 
assign ghc = ~GHC;  //complement 
assign ghd = ~GHD;  //complement 
assign CGB =  BBC & BDC & tkx  |  BBD & BDD & TKX  ; 
assign cgb = ~CGB;  //complement 
assign dgb =  bbc & bdc & tkx  |  bbd & bdd & TKX  ; 
assign DGB = ~dgb;  //complement 
assign oaw = ~OAW;  //complement 
assign oax = ~OAX;  //complement 
assign MBO =  LJC & paj  |  LJG & PAJ  ; 
assign mbo = ~MBO;  //complement 
assign MBP =  LJD & paj  |  LJH & PAJ  ; 
assign mbp = ~MBP;  //complement 
assign hjc = ~HJC;  //complement 
assign CJC =  BBP & BDP & tko  |  BBQ & BDQ & TKO  ; 
assign cjc = ~CJC;  //complement 
assign djc =  bbp & bdp & tko  |  bbq & bdq & TKO  ; 
assign DJC = ~djc;  //complement 
assign bbp = ~BBP;  //complement 
assign bbq = ~BBQ;  //complement 
assign bdp = ~BDP;  //complement 
assign bdq = ~BDQ;  //complement 
assign glb = ~GLB;  //complement 
assign glc = ~GLC;  //complement 
assign gld = ~GLD;  //complement 
assign CKB =  BBS & BDS & tko  |  BBT & BDT & TKO  ; 
assign ckb = ~CKB;  //complement 
assign dkb =  bbs & bds & tko  |  bbt & bdt & TKO  ; 
assign DKB = ~dkb;  //complement 
assign obo = ~OBO;  //complement 
assign obp = ~OBP;  //complement 
assign qlp = ~QLP;  //complement 
assign ghb = ~GHB;  //complement 
assign afp = ~AFP;  //complement 
assign fhc = ~FHC;  //complement 
assign ola = ~OLA;  //complement 
assign fia = ~FIA;  //complement 
assign EAO =  AEO & AFO  ; 
assign eao = ~EAO;  //complement 
assign ebo =  aeo & afo  ; 
assign EBO = ~ebo;  //complement 
assign aeo = ~AEO;  //complement 
assign aep = ~AEP;  //complement 
assign qlo = ~QLO;  //complement 
assign qls = ~QLS;  //complement 
assign aco = ~ACO;  //complement 
assign acp = ~ACP;  //complement 
assign qmf = ~QMF;  //complement 
assign qmh = ~QMH;  //complement 
assign qoa = ~QOA;  //complement 
assign qoe = ~QOE;  //complement 
assign qkt = ~QKT;  //complement 
assign qkv = ~QKV;  //complement 
assign qkx = ~QKX;  //complement 
assign qlh = ~QLH;  //complement 
assign afo = ~AFO;  //complement 
assign ado = ~ADO;  //complement 
assign adp = ~ADP;  //complement 
assign qmg = ~QMG;  //complement 
assign qod = ~QOD;  //complement 
assign qob = ~QOB;  //complement 
assign qof = ~QOF;  //complement 
assign qku = ~QKU;  //complement 
assign qkw = ~QKW;  //complement 
assign qky = ~QKY;  //complement 
assign qli = ~QLI;  //complement 
assign QKS = ~qks;  //complement 
assign QME = ~qme;  //complement 
assign EFC =  FHC & fdc  |  fhc & FDC  ; 
assign efc = ~EFC;  //complement 
assign EFF =  FHC & fdg  |  fhc & FDG  ; 
assign eff = ~EFF;  //complement 
assign qlk = ~QLK;  //complement 
assign qlm = ~QLM;  //complement 
assign QGD = ~qgd;  //complement 
assign QGF = ~qgf;  //complement 
assign QGH = ~qgh;  //complement 
assign QGJ = ~qgj;  //complement 
assign QGC = ~qgc;  //complement 
assign QGE = ~qge;  //complement 
assign QGG = ~qgg;  //complement 
assign QGI = ~qgi;  //complement 
assign aho = ~AHO;  //complement 
assign ahp = ~AHP;  //complement 
assign ago = ~AGO;  //complement 
assign qlg = ~QLG;  //complement 
assign qll = ~QLL;  //complement 
assign qpd = ~QPD;  //complement 
assign omd = ~OMD;  //complement 
assign pdo = ~PDO;  //complement 
assign pdn = ~PDN;  //complement 
assign TND = ~tnd;  //complement 
assign TNE = ~tne;  //complement 
assign TNF = ~tnf;  //complement 
assign qjp = ~QJP;  //complement 
assign oja = ~OJA;  //complement 
assign ako = ~AKO;  //complement 
assign jea = ~JEA;  //complement 
assign QEM = ~qem;  //complement 
assign QBM = ~qbm;  //complement 
assign QDM = ~qdm;  //complement 
assign QDO = ~qdo;  //complement 
assign QDN = ~qdn;  //complement 
assign QGB = ~qgb;  //complement 
assign qlj = ~QLJ;  //complement 
assign aio = ~AIO;  //complement 
assign aip = ~AIP;  //complement 
assign ajo = ~AJO;  //complement 
assign ajp = ~AJP;  //complement 
assign alo = ~ALO;  //complement 
assign alp = ~ALP;  //complement 
assign amo = ~AMO;  //complement 
assign amp = ~AMP;  //complement 
assign anp = ~ANP;  //complement 
assign aoo = ~AOO;  //complement 
assign bfo = ~BFO;  //complement 
assign bfp = ~BFP;  //complement 
assign bho = ~BHO;  //complement 
assign bhp = ~BHP;  //complement 
assign ano = ~ANO;  //complement 
assign BEO = ~beo;  //complement 
assign BEP = ~bep;  //complement 
assign bgo = ~BGO;  //complement 
assign bgp = ~BGP;  //complement 
assign aop = ~AOP;  //complement 
assign kbd =  gbd & hbd  |  GBD & HBD  ; 
assign KBD = ~kbd;  //complement 
assign kbh =  gbh & hbd  |  GBH & HBD  ; 
assign KBH = ~kbh;  //complement 
assign akp = ~AKP;  //complement 
assign lca = ~LCA;  //complement 
assign lce = ~LCE;  //complement 
assign lbd = ~LBD;  //complement 
assign lbh = ~LBH;  //complement 
assign TOB =  PBA  |  PCA  ; 
assign tob = ~TOB;  //complement 
assign qln = ~QLN;  //complement 
assign qlt = ~QLT;  //complement 
assign qno = ~QNO;  //complement 
assign PCA = ~pca;  //complement 
assign hca = ~HCA;  //complement 
assign kfd =  gfd & hfd  |  GFD & HFD  ; 
assign KFD = ~kfd;  //complement 
assign kfh =  gfh & hfd  |  GFH & HFD  ; 
assign KFH = ~kfh;  //complement 
assign qoj = ~QOJ;  //complement 
assign lga = ~LGA;  //complement 
assign lge = ~LGE;  //complement 
assign lfd = ~LFD;  //complement 
assign lfh = ~LFH;  //complement 
assign GEH = ~geh;  //complement 
assign QOC = ~qoc;  //complement 
assign qol = ~QOL;  //complement 
assign tok =  pba & pca  ; 
assign TOK = ~tok;  //complement 
assign tol =  pba & pca  ; 
assign TOL = ~tol;  //complement 
assign tof =  pba & pca  ; 
assign TOF = ~tof;  //complement 
assign hga = ~HGA;  //complement 
assign kjd =  gjd & hjd  |  GJD & HJD  ; 
assign KJD = ~kjd;  //complement 
assign kjh =  gjh & hjd  |  GJH & HJD  ; 
assign KJH = ~kjh;  //complement 
assign tod =  pba & pca  ; 
assign TOD = ~tod;  //complement 
assign ton =  pba & pca  ; 
assign TON = ~ton;  //complement 
assign too =  pba & pca  ; 
assign TOO = ~too;  //complement 
assign lka = ~LKA;  //complement 
assign lke = ~LKE;  //complement 
assign ljd = ~LJD;  //complement 
assign ljh = ~LJH;  //complement 
assign GIH = ~gih;  //complement 
assign qmj = ~QMJ;  //complement 
assign jed = ~JED;  //complement 
assign qnj = ~QNJ;  //complement 
assign qnk = ~QNK;  //complement 
assign hka = ~HKA;  //complement 
assign qog = ~QOG;  //complement 
assign agp = ~AGP;  //complement 
assign JEE =  AKN & AKO  |  QMO  ; 
assign jee = ~JEE;  //complement 
assign tha = ~THA;  //complement 
assign thb = ~THB;  //complement 
assign aao = ~AAO;  //complement 
assign aap = ~AAP;  //complement 
assign abo = ~ABO;  //complement 
assign abp = ~ABP;  //complement 
assign MAI =  LCA & pac  |  LCE & PAC  ; 
assign mai = ~MAI;  //complement 
assign MAJ =  LCB & pac  |  LCF & PAC  ; 
assign maj = ~MAJ;  //complement 
assign hbd = ~HBD;  //complement 
assign CBD =  BAK & BCK & tkh  |  BAL & BCL & TKH  ; 
assign cbd = ~CBD;  //complement 
assign dbd =  bak & bck & tkh  |  bal & bcl & TKH  ; 
assign DBD = ~dbd;  //complement 
assign oai = ~OAI;  //complement 
assign oaj = ~OAJ;  //complement 
assign GDF = ~gdf;  //complement 
assign GDG = ~gdg;  //complement 
assign GDH = ~gdh;  //complement 
assign CCA =  BAL & BCL & tks  |  BAM & BCM & TKS  ; 
assign cca = ~CCA;  //complement 
assign dca =  bal & bcl & tks  |  bam & bcm & TKS  ; 
assign DCA = ~dca;  //complement 
assign bal = ~BAL;  //complement 
assign bam = ~BAM;  //complement 
assign bcl = ~BCL;  //complement 
assign bcm = ~BCM;  //complement 
assign MBA =  LGA & pag  |  LGE & PAG  ; 
assign mba = ~MBA;  //complement 
assign MBB =  LGB & pag  |  LGF & PAG  ; 
assign mbb = ~MBB;  //complement 
assign hfd = ~HFD;  //complement 
assign CFD =  BBA & BDA & tkh  |  BBB & BDB & TKH  ; 
assign cfd = ~CFD;  //complement 
assign dfd =  bba & bda & tkh  |  bbb & bdb & TKH  ; 
assign DFD = ~dfd;  //complement 
assign oba = ~OBA;  //complement 
assign obb = ~OBB;  //complement 
assign GHG = ~ghg;  //complement 
assign GHH = ~ghh;  //complement 
assign CGA =  BBB & BDB & tkh  |  BBC & BDC & TKH  ; 
assign cga = ~CGA;  //complement 
assign bbb = ~BBB;  //complement 
assign bbc = ~BBC;  //complement 
assign bdb = ~BDB;  //complement 
assign bdc = ~BDC;  //complement 
assign MBQ =  LKA & pak  |  LKE & PAK  ; 
assign mbq = ~MBQ;  //complement 
assign MBR =  LKB & pak  |  LKF & PAK  ; 
assign mbr = ~MBR;  //complement 
assign hjd = ~HJD;  //complement 
assign CJD =  BBQ & BDQ & tkp  |  BBR & BDR & TKP  ; 
assign cjd = ~CJD;  //complement 
assign djd =  bbq & bdq & tkp  |  bbr & bdr & TKP  ; 
assign DJD = ~djd;  //complement 
assign obq = ~OBQ;  //complement 
assign obr = ~OBR;  //complement 
assign GLF = ~glf;  //complement 
assign GLG = ~glg;  //complement 
assign GLH = ~glh;  //complement 
assign CKA =  BBR & BDR & tkp  |  BBS & BDS & TKP  ; 
assign cka = ~CKA;  //complement 
assign dka =  bbr & bdr & tkp  |  bbs & bds & TKP  ; 
assign DKA = ~dka;  //complement 
assign bbr = ~BBR;  //complement 
assign bbs = ~BBS;  //complement 
assign bdr = ~BDR;  //complement 
assign bds = ~BDS;  //complement 
assign ocm = ~OCM;  //complement 
assign ocn = ~OCN;  //complement 
assign oco = ~OCO;  //complement 
assign ocp = ~OCP;  //complement 
assign GHF = ~ghf;  //complement 
assign dga =  bbb & bdb & tkw  |  bbc & bdc & TKW  ; 
assign DGA = ~dga;  //complement 
assign iab = ~IAB; //complement 
assign iac = ~IAC; //complement 
assign iad = ~IAD; //complement 
assign iae = ~IAE; //complement 
assign iaf = ~IAF; //complement 
assign iag = ~IAG; //complement 
assign iah = ~IAH; //complement 
assign iai = ~IAI; //complement 
assign iaj = ~IAJ; //complement 
assign iak = ~IAK; //complement 
assign ial = ~IAL; //complement 
assign iam = ~IAM; //complement 
assign ian = ~IAN; //complement 
assign iao = ~IAO; //complement 
assign iap = ~IAP; //complement 
assign iaq = ~IAQ; //complement 
assign iar = ~IAR; //complement 
assign ias = ~IAS; //complement 
assign iat = ~IAT; //complement 
assign iau = ~IAU; //complement 
assign iav = ~IAV; //complement 
assign iaw = ~IAW; //complement 
assign iax = ~IAX; //complement 
assign iay = ~IAY; //complement 
assign iaz = ~IAZ; //complement 
assign iba = ~IBA; //complement 
assign ibb = ~IBB; //complement 
assign ibc = ~IBC; //complement 
assign ibd = ~IBD; //complement 
assign ibe = ~IBE; //complement 
assign ibf = ~IBF; //complement 
assign ibg = ~IBG; //complement 
assign ibh = ~IBH; //complement 
assign ibi = ~IBI; //complement 
assign ibj = ~IBJ; //complement 
assign ibk = ~IBK; //complement 
assign ibl = ~IBL; //complement 
assign ibm = ~IBM; //complement 
assign ibn = ~IBN; //complement 
assign ibo = ~IBO; //complement 
assign ibp = ~IBP; //complement 
assign ibq = ~IBQ; //complement 
assign ibr = ~IBR; //complement 
assign ibs = ~IBS; //complement 
assign ibt = ~IBT; //complement 
assign ibu = ~IBU; //complement 
assign ibv = ~IBV; //complement 
assign ibw = ~IBW; //complement 
assign ibx = ~IBX; //complement 
assign iby = ~IBY; //complement 
assign ibz = ~IBZ; //complement 
assign icb = ~ICB; //complement 
assign icc = ~ICC; //complement 
assign icd = ~ICD; //complement 
assign ice = ~ICE; //complement 
assign icf = ~ICF; //complement 
assign icg = ~ICG; //complement 
assign ich = ~ICH; //complement 
assign ici = ~ICI; //complement 
assign ick = ~ICK; //complement 
assign icl = ~ICL; //complement 
assign icm = ~ICM; //complement 
assign icn = ~ICN; //complement 
assign ico = ~ICO; //complement 
assign icp = ~ICP; //complement 
assign icq = ~ICQ; //complement 
assign ics = ~ICS; //complement 
assign ict = ~ICT; //complement 
assign icu = ~ICU; //complement 
assign icv = ~ICV; //complement 
assign icw = ~ICW; //complement 
assign icx = ~ICX; //complement 
assign icy = ~ICY; //complement 
assign icz = ~ICZ; //complement 
assign ida = ~IDA; //complement 
assign idb = ~IDB; //complement 
assign idc = ~IDC; //complement 
assign idd = ~IDD; //complement 
assign ide = ~IDE; //complement 
assign idf = ~IDF; //complement 
assign idg = ~IDG; //complement 
assign idh = ~IDH; //complement 
assign idi = ~IDI; //complement 
assign idj = ~IDJ; //complement 
assign idk = ~IDK; //complement 
assign idl = ~IDL; //complement 
assign idm = ~IDM; //complement 
assign idn = ~IDN; //complement 
assign ido = ~IDO; //complement 
assign idp = ~IDP; //complement 
assign idq = ~IDQ; //complement 
assign idr = ~IDR; //complement 
assign ids = ~IDS; //complement 
assign idt = ~IDT; //complement 
assign idu = ~IDU; //complement 
assign idv = ~IDV; //complement 
assign idw = ~IDW; //complement 
assign idx = ~IDX; //complement 
assign idy = ~IDY; //complement 
assign idz = ~IDZ; //complement 
assign ief = ~IEF; //complement 
assign ieg = ~IEG; //complement 
assign ieh = ~IEH; //complement 
assign iei = ~IEI; //complement 
assign ieo = ~IEO; //complement 
assign iep = ~IEP; //complement 
assign ieq = ~IEQ; //complement 
assign ifff  = ~IFFF ; //complement 
assign ifo = ~IFO; //complement 
assign iga = ~IGA; //complement 
assign igb = ~IGB; //complement 
assign igc = ~IGC; //complement 
assign igd = ~IGD; //complement 
assign ige = ~IGE; //complement 
assign igf = ~IGF; //complement 
assign igg = ~IGG; //complement 
assign igh = ~IGH; //complement 
assign igi = ~IGI; //complement 
assign igj = ~IGJ; //complement 
assign igk = ~IGK; //complement 
assign igl = ~IGL; //complement 
assign igm = ~IGM; //complement 
assign ign = ~IGN; //complement 
assign igo = ~IGO; //complement 
assign igp = ~IGP; //complement 
assign iha = ~IHA; //complement 
assign ihb = ~IHB; //complement 
assign ihc = ~IHC; //complement 
assign ihd = ~IHD; //complement 
assign ihe = ~IHE; //complement 
assign ihf = ~IHF; //complement 
assign ihg = ~IHG; //complement 
assign ihh = ~IHH; //complement 
assign ihi = ~IHI; //complement 
assign ihj = ~IHJ; //complement 
assign ihk = ~IHK; //complement 
assign ihl = ~IHL; //complement 
assign ihm = ~IHM; //complement 
assign ihn = ~IHN; //complement 
assign iho = ~IHO; //complement 
assign ihp = ~IHP; //complement 
assign iua = ~IUA; //complement 
assign iub = ~IUB; //complement 
assign iva = ~IVA; //complement 
assign ivb = ~IVB; //complement 
assign ivc = ~IVC; //complement 
assign ivd = ~IVD; //complement 
assign ive = ~IVE; //complement 
assign ivf = ~IVF; //complement 
always@(posedge IZZ )
   begin 
 FEA <=  EBA & eaa  ; 
 AEA <=  ACA  |  QNI  |  QNH  ; 
 AEB <=  ACB  |  QNI  |  QNH  ; 
 ACA <=  AAA & TAA  |  ADA & TBA  |  ACA & TCA  ; 
 ACB <=  AAB & TAA  |  ADB & TBA  |  ACB & TCA  ; 
 QNF <=  QMI & qne  |  JEC  ; 
 AFA <=  ada & TFA  |  ADA & tfa  ; 
 AFB <=  adb & TFA  |  ADB & tfa  ; 
 ADA <=  IHA & TDA  |  BHA & TEA  ; 
 ADB <=  ABB & TDA  |  BHB & TEA  ; 
 FAD <=  EAA & EBB & EBC  |  EAB & EBC  |  EAC  ; 
 FAC <=  EBB & EAA  |  EAB  ; 
 qma <=  jba  |  jbb  |  jbc  ; 
 QNE <= QMH & QMD ; 
 QKA <=  QAA & QFA & qea  ; 
 QJB <= QJA ; 
 QJC <= QJB ; 
 QJE <= QJD ; 
 QJF <= QJE ; 
 AHA <=  AGB & TGA  |  AGA & tga  ; 
 AHB <=  AGC & TGA  |  AGB & tga  ; 
 AGA <=  FEA  ; 
 AGB <=  ECB  ; 
 QKB <=  QAA & QFA & QEA  ; 
 QJJ <=  QCB & QFB  |  QCB & QEB  |  QJJ & QGA  ; 
 PDB <= aha ; 
 qbb <= qba ; 
 FEB <=  EBB & eab  ; 
 QJD <=  QCA & qfa & qea  |  QAA  ; 
 AKA <=  aia  ; 
 AKB <=  aib & PDB  |  AIB & pdb  ; 
 FAB <= EAA ; 
 AIA <= AHA ; 
 AIB <= AHB ; 
 AJA <= AIA ; 
 AJB <= AIB ; 
 ALA <= AJA ; 
 ALB <= AJB ; 
 AMA <= AKA ; 
 AMB <= AKB ; 
 ANA <=  ALA & tha  |  QNO & THA  |  QNK & THA  ; 
 ANB <=  ALB & tha  |  QOC & THA  ; 
 AOA <=  AMA & thb  |  QNO & THB  ; 
 AOB <=  AMB & thb  |  QOC & THB  ; 
 BFA <= BEA ; 
 BFB <= BEB ; 
 BHA <= BGA ; 
 BHB <= BGG ; 
 bea <= iha ; 
 beb <= abb ; 
 BGA <= BFA ; 
 BGB <= BFB ; 
 TLA <= QNA ; 
 TLB <= QNA ; 
 TLC <= QNA ; 
 TLD <= QNA ; 
 qba <= ivb ; 
 qda <= ivd ; 
 QMB <= QMA ; 
 QMD <= QMC ; 
 QMC <= QMB ; 
 HAA <=  DAA & caa & tla  |  daa & TLA  |  CAA & TLA  ; 
 LDD <= tnb & KDD ; 
 LDH <= tnb & KDH ; 
 gch <=  dca & ccb & ccc  |  dcb & ccc  |  dcc  ; 
 qaa <= iva ; 
 qca <= ivc ; 
 qfa <= ivf ; 
 qea <= ive ; 
 QJA <=  IVC & ivf & ive  |  IVA  |  JGA  ; 
 ODC <=  IVC & ivf & ive  |  IVA  |  JGA  ; 
 ODA <=  IVC & ivf & ive  |  IVA  |  JGA  ; 
 ODB <=  IVC & ivf & ive  |  IVA  |  JGA  ; 
 HEA <=  DEA & cea & tla  |  dea & TLA  |  CEA & TLA  ; 
 LEA <= tnd & HEA ; 
 LEE <= tnd & hea ; 
 LHD <= tnd & KHD ; 
 LHH <= tnd & KHH ; 
 ggh <=  dga & cgb & cgc  |  dgb & cgc  |  dgc  ; 
 OEA <=  QCA & qfa & qea  |  QAA  ; 
 OEB <=  QCA & qfa & qea  |  QAA  ; 
 OEC <=  QCA & qfa & qea  |  QAA  ; 
 BBZ <= IBZ ; 
 PAM <=  KMA & KPA & KQA  |  KNA & KQA  |  KOA  ; 
 HIA <=  DIA & cia & tla  |  dia & TLA  |  CIA & TLA  ; 
 LIA <= tnf & HIA ; 
 LIE <= tnf & hia ; 
 LLD <= tnf & KLD ; 
 LLH <= tnf & KLH ; 
 gkh <=  dka & ckb & ckc  |  dkb & ckc  |  dkc  ; 
 LMA <= tnf & HMA ; 
 LME <= tnf & hma ; 
 HMA <=  DMA & cma & tla  |  dma & TLA  |  CMA & TLA  ; 
 AAA <= IGA ; 
 AAB <= IGB ; 
 ABB <= IHB ; 
 bac <=  iac & tib  |  icc & tib  |  iad & TIB  |  icd & TIB  ; 
 BCC <=  IAC & tia  |  ICC & tia  |  IAD & TIA  |  ICD & TIA  ; 
 gbf <=  dba & dba  ; 
 gbg <=  cbb & dba  |  dbb  ; 
 gbh <=  dba & cbb & cbc  |  dbb & cbc  |  dbc  ; 
 BAD <= IAD ; 
 BAE <= IAE ; 
 BCD <= ICD ; 
 BCE <= ICE ; 
 HDD <=  DDD & cdd & tlb  |  ddd & TLB  |  CDD & TLB  ; 
 OAA <=  LAA & TOC  |  LAB & toc  ; 
 OAB <=  LAB & TOC  |  LAC & toc  ; 
 gff <=  dfa & dfa  ; 
 gfg <=  cfb & dfa  |  dfb  ; 
 gfh <=  dfa & cfb & cfc  |  dfb & cfc  |  dfc  ; 
 BAT <= IAT ; 
 BAU <= IAU ; 
 BCT <= ICT ; 
 BCU <= ICU ; 
 HHD <=  DHD & chd & tlb  |  dhd & TLB  |  CHD & TLB  ; 
 OAQ <=  MAQ & TOE  |  MAR & toe  ; 
 OAR <=  MAR & TOE  |  MAS & toe  ; 
 gjf <=  dja & dja  ; 
 gjg <=  cjb & dja  |  djb  ; 
 gjh <=  dja & cjb & cjc  |  djb & cjc  |  djc  ; 
 BBJ <= IBJ ; 
 BBK <= IBK ; 
 BDJ <= IDJ ; 
 BDK <= IDK ; 
 HLD <=  DLD & cld & tlb  |  dld & TLB  |  CLD & TLA  ; 
 OBI <=  MBI & TOG  |  MBJ & tog  ; 
 OBJ <=  MBJ & TOG  |  MBK & tog  ; 
 gmf <= dma ; 
 GMB <= CMA ; 
 BDZ <=  IDZ & tib  ; 
 FEC <=  EBC & eac  ; 
 AEC <= ACC ; 
 AED <= ACD ; 
 ACC <=  AAC & TAA  |  ADC & TBA  |  ACC & TCA  ; 
 ACD <=  AAD & TAA  |  ADD & TBA  |  ACD & TCA  ; 
 FED <=  EBD & ead  ; 
 AFC <=  adc & TFA  |  ADC & tfa  ; 
 AFD <=  add & TFA  |  ADD & tfa  ; 
 ADC <=  ABC & TDA  |  BHC & TEA  ; 
 ADD <=  ABD & TDA  |  BHD & TEA  ; 
 FAE <=  EAA & EBB & EBC & EBD  |  EAB & EBC & EBD  |  EAC & EBD  |  EAD  ; 
 qdb <= qda ; 
 qbc <= qbb ; 
 qdc <= qdb ; 
 AHC <=  AGD & TGA  |  AGC & tga  ; 
 AHD <=  AGE & TGA  |  AGD & tga  ; 
 AGC <=  ECC  ; 
 AGD <=  ECD  ; 
 QKC <=  QCB & QFB & qeb  ; 
 OGA <=  QCB & QFB  |  QCB & QEB  |  QJJ & QGA  ; 
 OGB <=  QCB & QFB  |  QCB & QEB  |  QJJ & QGA  ; 
 OGC <=  QCB & QFB  |  QCB & QEB  |  QJJ & QGA  ; 
 PDC <= JDC ; 
 PDD <= JDD ; 
 QKD <=  QCB & QFB & QEB  ; 
 qab <= qaa ; 
 qeb <= qea ; 
 qfb <= qfa ; 
 qcb <= qca ; 
 AKC <=  aic & PDC  |  AIC & pdc  ; 
 AKD <=  aid & PDD  |  AID & pdd  ; 
 qac <= qab ; 
 qec <= qeb ; 
 qfc <= qfb ; 
 qcc <= qcb ; 
 AIC <= AHC ; 
 AID <= AHD ; 
 AJC <= AIC ; 
 AJD <= AID ; 
 ALC <= AJC ; 
 ALD <= AJD ; 
 AMC <= AKC ; 
 AMD <= AKD ; 
 ANC <=  ALC & tha  |  QOF & THA  ; 
 ANDD  <=  ALD & tha  ; 
 AOC <=  AMC & thb  |  QOF & THB  ; 
 AOD <=  AMD & thb  ; 
 BFC <= BEC ; 
 BFD <= BED ; 
 BHC <= BGC ; 
 BHD <= BGD ; 
 bec <= abc ; 
 bed <= abd ; 
 BGC <= BFC ; 
 BGD <= BFD ; 
 QPA <=  QPA & qba & qdc  |  QBA & qea  |  QDC & qec  ; 
 OMA <=  QPA & qba & qdc  |  QBA & qea  |  QDC & qec  ; 
 HAB <=  DAB & cab & tlc  |  dab & TLC  |  CAB & TLC  ; 
 LDC <= tnb & KDC ; 
 LDG <= tnb & KDG ; 
 LAA <= tnb & KAA ; 
 LAB <= tnb & KAB ; 
 gcf <=  dca & dca  ; 
 gcg <=  ccb & dca  |  dcb  ; 
 pai <=  kma & kna  |  kpa & kna  ; 
 HEB <=  DEB & ceb & tlc  |  deb & TLC  |  CEB & TLC  ; 
 LEB <= tnd & KEB ; 
 LEF <= tnd & KEF ; 
 LHC <= tnd & KHC ; 
 LHG <= tnd & KHG ; 
 ggf <=  dga & dga  ; 
 ggg <=  cgb & dga  |  dgb  ; 
 PAL <=  KMA & KPA & NEC  |  KNA & NEC  |  NCC  ; 
 HIB <=  DIB & cib & tlc  |  dib & TLC  |  CIB & TLC  ; 
 LIB <= tnf & KIB ; 
 LIF <= tnf & KIF ; 
 LLC <= tnf & KLC ; 
 LLG <= tnf & KLG ; 
 gkf <=  dka & dka  ; 
 gkg <=  ckb & dka  |  dkb  ; 
 AAC <= IGC ; 
 AAD <= IGD ; 
 ABC <= IHC ; 
 ABD <= IHD ; 
 bab <=  iab & tib  |  icb & tib  |  iac & TIB  |  icc & TIB  ; 
 BCB <=  IAB & tia  |  ICB & tia  |  IAC & TIA  |  ICC & TIA  ; 
 GBB <=  CBA & CBA  ; 
 GBC <=  DBB & CBA  |  CBB  ; 
 GBD <=  CBA & DBB & DBC  |  CBB & DBC  |  CBC  ; 
 OAO <=  MAO & TOB  |  MAP & tob  ; 
 OAP <=  MAP & TOB  |  MAQ & tob  ; 
 HDC <=  DDC & cdc & tld  |  ddc & TLD  |  CDC & TLD  ; 
 BAR <= IAR ; 
 BAS <= IAS ; 
 BCS <= ICS ; 
 GFB <=  CFA & CFA  ; 
 GFC <=  DFB & CFA  |  CFB  ; 
 GFD <=  CFA & DFB & DFC  |  CFB & DFC  |  CFC  ; 
 OBG <=  MBG & TOD  |  MBH & tod  ; 
 OBH <=  MBH & TOD  |  MBI & tod  ; 
 HHC <=  DHC & chc & tld  |  dhc & TLD  |  CHC & TLD  ; 
 BBH <= IBH ; 
 BBI <= IBI ; 
 BDH <= IDH ; 
 BDI <= IDI ; 
 GJB <=  CJA & CJA  ; 
 GJC <=  DJB & CJA  |  CJB  ; 
 GJD <=  CJA & DJB & DJC  |  CJB & DJC  |  CJC  ; 
 OBW <=  MBW & TOF  |  MBX & tof  ; 
 OBX <=  MBX & TOF  |  MBY & tof  ; 
 HLC <=  DLC & clc & tld  |  dlc & TLD  |  CLC & TLD  ; 
 BBX <= IBX ; 
 BBY <= IBY ; 
 BDX <= IDX ; 
 BDY <= IDY ; 
 OCA <=  AOA & TOL  |  ANA & tol  ; 
 OCB <=  AOB & TOL  |  ANB & tol  ; 
 OCC <=  AOC & TOL  |  ANC & tol  ; 
 OCD <=  AOD & TOL  |  ANDD  & tol  ; 
 QIA <=  QCA  |  QIA & IUA  ; 
 qga <= iua ; 
 FFA <=  EBE & eae  ; 
 AEE <= ACE ; 
 AEF <= ACF ; 
 ACE <=  AAE & TAA  |  ADE & TBA  |  ACE & TCA  ; 
 ACF <=  AAF & TAA  |  ADF & TBA  |  ACF & TCA  ; 
 FBE <=  EAE & EBF & EBG & EBH  |  EAF & EBG & EBH  |  EAG & EBH  |  EAH  ; 
 AFE <=  ade & TFA  |  ADE & tfa  ; 
 AFF <=  adf & TFA  |  ADF & tfa  ; 
 ADE <=  ABE & TDA  |  BHE & TEA  ; 
 ADF <=  ABF & TDA  |  BHF & TEA  ; 
 FBD <=  EAE & EBF & EBG  |  EAF & EBG  |  EAG  ; 
 FBC <=  EBF & EAE  |  EAF  ; 
 qbd <= qbc ; 
 qdd <= qdc ; 
 QRB <= QRA ; 
 QRE <= QRD ; 
 QRA <=  QQA  |  QQB  ; 
 QRC <= QRB ; 
 QRF <= QRE ; 
 QRH <= QRG ; 
 QRJ <= QRI ; 
 QJH <= QJG ; 
 QJI <= QJH ; 
 AHE <=  AGF & TGA  |  AGE & tga  ; 
 AHF <=  AGG & TGA  |  AGF & tga  ; 
 AGE <=  FFA & egb  |  ffa & EGB  ; 
 AGF <=  EDB & egb  |  EDE & EGB  ; 
 QRD <= QRC ; 
 QRG <= QRF ; 
 QRI <= QRH ; 
 QRK <= QRJ ; 
 QJG <=  QCB & qfb & qeb  |  QJG & QGA  ; 
 PDE <= JDE ; 
 PDF <= JDF ; 
 QQB <=  QBE & QHE  |  QQB & QGB  |  QDG & QHG  ; 
 QKE <=  QKE & QGB  |  QDG & QEG  |  QBE & QEE  ; 
 OKA <=  QKE & QGB  |  QDG & QEG  |  QBE & QEE  ; 
 AKE <=  aie & PDE  |  AIE & pde  ; 
 AKF <=  aif & PDF  |  AIF & pdf  ; 
 qad <= qac ; 
 qed <= qec ; 
 qfd <= qfc ; 
 QCD <= QCC ; 
 qhc <= qhb ; 
 qhe <= qhd ; 
 qhg <= qhf ; 
 AIE <= AHE ; 
 AIF <= AHF ; 
 AJE <= AIE ; 
 AJF <= AIF ; 
 ALE <= AJE ; 
 ALF <= AJF ; 
 AME <= AKE ; 
 AMF <= AKF ; 
 ANE <=  ALE & tha  ; 
 ANF <=  ALF & tha  ; 
 AOE <=  AME & thb  ; 
 AOF <=  AMF & thb  ; 
 BFE <= BEE ; 
 BFF <= BEF ; 
 BHE <= BGE ; 
 BHF <= BGF ; 
 FFB <=  EBF & eaf  ; 
 bee <= abe ; 
 bef <= abf ; 
 BGE <= BFE ; 
 BGF <= BFF ; 
 TLE <= QNA ; 
 TLF <= QNA ; 
 TLG <= QNA ; 
 TLH <= QNA ; 
 pae <=  kma  ; 
 pad <=  ZZI & gae & gbe & gce  |  hbe & gbe & gce  |  hce & gce  ; 
 GAA <=  CNA & CNA  ; 
 GAB <=  DAA & CNA  |  CAA  ; 
 FBB <= EAE ; 
 LDB <= tnb & KDB ; 
 LDF <= tnb & KDF ; 
 LAC <= tnb & KAC ; 
 LAD <= tnb & KAD ; 
 GCB <=  CCA & CCA  ; 
 GCC <=  DCB & CCA  |  CCB  ; 
 paf <=  gee & kma  |  hee & gee  ; 
 hee <=  dea  |  deb  |  dec  |  ded  ; 
 LEC <= tnd & KEC ; 
 LEG <= tnd & KEG ; 
 LHB <= tnd & KHB ; 
 LHF <= tnd & KHF ; 
 GGB <=  CGA & CGA  ; 
 GGC <=  DGB & CGA  |  CGB  ; 
 PAJ <=  KMA & KPA & HIE  |  KNA & HIE  |  GIE  ; 
 hie <=  dia  |  dib  |  dic  |  did  ; 
 qmo <=  qkw  |  qli  ; 
 LIC <= tnf & KIC ; 
 LIG <= tnf & KIG ; 
 LLB <= tnf & KLB ; 
 LLF <= tnf & KLF ; 
 GKB <=  CKA & CKA  ; 
 GKC <=  DKB & CKA  |  CKB  ; 
 qhb <= qha ; 
 qhd <= qhc ; 
 qhf <= qhe ; 
 QQA <=  QAB & QHB  |  QCC & QHC  |  QQA & QGB  ; 
 AAE <= IGE ; 
 AAF <= IGF ; 
 ABE <= IHE ; 
 ABF <= IHF ; 
 BAA <=  IAB & ICB & TIA  ; 
 OAC <=  LAC & TOA  |  LAD & toa  ; 
 OAD <=  LAD & TOA  |  MAE & toa  ; 
 HAC <=  DAC & cac & tle  |  dac & TLE  |  CAC & TLE  ; 
 GBE <=  CBA & DBB & DBC & DBD  |  CBB & DBC & DBD  |  CBC & DBD  |  CBD  ; 
 BAF <=  IAF & icf & ief  |  iaf & ICF & ief  |  iaf & icf & IEF  |  IAF & ICF & IEF  ;
 bcg <=  IAF & icf & ief  |  iaf & ICF & ief  |  iaf & icf & IEF  |  iaf & icf & ief  ;
 BCF <= IFFF  ; 
 HDB <=  DDB & cdb & tlf  |  ddb & TLF  |  CDB & TLF  ; 
 BAQ <=  IAQ & icq & ieq  |  iaq & ICQ & ieq  |  iaq & icq & IEQ  |  IAQ & ICQ & IEQ  ;
 bcr <=  IAQ & icq & ieq  |  iaq & ICQ & ieq  |  iaq & icq & IEQ  |  iaq & icq & ieq  ;
 HEC <=  DEC & cec & tle  |  dec & TLE  |  CEC & TLE  ; 
 GFE <=  CFA & DFB & DFC & DFD  |  CFB & DFC & DFD  |  CFC & DFD  |  CFD  ; 
 BAV <= IAV ; 
 BAW <= IAW ; 
 BCV <= ICV ; 
 BCW <= ICW ; 
 HHB <=  DHB & chb & tlf  |  dhb & TLF  |  CHB & TLF  ; 
 OAS <=  MAS & TOE  |  MAT & toe  ; 
 OAT <=  MAT & TOE  |  MAU & toe  ; 
 HIC <=  DIC & cic & tle  |  dic & TLE  |  CIC & TLE  ; 
 GJE <=  CJA & DJB & DJC & DJD  |  CJB & DJC & DJD  |  CJC & DJD  |  CJD  ; 
 BBL <= IBL ; 
 BBM <= IBM ; 
 BDL <= IDL ; 
 BDM <= IDM ; 
 HLB <=  DLB & clb & tlf  |  dlb & TLF  |  CLB & TLF  ; 
 OBK <=  MBK & TOG  |  MBL & tog  ; 
 OBL <=  MBL & TOG  |  MBM & tog  ; 
 FFD <=  EBH & eah  ; 
 QPC <=  QBC  |  QDE  |  QPC & IUA  ; 
 OMC <=  QBC  |  QDE  |  QPC & IUA  ; 
 qha <= iub ; 
 FFC <= eag & EBG ; 
 AEG <= ACG ; 
 AEH <= ACH ; 
 ACG <=  AAG & TAA  |  ADG & TBA  |  ACG & TCA  ; 
 ACH <=  AAH & TAA  |  ADH & TBA  |  ACH & TCA  ; 
 FFE <=  EBE & EBF & EBG & EBH  ; 
 AFG <=  adg & TFA  |  ADG & tfa  ; 
 AFH <=  adh & TFA  |  ADH & tfa  ; 
 ADG <=  ABG & TDA  |  BHG & TEA  ; 
 ADH <=  ABH & TDA  |  BHH & TEA  ; 
 fbh <=  ebe & eaf & eag  |  ebf & eag  |  ebg  ; 
 fbf <=  ebe & ebe  ; 
 fbg <=  eaf & ebe  |  ebf  ; 
 TBA <= QJF ; 
 TBB <= QJF ; 
 TCA <= QJI ; 
 TCB <= QJI ; 
 qbe <= qbd ; 
 qde <= qdd ; 
 qbf <= qbe ; 
 qdf <= qde ; 
 AHG <=  AGH & TGA  |  AGG & tga  ; 
 AHH <=  AGI & TGA  |  AGH & tga  ; 
 AGG <=  EDC & egb  |  EDF & EGB  ; 
 AGH <=  EDD & egb  |  EDG & EGB  ; 
 TGA <= QKL ; 
 TGB <= QKL ; 
 OFA <=  QCB & qfb & qeb  |  QJG & QGA  ; 
 OFB <=  QCB & qfb & qeb  |  QJG & QGA  ; 
 OFC <=  QCB & qfb & qeb  |  QJG & QGA  ; 
 pdg <=  jdg  ; 
 pdh <=  AHG  |  jdg  ; 
 QJS <=  QJS & QGB  |  JGB  ; 
 AKG <=  aig & PDG  |  AIG & pdg  ; 
 AKH <=  aih & PDH  |  AIH & pdh  ; 
 qaf <= qae ; 
 qef <= qee ; 
 qff <= qfe ; 
 qcf <= qce ; 
 qae <= qad ; 
 qee <= qed ; 
 qfe <= qfd ; 
 qce <= qcd ; 
 AIG <= AHG ; 
 AIH <= AHH ; 
 AJG <= AIG ; 
 AJH <= AIH ; 
 ALG <= AJG ; 
 ALH <= AJH ; 
 AMG <= AKG ; 
 AMH <= AKH ; 
 ANG <=  ALG & tha  ; 
 ANH <=  ALH & tha  ; 
 AOG <=  AMG & thb  ; 
 AOH <=  AMH & thb  ; 
 BFG <= BEG ; 
 BFH <= BEH ; 
 BHG <= BGG ; 
 BHH <= BGH ; 
 pah <=  nbc & kma  |  ndc & nbc  ; 
 beg <= abg ; 
 beh <= abh ; 
 BGG <= BFG ; 
 BGH <= BFH ; 
 pab <=  gae  ; 
 pac <=  gbe & gae  |  hbe & gbe  ; 
 GAC <=  CNA & DAA & DAB  |  CAA & DAB  |  CAB  ; 
 TAA <= QJL ; 
 TAB <= QJL ; 
 QJK <= QJJ ; 
 QJL <= QJK ; 
 LDA <= tnb & HDA ; 
 LDE <= tnb & hda ; 
 GCD <=  CCA & DCB & DCC  |  CCB & DCC  |  CCC  ; 
 pag <=  nbb & kma  |  ndb & nbb  ; 
 GEE <=  CEA & DEB & DEC & DED  |  CEB & DEC & DED  |  CEC & DED  |  CED  ; 
 LHA <= tnd & HHA ; 
 LHE <= tnd & hha ; 
 LED <= tnd & KED ; 
 LEH <= tnd & KEH ; 
 GGD <=  CGA & DGB & DGC  |  CGB & DGC  |  CGC  ; 
 PAK <=  KMA & KPA & NEB  |  KNA & NEB  |  NCB  ; 
 gib <=  cia  ; 
 GIC <=  CIB  |  CIA & DIB  ; 
 qnm <=  qnl  |  QMI  |  JEB  ; 
 LLA <= tnf & HLA ; 
 LLE <= tnf & hla ; 
 LID <= tnf & KID ; 
 LIH <= tnf & KIH ; 
 GKD <=  CKA & DKB & DKC  |  CKB & DKC  |  CKC  ; 
 AAG <= IGG ; 
 AAH <= IGH ; 
 ABG <= IHG ; 
 ABH <= IHH ; 
 TKQ <= QMM ; 
 TKR <= QMM ; 
 TKA <= QMM ; 
 TKB <= QMM ; 
 HAD <=  DAD & cad & tlg  |  dad & TLG  |  CAD & TLG  ; 
 HBE <=  DBA & DBB & DBC & DBD  ; 
 BAG <=  IAG & icg & ieg  |  iag & ICG & ieg  |  iag & icg & IEG  |  IAG & ICG & IEG  ;
 bch <=  IAG & icg & ieg  |  iag & ICG & ieg  |  iag & icg & IEG  |  iag & icg & ieg  ;
 HDA <=  DDA & cda & tlh  |  dda & TLH  |  CDA & TLH  ; 
 BAP <=  IAP & icp & iep  |  iap & ICP & iep  |  iap & icp & IEP  |  IAP & ICP & IEP  ;
 bcq <=  IAP & icp & iep  |  iap & ICP & iep  |  iap & icp & IEP  |  iap & icp & iep  ;
 HED <=  DED & ced & tlg  |  ded & TLG  |  CED & TLG  ; 
 hfe <=  dfa  |  dfb  |  dfc  |  dfd  ; 
 hff <=  dfa  |  dfb  |  dfc  |  dfd  ; 
 OAM <=  MAM & TOD  |  MAN & tod  ; 
 OAN <=  MAN & TOD  |  MAO & tod  ; 
 HHA <=  DHA & cha & tlh  |  dha & TLH  |  CHA & TLH  ; 
 BBF <= IBF ; 
 BBG <= IBG ; 
 BDF <= IDF ; 
 BDG <= IDG ; 
 HID <=  DID & cid & tlg  |  did & TLG  |  CID & TLG  ; 
 hje <=  dja  |  djb  |  djc  |  djd  ; 
 hjf <=  dja  |  djb  |  djc  |  djd  ; 
 OBE <=  MBE & TOF  |  MBF & tof  ; 
 OBF <=  MBF & TOF  |  MBG & tof  ; 
 HLA <=  DLA & cla & tlh  |  dla & TLH  |  CLA & TLH  ; 
 BBV <= IBV ; 
 BBW <= IBW ; 
 BDV <= IDV ; 
 BDW <= IDW ; 
 OCE <=  AOE & TOM  |  ANE & tom  ; 
 OCF <=  AOF & TOM  |  ANF & tom  ; 
 OCG <=  AOG & TOM  |  ANG & tom  ; 
 OCH <=  AOH & TOM  |  ANH & tom  ; 
 tki <= qmm ; 
 tkj <= qmm ; 
 tku <= qmm ; 
 tkv <= qmm ; 
 OBU <=  MBU & TOH  |  MBV & toh  ; 
 OBV <=  MBV & TOH  |  MBW & toh  ; 
 FGA <=  EBI & eai  ; 
 AEI <= ACI ; 
 AEJ <= ACJ ; 
 ACI <=  AAI & TAB  |  ADI & TBB  |  ACI & TCB  ; 
 ACJ <=  AAJ & TAB  |  ADJ & TBB  |  ACJ & TCB  ; 
 FCE <=  EAI & EBJ & EBK & EBL  |  EAJ & EBK & EBL  |  EAK & EBL  |  EAL  ; 
 AFI <=  adi & TFB  |  ADI & tfb  ; 
 AFJ <=  adj & TFB  |  ADJ & tfb  ; 
 ADI <=  ABI & TDB  |  BHI & TEB  ; 
 ADJ <=  ABJ & TDB  |  BHJ & TEB  ; 
 FCD <=  EAI & EBJ & EBK  |  EAJ & EBK  |  EAK  ; 
 FCB <=  EAI & EAI  ; 
 FCC <=  EBJ & EAI  |  EAJ  ; 
 TEA <= QJO ; 
 TEB <= QJO ; 
 TDA <= QJC ; 
 TDB <= QJC ; 
 TFA <= QKF ; 
 TFB <= QKF ; 
 QLC <= QLB ; 
 QLE <= QLD ; 
 QJN <= QJM ; 
 QJO <= QJN ; 
 QLD <= QLC ; 
 AHI <=  AGJ & TGB  |  AGI & tgb  ; 
 AHJ <=  AGK & TGB  |  AGJ & tgb  ; 
 AGI <=  FGA & egc  |  fga & EGC  ; 
 AGJ <=  EEB & egc  |  EEE & EGC  ; 
 qbg <= qbf ; 
 qdg <= qdf ; 
 qbh <= qbg ; 
 qdh <= qdg ; 
 QJM <=  QBD  |  QDF  |  QJM & QGA  ; 
 pdi <=  jdi  |  jdg  ; 
 pdj <=  jdj  |  jdg  ; 
 QLB <=  QAH & qfh  |  QCI & qfi  |  QLB & QGH  ; 
 OJD <=  QJS & QGB  |  JGB  ; 
 OJE <=  QJS & QGB  |  JGB  ; 
 OJF <=  QJS & QGB  |  JGB  ; 
 AKI <=  aii & PDI  |  AII & pdi  ; 
 AKJ <=  aij & PDJ  |  AIJ & pdj  ; 
 qah <= qag ; 
 qeh <= qeg ; 
 qfh <= qfg ; 
 qch <= qcg ; 
 qag <= qaf ; 
 qeg <= qef ; 
 qfg <= qff ; 
 qcg <= qcf ; 
 AII <= AHI ; 
 AIJ <= AHJ ; 
 AJI <= AII ; 
 AJJ <= AIJ ; 
 ALI <= AJI ; 
 ALJ <= AJJ ; 
 AMI <= AKI ; 
 AMJ <= AKJ ; 
 ANI <=  ALI & tha  ; 
 ANJ <=  ALJ & tha  ; 
 AOI <=  AMI & thb  ; 
 AOJ <=  AMJ & thb  ; 
 BFI <= BEI ; 
 BFJ <= BEJ ; 
 BHI <= BGI ; 
 BHJ <= BGJ ; 
 FGB <=  EBJ & eaj  ; 
 bei <= abi ; 
 bej <= abj ; 
 BGI <= BFI ; 
 BGJ <= BFJ ; 
 TLI <= QNA ; 
 TLJ <= QNA ; 
 TLK <= QNA ; 
 TLL <= QNA ; 
 QLF <=  QLB & QKO  |  QLB & QKR  ; 
 LBA <= tna & HBA ; 
 LBE <= tna & hba ; 
 LCD <= tna & KCD ; 
 LCH <= tna & KCH ; 
 GAD <=  CNA & DAA & DAB & DAC  |  CAA & DAB & DAC  |  CAB & DAC  |  CAC  ; 
 GCE <=  CCA & DCB & DCC & DCD  |  CCB & DCC & DCD  |  CCC & DCD  |  CCD  ; 
 OIA <= QJM ; 
 OIB <= QJM ; 
 OIC <= QJM ; 
 OID <= QJM ; 
 LFA <= tnc & HFA ; 
 LFE <= tnc & hfa ; 
 LGD <= tnc & KGD ; 
 LGH <= tnc & KGH ; 
 GED <=  CEA & DEB & DEC  |  CEB & DEC  |  CEC  ; 
 GGE <=  CGA & DGB & DGC & DGD  |  CGB & DGC & DGD  |  CGC & DGD  |  CGD  ; 
 QNH <=  qeh & QBH  |  qej & QDJ  |  QNH & QGE  ; 
 QNI <=  QEH & QBH  |  QEJ & QDJ  |  QNI & QGE  ; 
 LJA <= tne & HJA ; 
 LJE <= tne & hja ; 
 LKD <= tne & KKD ; 
 LKH <= tne & KKH ; 
 GID <=  CIA & DIB & DIC  |  CIB & DIC  |  CIC  ; 
 GKE <=  CKA & DKB & DKC & DKD  |  CKB & DKC & DKD  |  CKC & DKD  |  CKD  ; 
 qnl <=  qlf & qle  |  qlf & jed  ; 
 AAI <= IGI ; 
 AAJ <= IGJ ; 
 ABI <= IHI ; 
 ABJ <= IHJ ; 
 TKC <= QMM ; 
 TKD <= QMM ; 
 TKE <= QMM ; 
 TKF <= QMM ; 
 OAE <=  MAE & TOA  |  MAF & toa  ; 
 OAF <=  MAF & TOA  |  MAG & toa  ; 
 HBA <=  DBA & cba & tlj  |  dba & TLJ  |  CBA & TLJ  ; 
 BAH <=  IAH & ich & ieh  |  iah & ICH & ieh  |  iah & ich & IEH  |  IAH & ICH & IEH  ;
 bci <=  IAH & ich & ieh  |  iah & ICH & ieh  |  iah & ich & IEH  |  iah & ich & ieh  ;
 HCD <=  DCD & ccd & tli  |  dcd & TLI  |  CCD & TLI  ; 
 HDE <=  DDA & DDB & DDC & DDD  ; 
 BAO <=  IAO & ico & ieo  |  iao & ICO & ieo  |  iao & ico & IEO  |  IAO & ICO & IEO  ;
 bcp <=  IAO & ico & ieo  |  iao & ICO & ieo  |  iao & ico & IEO  |  iao & ico & ieo  ;
 HFA <=  DFA & cfa & tlj  |  dfa & TLJ  |  CFA & TLJ  ; 
 BAX <= IAX ; 
 BAY <= IAY ; 
 BCX <= ICX ; 
 BCY <= ICY ; 
 HGD <=  DGD & cgd & tli  |  dgd & TLI  |  CGD & TLI  ; 
 hhe <=  dha  |  dhb  |  dhc  |  dhd  ; 
 hhf <=  dha  |  dhb  |  dhc  |  dhd  ; 
 OAU <=  MAU & TOE  |  MAV & toe  ; 
 OAV <=  MAV & TOE  |  MAW & toe  ; 
 HJA <=  DJA & cja & tlj  |  dja & TLJ  |  CJA & TLJ  ; 
 BBN <= IBN ; 
 BBO <= IBO ; 
 BDN <= IDN ; 
 BDO <= IDO ; 
 HKD <=  DKD & ckd & tli  |  dkd & TLI  |  CKD & TLI  ; 
 hle <=  dla  |  dlb  |  dlc  |  dld  ; 
 hlf <=  dla  |  dlb  |  dlc  |  dld  ; 
 OBM <=  MBM & TOK  |  MBN & tok  ; 
 OBN <=  MBN & TOK  |  MBO & tok  ; 
 FGD <=  EBL & eal  ; 
 tkk <= qmm ; 
 tkl <= qmm ; 
 tkm <= qmm ; 
 tkn <= qmm ; 
 FGC <=  EBK & eak  ; 
 AEK <= ACK ; 
 AEL <= ACL ; 
 ACK <=  AAK & TAB  |  ADK & TBB  |  ACK & TCB  ; 
 ACL <=  AAL & TAB  |  ADL & TBB  |  ACL & TCB  ; 
 FGE <=  EBI & EBJ & EBK & EBL  ; 
 AFK <=  adk & TFB  |  ADK & tfb  ; 
 AFL <=  adl & TFB  |  ADL & tfb  ; 
 ADK <=  ABK & TDB  |  BHK & TEB  ; 
 ADL <=  ABL & TDB  |  BHL & TEB  ; 
 fch <=  ebi & eaj & eak  |  ebj & eak  |  ebk  ; 
 fcf <=  ebi & ebi  ; 
 fcg <=  eaj & ebi  |  ebi  ; 
 qbi <= qbh ; 
 qdi <= qdh ; 
 qbj <= qbi ; 
 qdj <= qdi ; 
 QKF <=  QBG  |  QDI  |  QKF & QGD  ; 
 qmk <=  qai  |  qfi  |  qei  ; 
 QNA <=  QNA & QGJ  |  QCJ & QFJ  |  QCK & QFK  |  QBM  |  QDO  ; 
 AHK <=  AGL & TGB  |  AGK & tgb  ; 
 AHL <=  AGM & TGB  |  AGL & tgb  ; 
 AGK <=  EEC & egc  |  EEF & EGC  ; 
 AGL <=  EED & egc  |  EEG & EGC  ; 
 qml <=  qcj  |  qfj  |  qej  ; 
 OHA <=  QBD  |  QDF  |  QJM & QGA  ; 
 OHB <=  QBD  |  QDF  |  QJM & QGA  ; 
 OHC <=  QBD  |  QDF  |  QJM & QGA  ; 
 pdk <=  jdk  |  jdg  ; 
 pdl <=  jdl  |  jdg  ; 
 QLA <=  QAJ & QFJ  |  QCK & QFK  |  QLA & QGJ  ; 
 QJR <=  QJR & QGB  |  JGE  ; 
 OJC <=  QJR & QGB  |  JGE  ; 
 AKK <=  aik & PDK  |  AIK & pdk  ; 
 AKL <=  ail & PDL  |  AIL & pdl  ; 
 qaj <= qai ; 
 qej <= qei ; 
 qfj <= qfi ; 
 qcj <= qci ; 
 qai <= qah ; 
 qei <= qeh ; 
 qfi <= qfh ; 
 qci <= qch ; 
 AIK <= AHK ; 
 AIL <= AHL ; 
 AJK <= AIK ; 
 AJL <= AIL ; 
 ALK <= AJK ; 
 ALL <= AJL ; 
 AMK <= AKK ; 
 AML <= AKL ; 
 ANK <=  ALK & tha  ; 
 ANL <=  ALL & tha  ; 
 AOK <=  AMK & thb  ; 
 AOL <=  AML & thb  ; 
 BFK <= BEK ; 
 BFL <= BEL ; 
 BHK <= BGK ; 
 BHL <= BGL ; 
 bek <= abk ; 
 bel <= abl ; 
 BGK <= BFK ; 
 BGL <= BFL ; 
 LBB <= tna & KBB ; 
 LBF <= tna & KBF ; 
 LCC <= tna & KCC ; 
 LCG <= tna & KCG ; 
 GAE <=  CNA & DAA & DAB & DAC & DAD  |  CAA & DAB & DAC & DAD  |  CAB & DAC & DAD  |  CAC & DAD & DAD  ; 
 hce <=  dca  |  dcb  |  dcc  |  dcd  ; 
 LFB <= tnc & KFB ; 
 LFF <= tnc & KFF ; 
 LGC <= tnc & KGC ; 
 LGG <= tnc & KGG ; 
 GEB <=  CEA & CEA  ; 
 GEC <=  DEB & CEA  |  CEB  ; 
 qmm <=  QMK  |  QML  |  QMM & QGJ  ; 
 TIA <=  QMK  |  QML  |  QMM & QGJ  ; 
 TIB <=  QMK  |  QML  |  QMM & QGJ  ; 
 hge <=  dga  |  dgb  |  dgc  |  dgd  ; 
 hgf <=  dga  |  dgb  |  dgc  |  dgd  ; 
 LJB <= tne & KJB ; 
 LJF <= tne & KJF ; 
 LKC <= tne & KKC ; 
 LKG <= tne & KKG ; 
 GIE <=  CIA & DIB & DIC & DID  |  CIB & DIC & DID  |  CIC & DID  |  CID  ; 
 hke <=  dka  |  dkb  |  dkc  |  dkd  ; 
 hkf <=  dka  |  dkb  |  dkc  |  dkd  ; 
 AAK <= IGK ; 
 AAL <= IGL ; 
 ABK <= IHK ; 
 ABL <= IHL ; 
 TKS <= QMM ; 
 TKT <= QMM ; 
 TKG <= QMM ; 
 TKH <= QMM ; 
 OAK <=  MAK & TOA  |  MAL & toa  ; 
 OAL <=  MAL & TOA  |  MAM & toa  ; 
 HBB <=  DBB & cbb & tll  |  dbb & TLL  |  CBB & TLL  ; 
 BAI <=  IAI & ici & iei  |  iai & ICI & iei  |  iai & ici & IEI  |  IAI & ICI & IEI  ;
 bcj <=  IAI & ici & iei  |  iai & ICI & iei  |  iai & ici & IEI  |  iai & ici & iei  ;
 HCC <=  DCC & ccc & tlk  |  dcc & TLK  |  CCC & TLK  ; 
 GDE <=  CDA & DDB & DDC & DDD  |  CDB & DDC & DDD  |  CDC & DDD  |  CDD  ; 
 BAN <= IAN ; 
 BCN <= ICN ; 
 BCO <= IFO ; 
 HFB <=  DFB & cfb & tll  |  dfb & TLL  |  CFB & TLL  ; 
 OBC <=  MBC & TOI  |  MBD & toi  ; 
 OBD <=  MBD & TOI  |  MBE & toi  ; 
 HGC <=  DGC & cgc & tlk  |  dgc & TLK  |  CGC & TLK  ; 
 GHE <=  CHA & DHB & DHC & DHD  |  CHB & DHC & DHD  |  CHC & DHD  |  CHD  ; 
 BBD <= IBD ; 
 BBE <= IBE ; 
 BDD <= IDD ; 
 BDE <= IDE ; 
 HJB <=  DJB & cjb & tll  |  djb & TLL  |  CJB & TLL  ; 
 OBS <=  MBS & TOJ  |  MBT & toj  ; 
 OBT <=  MBT & TOJ  |  MBU & toj  ; 
 HKC <=  DKC & ckc & tlk  |  dkc & TLK  |  CKC & TLK  ; 
 GLE <=  CLA & DLB & DLC & DLD  |  CLB & DLC & DLD  |  CLC & DLD  |  CLD  ; 
 BBT <= IBT ; 
 BBU <= IBU ; 
 BDT <= IDT ; 
 BDU <= IDU ; 
 OCI <=  AOI & TON  |  ANI & ton  ; 
 OCJ <=  AOJ & TON  |  ANJ & ton  ; 
 OCK <=  AOK & TON  |  ANK & ton  ; 
 OCL <=  AOL & TON  |  ANL & ton  ; 
 tko <= qmm ; 
 tkp <= qmm ; 
 tkw <= qmm ; 
 tkx <= qmm ; 
 FHB <=  EBN & ean  ; 
 FHA <=  EBM & eam  ; 
 AEM <= ACM ; 
 AEN <= ACN ; 
 QLQ <= QLP ; 
 QLU <= QLT ; 
 ACM <=  AAM & TAB  |  ADM & TBB  |  ACM & TCB  ; 
 ACN <=  AAN & TAB  |  ADN & TBB  |  ACN & TCB  ; 
 QMI <=  QLC & QMD  |  QMH & QLC  ; 
 QOH <=  QMH & QMD  ; 
 AFM <=  adm & TFB  |  ADM & tfb  ; 
 AFN <=  adn & TFB  |  ADN & tfb  ; 
 ADM <=  ABM & TDB  |  BHM & TEB  ; 
 ADN <=  ABN & TDB  |  BHN & TEB  ; 
 fdf <=  ebm & ebm  ; 
 fdg <=  ean & ebm  |  ebn  ; 
 FDB <=  EAM & EAM  ; 
 FDC <=  EBN & EAM  |  EAN  ; 
 QKN <= QKM ; 
 QKQ <= QKP ; 
 QOI <= QOH ; 
 qmn <= jeb ; 
 qbk <= qbj ; 
 qdk <= qdj ; 
 qbl <= qbk ; 
 qdl <= qdk ; 
 QKM <= JAA ; 
 QKP <= JAB ; 
 QKO <= QKN ; 
 QKR <= QKQ ; 
 AHM <=  AGN & TGB  |  AGM & tgb  ; 
 AHN <=  AGO & TGB  |  AGN & tgb  ; 
 AGM <=  FHA & egd  |  fha & EGD  ; 
 AGN <=  EFB & egd  |  EFE & EGD  ; 
 QKL <=  QKL & QGG  |  QBJ & QEJ  |  QDL & QEL  ; 
 QPB <=  QBD & qed  |  QDF & qef  |  QPB & QGA  ; 
 OMB <=  QBD & qed  |  QDF & qef  |  QPB & QGA  ; 
 PDM <=  JDM & JDG  ; 
 tna <=  qnf & qle  |  qnf & qmn  ; 
 tnb <=  qnf & qle  |  qnf & qmn  ; 
 tnc <=  qnf & qle  |  qnf & qmn  ; 
 QJQ <=  QJQ & QGB  |  JGD  ; 
 OJB <=  QJQ & QGB  |  JGD  ; 
 AKM <=  aim & PDM  |  AIM & pdm  ; 
 AKN <=  ain & PDN  |  AIN & pdn  ; 
 qck <= qcj ; 
 qek <= qej ; 
 qfk <= qfj ; 
 qel <= qek ; 
 AIM <= AHM ; 
 AIN <= AHN ; 
 AJM <= AIM ; 
 AJN <= AIN ; 
 ALM <= AJM ; 
 ALN <= AJN ; 
 AMN <= AKN ; 
 AMM <= AKM ; 
 ANM <=  ALM & tha  ; 
 ANN <=  ALN & tha  |  QOG & THA  ; 
 AOM <=  AMM & thb  ; 
 AON <=  AMN & thb  |  QOG & THB  ; 
 BFM <= BEM ; 
 BFN <= BEN ; 
 BHM <= BGM ; 
 BHN <= BGN ; 
 QLV <= QLU ; 
 QLR <= QLQ ; 
 bem <= abm ; 
 ben <= abn ; 
 BGM <= BFM ; 
 BGN <= BFN ; 
 TLM <= QNA ; 
 TLN <= QNA ; 
 TLO <= QNA ; 
 TLP <= QNA ; 
 LBC <= tna & KBC ; 
 LBG <= tna & KBG ; 
 LCB <= tna & KCB ; 
 LCF <= tna & KCF ; 
 PBA <=  KMB & KPB & KQB & HMA & QOJ  |  KNB & KQB & HMA & QOJ  |  KOB & HMA & QOJ  ; 
 HCB <=  DCB & ccb & tlm  |  dcb & TLM  |  CCB & TLM  ; 
 LFC <= tnc & KFC ; 
 LFG <= tnc & KFG ; 
 LGB <= tnc & KGB ; 
 LGF <= tnc & KGF ; 
 gef <=  dea & dea  ; 
 geg <=  ceb & dea  |  deb  ; 
 HGB <=  DGB & cgb & tlm  |  dgb & TLM  |  CGB & TLM  ; 
 LJC <= tne & KJC ; 
 LJG <= tne & KJG ; 
 LKB <= tne & KKB ; 
 LKF <= tne & KKF ; 
 gif <=  dia & dia  ; 
 gig <=  cib & dia  |  dib  ; 
 HKB <=  DKB & ckb & tlm  |  dkb & TLM  |  CKB & TLM  ; 
 AAM <= IGM ; 
 AAN <= IGN ; 
 ABM <= IHM ; 
 ABN <= IHN ; 
 HBC <=  DBC & cbc & tln  |  dbc & TLN  |  CBC & TLN  ; 
 BAJ <= IAJ ; 
 BAK <= IAK ; 
 BCK <= ICK ; 
 GDB <=  CDA & CDA  ; 
 GDC <=  DDB & CDA  |  CDB  ; 
 GDD <=  CDA & DDB & DDC  |  CDB & DDC  |  CDC  ; 
 OAG <=  MAG & TOC  |  MAH & toc  ; 
 OAH <=  MAH & TOC  |  MAI & toc  ; 
 HFC <=  DFC & cfc & tln  |  dfc & TLN  |  CFC & TLN  ; 
 BAZ <= IAZ ; 
 BBA <= IBA ; 
 BCZ <= ICZ ; 
 BDA <= IDA ; 
 GHC <=  DHB & CHA  |  CHB  ; 
 GHD <=  CHA & DHB & DHC  |  CHB & DHC  |  CHC  ; 
 OAW <=  MAW & TOE  |  MAX & toe  ; 
 OAX <=  MAX & TOE  |  MBA & toe  ; 
 HJC <=  DJC & cjc & tln  |  djc & TLN  |  CJC & TLM  ; 
 BBP <= IBP ; 
 BBQ <= IBQ ; 
 BDP <= IDP ; 
 BDQ <= IDQ ; 
 GLB <=  CLA & CLA  ; 
 GLC <=  DLB & CLA  |  CLB  ; 
 GLD <=  CLA & DLB & DLC  |  CLB & DLC  |  CLC  ; 
 OBO <=  MBO & TOK  |  MBP & tok  ; 
 OBP <=  MBP & TOK  |  MBQ & tok  ; 
 QLP <= QLO ; 
 GHB <= CHA ; 
 AFP <= ADP ; 
 FHC <=  EBO & eao  ; 
 OLA <=  QOL & QRK  ; 
 FIA <=  AEP & afp  |  aep & AFP  ; 
 AEO <= ACO ; 
 AEP <= ACP ; 
 QLO <= EAO ; 
 QLS <= ebo ; 
 ACO <=  aao & TAB  |  ADO & TBB  |  ACO & TCB  ; 
 ACP <=  AAP & TAB  |  ADP & TBB  |  ACP & TCB  ; 
 QMF <= QME ; 
 QMH <= QMG ; 
 QOA <= QLK ; 
 QOE <= QOD ; 
 QKT <= QKS ; 
 QKV <= QKU ; 
 QKX <= QKW ; 
 QLH <= QLG ; 
 AFO <=  ado & TFB  |  ADO & tfb  ; 
 ADO <=  abo & TDB  |  bho & TEB  ; 
 ADP <=  ABP & TDB  |  BHP & TEB  ; 
 QMG <= QMF ; 
 QOD <= QLM ; 
 QOB <= QOA ; 
 QOF <= QOE ; 
 QKU <= QKT ; 
 QKW <= QKV ; 
 QKY <= QKX ; 
 QLI <= QLH ; 
 qks <=  jcb  |  jcc  |  jcd  ; 
 qme <=  jca  |  jcb  |  jcc  |  jcd  ; 
 QLK <=  QLG & QKR  ; 
 QLM <=  QLL & QKR  |  QLL & AGP  |  QLL & QKU  ; 
 qgd <= qgc ; 
 qgf <= qge ; 
 qgh <= qgg ; 
 qgj <= qgi ; 
 qgc <= qgb ; 
 qge <= qgd ; 
 qgg <= qgf ; 
 qgi <= qgh ; 
 AHO <=  AGO  ; 
 AHP <=  AGP  ; 
 AGO <=  EFC & egd  |  EFF & EGD  ; 
 QLG <=  qek & QBK  |  qem & QDM  |  QLG & QGH  ; 
 QLL <=  QEK & QBK  |  QEM & QDM  |  QLL & QGH  ; 
 QPD <=  QBD & QED  |  QDF & QEF  |  QPD & QGA  ; 
 OMD <=  QBD & QED  |  QDF & QEF  |  QPD & QGA  ; 
 PDO <=  JDO & JDM & JDG  ; 
 PDN <=  ahm & JDM & JDG  ; 
 tnd <=  qnf & qle  |  qnf & qmn  ; 
 tne <=  qnf & qle  |  qnf & qmn  ; 
 tnf <=  qnf & qle  |  qnf & qmn  ; 
 QJP <=  QJP & QGB & jgb  |  jgb & qgc  ; 
 OJA <=  QJP & QGB & jgb  |  jgb & qgc  ; 
 AKO <=  AIO & PDO  |  aio & pdo  ; 
 JEA <=  AIN & aio  ; 
 qem <= qel ; 
 qbm <= qbl ; 
 qdm <= qdl ; 
 qdo <= qdn ; 
 qdn <= qdm ; 
 qgb <= qga ; 
 QLJ <= QLI ; 
 AIO <= AHO ; 
 AIP <= AHP ; 
 AJO <= aio ; 
 AJP <= AIP ; 
 ALO <= AJO ; 
 ALP <= AJP ; 
 AMO <= AKO ; 
 AMP <= AKP ; 
 ANP <=  ALP & tha  |  ALP & QNK  ; 
 AOO <=  AMO & thb  |  QOG & THB  |  THB & QNK  ; 
 BFO <= BEO ; 
 BFP <= BEP ; 
 BHO <= BGO ; 
 BHP <= BGP ; 
 ANO <=  ALO & tha  |  QOG & THA  |  THA & QNK  ; 
 beo <= abo ; 
 bep <= abp ; 
 BGO <= BFO ; 
 BGP <= BFP ; 
 AOP <=  AMP & thb  |  AMP & QNK  ; 
 AKP <=  AIP  ; 
 LCA <= tna & HCA ; 
 LCE <= tna & hca ; 
 LBD <= tna & KBD ; 
 LBH <= tna & KBH ; 
 QLN <=  QLF  |  QLK  |  QLM  ; 
 QLT <=  QLS  ; 
 QNO <= qnf & QNM ; 
 pca <=  KMB & KPB & KQB  |  KNB & KQB  |  KOB  |  HMA  |  qoj  ; 
 HCA <=  DCA & cca & tlo  |  dca & TLO  |  CCA & TLO  ; 
 QOJ <=  qoi  |  qle  ; 
 LGA <= tnc & HGA ; 
 LGE <= tnc & hga ; 
 LFD <= tnc & KFD ; 
 LFH <= tnc & KFH ; 
 geh <=  dea & ceb & cec  |  deb & cec  |  dec  ; 
 qoc <=  qob & qlj  |  qob & jee  ; 
 QOL <=  QNO  |  QOC  |  QOF & qky  ; 
 HGA <=  DGA & cga & tlo  |  dga & TLO  |  CGA & TLO  ; 
 LKA <= tne & HKA ; 
 LKE <= tne & hka ; 
 LJD <= tne & KJD ; 
 LJH <= tne & KJH ; 
 gih <=  dia & cib & cic  |  dib & cic  |  dic  ; 
 QMJ <=  QMI  |  QLN  |  QLA  ; 
 JED <= ago & AGN ; 
 QNJ <= QLA ; 
 QNK <= QNJ ; 
 HKA <=  DKA & cka & tlo  |  dka & TLO  |  CKA & TLO  ; 
 QOG <=  QLJ & JEE  |  QNM & qnf  |  QOB  |  QOE  ; 
 AGP <=  FIA  ; 
 THA <=  QMJ  |  JEA & QLE  |  JEE & QLJ  |  QMN & QLE  |  QNF  ; 
 THB <=  QMJ  |  JEA & QLE  |  JEE & QLJ  |  QMN & QLE  |  QNF  ; 
 AAO <= IGO ; 
 AAP <= IGP ; 
 ABO <= IHO ; 
 ABP <= IHP ; 
 HBD <=  DBD & cbd & tle  |  dbd & TLP  |  CBD & TLP  ; 
 OAI <=  MAI & TOB  |  MAJ & tob  ; 
 OAJ <=  MAJ & TOB  |  MAK & tob  ; 
 gdf <=  dda & dda  ; 
 gdg <=  cdb & dda  |  ddb  ; 
 gdh <=  dda & cdb & cdc  |  ddb & cdc  |  ddc  ; 
 BAL <= IAL ; 
 BAM <= IAM ; 
 BCL <= ICL ; 
 BCM <= ICM ; 
 HFD <=  DFD & cfd & tlp  |  dfd & TLP  |  CFD & TLP  ; 
 OBA <=  MBA & TOI  |  MBB & toi  ; 
 OBB <=  MBB & TOI  |  MBC & toi  ; 
 ghg <=  chb & dha  |  dhb  ; 
 ghh <=  dha & chb & chc  |  dhb & chc  |  dhc  ; 
 BBB <= IBB ; 
 BBC <= IBC ; 
 BDB <= IDB ; 
 BDC <= IDC ; 
 HJD <=  DJD & cjd & tlp  |  djd & TLP  |  CJD & TLP  ; 
 OBQ <=  MBQ & TOJ  |  MBR & toj  ; 
 OBR <=  MBR & TOJ  |  MBS & toj  ; 
 glf <=  dla & dla  ; 
 glg <=  clb & dla  |  dlb  ; 
 glh <=  dla & clb & clc  |  dlb & clc  |  dlc  ; 
 BBR <= IBR ; 
 BBS <= IBS ; 
 BDR <= IDR ; 
 BDS <= IDS ; 
 OCM <=  AOM & TOO  |  ANM & too  ; 
 OCN <=  AON & TOO  |  ANN & too  ; 
 OCO <=  AOO & TOO  |  ANO & too  ; 
 OCP <=  AOP & TOO  |  ANP & too  ; 
 ghf <=  dha  ; 
end 
endmodule;
