module jb( IZZ,
 IAA, 
 IAB, 
 IAC, 
 IAD, 
 IAE, 
 IAF, 
 IAG, 
 IAH, 
 IAI, 
 IAJ, 
 IAK, 
 IAL, 
 IAM, 
 IAN, 
 IAO, 
 IAP, 
 IBA, 
 IBB, 
 IBC, 
 IBD, 
 IBE, 
 IBF, 
 IBG, 
 IBH, 
 IBI, 
 IBJ, 
 IBK, 
 IBL, 
 IBM, 
 IBN, 
 IBO, 
 IBP, 
 ICA, 
 ICB, 
 ICC, 
 ICD, 
 ICE, 
 ICF, 
 ICG, 
 ICH, 
 ICI, 
 ICJ, 
 ICK, 
 ICL, 
 ICM, 
 ICN, 
 ICO, 
 ICP, 
 IDA, 
 IDB, 
 IDC, 
 IDD, 
 IDE, 
 IDF, 
 IEA, 
 IEB, 
 IFA, 
 IGA, 
 IHA, 
 IHB, 
 IHF, 
 IJA, 
 IKA, 
 IKB, 
 IKC, 
 IKD, 
 IKE, 
 IKF, 
 IKG, 
 IKH, 
 ILA, 
 OAA, 
 OAB, 
 OAC, 
 OAD, 
 OAE, 
 OAF, 
 OAG, 
 OAH, 
 OAI, 
 OAJ, 
 OAK, 
 OAL, 
 OAM, 
 OAN, 
 OAO, 
 OAP, 
 OBA, 
 OBB, 
 OBC, 
 OBD, 
 OBE, 
 OBF, 
 OBG, 
 OBH, 
 OBI, 
 OBJ, 
 OBK, 
 OBL, 
 OBM, 
 OBN, 
 OBO, 
 OBP, 
 OCA, 
 OCB, 
 OCC, 
 OCD, 
 OCE, 
 OCF, 
 OCG, 
 OCH, 
 OCI, 
 OCJ, 
 OCK, 
 OCL, 
 OCM, 
 OCN, 
 OCO, 
 OCP, 
 ODA, 
 ODB, 
 ODC, 
 ODD, 
 ODE, 
 ODF, 
 ODG, 
 ODH, 
 ODI, 
 ODJ, 
 ODK, 
 ODL, 
 ODM, 
 ODN, 
 ODO, 
 ODP, 
 OEA, 
 OEB, 
 OEC, 
 OED, 
 OEE, 
 OEF, 
 OEG, 
 OEH, 
 OEI, 
 OEJ, 
 OEK, 
 OEL, 
 OEM, 
 OEN, 
 OEO, 
 OEP, 
 OFA, 
 OFB, 
 OFC, 
 OFD, 
 OFE, 
 OFF, 
 OFG, 
 OFH, 
 OFI, 
 OFJ, 
 OFK, 
 OFL, 
 OFM, 
 OFN, 
 OFO, 
 OFP, 
 OGA, 
 OGB, 
 OGC, 
 OGD, 
 OGE, 
 OGF, 
 OGG, 
 OGH, 
 OGI, 
 OGJ, 
 OGK, 
 OGL, 
 OGM, 
 OGN, 
 OGO, 
 OGP, 
 OHA, 
 OHB, 
 OHC, 
 OHD, 
 OHE, 
 OHF, 
 OHG, 
 OHH, 
 OHI, 
 OHJ, 
 OHK, 
 OHL, 
 OHM, 
 OHN, 
 OHO, 
 OHP, 
 OIA, 
 OIB, 
 OIC, 
 OID, 
 OIE, 
 OIF, 
 OIG, 
 OIH, 
 OJA, 
 OJB, 
 OJC, 
 OJD, 
 OJE, 
 OJF, 
 OJG, 
 OJH, 
 OJI, 
 OJJ, 
 OJK, 
 OJL, 
 OKA, 
 OKB, 
 OKC, 
 OKD, 
 OKE, 
 OKF, 
 OLA, 
 OLB, 
 OLC, 
 OLD, 
 OLF, 
 OMA, 
 OMB, 
 OMC, 
 OMD, 
 OMF, 
 ONA, 
 ONB, 
 ONC, 
 OND, 
 ONE, 
 ONF, 
 ORA, 
 ORB, 
 ORC, 
 ORD, 
 OSA, 
 OSB, 
 OSC, 
 OSD, 
 OSE, 
 OSF, 
 OSG, 
 OSH, 
 OTA, 
 OUA, 
 OUB, 
OUC ); 
    
 input IZZ; 
 input IAA; 
 input IAB; 
 input IAC; 
 input IAD; 
 input IAE; 
 input IAF; 
 input IAG; 
 input IAH; 
 input IAI; 
 input IAJ; 
 input IAK; 
 input IAL; 
 input IAM; 
 input IAN; 
 input IAO; 
 input IAP; 
 input IBA; 
 input IBB; 
 input IBC; 
 input IBD; 
 input IBE; 
 input IBF; 
 input IBG; 
 input IBH; 
 input IBI; 
 input IBJ; 
 input IBK; 
 input IBL; 
 input IBM; 
 input IBN; 
 input IBO; 
 input IBP; 
 input ICA; 
 input ICB; 
 input ICC; 
 input ICD; 
 input ICE; 
 input ICF; 
 input ICG; 
 input ICH; 
 input ICI; 
 input ICJ; 
 input ICK; 
 input ICL; 
 input ICM; 
 input ICN; 
 input ICO; 
 input ICP; 
 input IDA; 
 input IDB; 
 input IDC; 
 input IDD; 
 input IDE; 
 input IDF; 
 input IEA; 
 input IEB; 
 input IFA; 
 input IGA; 
 input IHA; 
 input IHB; 
 input IHF; 
 input IJA; 
 input IKA; 
 input IKB; 
 input IKC; 
 input IKD; 
 input IKE; 
 input IKF; 
 input IKG; 
 input IKH; 
 input ILA; 
 output OAA; 
 output OAB; 
 output OAC; 
 output OAD; 
 output OAE; 
 output OAF; 
 output OAG; 
 output OAH; 
 output OAI; 
 output OAJ; 
 output OAK; 
 output OAL; 
 output OAM; 
 output OAN; 
 output OAO; 
 output OAP; 
 output OBA; 
 output OBB; 
 output OBC; 
 output OBD; 
 output OBE; 
 output OBF; 
 output OBG; 
 output OBH; 
 output OBI; 
 output OBJ; 
 output OBK; 
 output OBL; 
 output OBM; 
 output OBN; 
 output OBO; 
 output OBP; 
 output OCA; 
 output OCB; 
 output OCC; 
 output OCD; 
 output OCE; 
 output OCF; 
 output OCG; 
 output OCH; 
 output OCI; 
 output OCJ; 
 output OCK; 
 output OCL; 
 output OCM; 
 output OCN; 
 output OCO; 
 output OCP; 
 output ODA; 
 output ODB; 
 output ODC; 
 output ODD; 
 output ODE; 
 output ODF; 
 output ODG; 
 output ODH; 
 output ODI; 
 output ODJ; 
 output ODK; 
 output ODL; 
 output ODM; 
 output ODN; 
 output ODO; 
 output ODP; 
 output OEA; 
 output OEB; 
 output OEC; 
 output OED; 
 output OEE; 
 output OEF; 
 output OEG; 
 output OEH; 
 output OEI; 
 output OEJ; 
 output OEK; 
 output OEL; 
 output OEM; 
 output OEN; 
 output OEO; 
 output OEP; 
 output OFA; 
 output OFB; 
 output OFC; 
 output OFD; 
 output OFE; 
 output OFF; 
 output OFG; 
 output OFH; 
 output OFI; 
 output OFJ; 
 output OFK; 
 output OFL; 
 output OFM; 
 output OFN; 
 output OFO; 
 output OFP; 
 output OGA; 
 output OGB; 
 output OGC; 
 output OGD; 
 output OGE; 
 output OGF; 
 output OGG; 
 output OGH; 
 output OGI; 
 output OGJ; 
 output OGK; 
 output OGL; 
 output OGM; 
 output OGN; 
 output OGO; 
 output OGP; 
 output OHA; 
 output OHB; 
 output OHC; 
 output OHD; 
 output OHE; 
 output OHF; 
 output OHG; 
 output OHH; 
 output OHI; 
 output OHJ; 
 output OHK; 
 output OHL; 
 output OHM; 
 output OHN; 
 output OHO; 
 output OHP; 
 output OIA; 
 output OIB; 
 output OIC; 
 output OID; 
 output OIE; 
 output OIF; 
 output OIG; 
 output OIH; 
 output OJA; 
 output OJB; 
 output OJC; 
 output OJD; 
 output OJE; 
 output OJF; 
 output OJG; 
 output OJH; 
 output OJI; 
 output OJJ; 
 output OJK; 
 output OJL; 
 output OKA; 
 output OKB; 
 output OKC; 
 output OKD; 
 output OKE; 
 output OKF; 
 output OLA; 
 output OLB; 
 output OLC; 
 output OLD; 
 output OLF; 
 output OMA; 
 output OMB; 
 output OMC; 
 output OMD; 
 output OMF; 
 output ONA; 
 output ONB; 
 output ONC; 
 output OND; 
 output ONE; 
 output ONF; 
 output ORA; 
 output ORB; 
 output ORC; 
 output ORD; 
 output OSA; 
 output OSB; 
 output OSC; 
 output OSD; 
 output OSE; 
 output OSF; 
 output OSG; 
 output OSH; 
 output OTA; 
 output OUA; 
 output OUB; 
 output OUC; 
  
  
reg  AAA ;
reg  AAB ;
reg  AAC ;
reg  AAD ;
reg  AAE ;
reg  AAF ;
reg  AAG ;
reg  AAH ;
reg  AAI ;
reg  AAJ ;
reg  AAK ;
reg  AAL ;
reg  AAM ;
reg  AAN ;
reg  AAO ;
reg  AAP ;
reg  ABA ;
reg  ABB ;
reg  ABC ;
reg  ABD ;
reg  ABE ;
reg  ABF ;
reg  ABG ;
reg  ABH ;
reg  ABI ;
reg  ABJ ;
reg  ABK ;
reg  ABL ;
reg  ABM ;
reg  ABN ;
reg  ABO ;
reg  ABP ;
reg  BAA ;
reg  BAB ;
reg  BAC ;
reg  BAD ;
reg  BAE ;
reg  BAF ;
reg  bai ;
reg  baj ;
reg  bak ;
reg  bal ;
reg  bam ;
reg  ban ;
reg  bba ;
reg  bbb ;
reg  bbc ;
reg  bbd ;
reg  bbe ;
reg  bbf ;
reg  bbg ;
reg  bbi ;
reg  bbj ;
reg  bbk ;
reg  bbl ;
reg  bbm ;
reg  bbn ;
reg  bbo ;
reg  bca ;
reg  bcb ;
reg  bcc ;
reg  bcd ;
reg  bce ;
reg  bcf ;
reg  bcg ;
reg  bda ;
reg  bdb ;
reg  bdc ;
reg  bdd ;
reg  bde ;
reg  bdf ;
reg  bdg ;
reg  bdi ;
reg  bdj ;
reg  bdk ;
reg  bdl ;
reg  bdm ;
reg  bdn ;
reg  bdo ;
reg  bdp ;
reg  bea ;
reg  beb ;
reg  bec ;
reg  bed ;
reg  bee ;
reg  bef ;
reg  beg ;
reg  beh ;
reg  CAA ;
reg  CAB ;
reg  CAC ;
reg  CAD ;
reg  CAE ;
reg  CAF ;
reg  CBA ;
reg  CBB ;
reg  CBC ;
reg  CBD ;
reg  CBE ;
reg  CBF ;
reg  CCA ;
reg  CCB ;
reg  CCC ;
reg  CCD ;
reg  CCE ;
reg  CCF ;
reg  CDA ;
reg  CDB ;
reg  CDC ;
reg  CDD ;
reg  CDE ;
reg  CDF ;
reg  CEA ;
reg  CEB ;
reg  CEC ;
reg  CED ;
reg  CEE ;
reg  CEF ;
reg  CFA ;
reg  CFB ;
reg  CFC ;
reg  CFD ;
reg  CFE ;
reg  CFF ;
reg  eaa ;
reg  eab ;
reg  eac ;
reg  ead ;
reg  eae ;
reg  eaf ;
reg  eag ;
reg  eah ;
reg  eai ;
reg  eaj ;
reg  eak ;
reg  eal ;
reg  eam ;
reg  ean ;
reg  eao ;
reg  eap ;
reg  ebj ;
reg  ebk ;
reg  ebl ;
reg  ebm ;
reg  ebn ;
reg  ebo ;
reg  ebp ;
reg  ecm ;
reg  ecn ;
reg  eco ;
reg  ecp ;
reg  GAA ;
reg  GAB ;
reg  GAC ;
reg  GAD ;
reg  GAE ;
reg  GAF ;
reg  GAG ;
reg  GAH ;
reg  GAI ;
reg  GAJ ;
reg  GAK ;
reg  gba ;
reg  gbb ;
reg  gbc ;
reg  gbd ;
reg  gbe ;
reg  gbf ;
reg  gbg ;
reg  gbh ;
reg  gbk ;
reg  gbl ;
reg  gbn ;
reg  gbo ;
reg  gca ;
reg  gcb ;
reg  gcc ;
reg  gcd ;
reg  gce ;
reg  gcf ;
reg  gch ;
reg  gci ;
reg  gcj ;
reg  gck ;
reg  gcl ;
reg  gcm ;
reg  gcn ;
reg  gco ;
reg  gcp ;
reg  gda ;
reg  gdb ;
reg  gdc ;
reg  LAA ;
reg  LAB ;
reg  LAC ;
reg  LAD ;
reg  LAE ;
reg  LAF ;
reg  LAG ;
reg  LAH ;
reg  LAI ;
reg  LAJ ;
reg  LAK ;
reg  LAL ;
reg  LAM ;
reg  LAN ;
reg  LAO ;
reg  LAP ;
reg  lba ;
reg  lbb ;
reg  lbc ;
reg  lbd ;
reg  lbe ;
reg  lbf ;
reg  lbg ;
reg  lbh ;
reg  lbi ;
reg  lbj ;
reg  lbk ;
reg  lbl ;
reg  lbm ;
reg  lbn ;
reg  lbo ;
reg  lbp ;
reg  lca ;
reg  lcb ;
reg  lcc ;
reg  lcd ;
reg  lce ;
reg  lcf ;
reg  lcg ;
reg  lch ;
reg  lci ;
reg  lcj ;
reg  lck ;
reg  lcl ;
reg  lcm ;
reg  lcn ;
reg  lco ;
reg  lcp ;
reg  lda ;
reg  ldb ;
reg  ldc ;
reg  ldd ;
reg  lde ;
reg  ldf ;
reg  ldg ;
reg  ldh ;
reg  ldi ;
reg  ldj ;
reg  ldk ;
reg  ldl ;
reg  ldm ;
reg  ldn ;
reg  ldo ;
reg  ldp ;
reg  lea ;
reg  leb ;
reg  lec ;
reg  led ;
reg  lee ;
reg  lef ;
reg  leg ;
reg  leh ;
reg  lfa ;
reg  lfb ;
reg  lfc ;
reg  lfd ;
reg  lfe ;
reg  lff ;
reg  lfg ;
reg  lfh ;
reg  lga ;
reg  lgb ;
reg  lgc ;
reg  lgd ;
reg  lge ;
reg  lgf ;
reg  lgg ;
reg  lgh ;
reg  MAA ;
reg  MAC ;
reg  MAD ;
reg  MAE ;
reg  MAF ;
reg  MAG ;
reg  MAH ;
reg  MAI ;
reg  MAJ ;
reg  MAK ;
reg  MAL ;
reg  MAM ;
reg  MAN ;
reg  MAO ;
reg  MAP ;
reg  MBA ;
reg  MBB ;
reg  MBC ;
reg  NAA ;
reg  NAC ;
reg  NAD ;
reg  NAE ;
reg  NAF ;
reg  NAG ;
reg  NAH ;
reg  NAI ;
reg  NAJ ;
reg  NAK ;
reg  NAL ;
reg  NAM ;
reg  NAN ;
reg  NBA ;
reg  NBB ;
reg  NBC ;
reg  NBD ;
reg  NBE ;
reg  NBF ;
reg  NBG ;
reg  NBH ;
reg  NBI ;
reg  NBJ ;
reg  NBK ;
reg  NBL ;
reg  NBM ;
reg  NBN ;
reg  NBO ;
reg  NBP ;
reg  NCA ;
reg  NCC ;
reg  NCD ;
reg  NCE ;
reg  NCF ;
reg  NCG ;
reg  NCH ;
reg  NCI ;
reg  NCJ ;
reg  NCK ;
reg  NCL ;
reg  NCM ;
reg  NCN ;
reg  OAA ;
reg  OAB ;
reg  OAC ;
reg  OAD ;
reg  OAE ;
reg  OAF ;
reg  OAG ;
reg  OAH ;
reg  OAI ;
reg  OAJ ;
reg  OAK ;
reg  OAL ;
reg  OAM ;
reg  OAN ;
reg  OAO ;
reg  OAP ;
reg  OBA ;
reg  OBB ;
reg  OBC ;
reg  OBD ;
reg  OBE ;
reg  OBF ;
reg  OBG ;
reg  OBH ;
reg  OBI ;
reg  OBJ ;
reg  OBK ;
reg  OBL ;
reg  OBM ;
reg  OBN ;
reg  OBO ;
reg  OBP ;
reg  OCA ;
reg  OCB ;
reg  OCC ;
reg  OCD ;
reg  OCE ;
reg  OCF ;
reg  OCG ;
reg  OCH ;
reg  OCI ;
reg  OCJ ;
reg  OCK ;
reg  OCL ;
reg  OCM ;
reg  OCN ;
reg  OCO ;
reg  OCP ;
reg  ODA ;
reg  ODB ;
reg  ODC ;
reg  ODD ;
reg  ODE ;
reg  ODF ;
reg  ODG ;
reg  ODH ;
reg  ODI ;
reg  ODJ ;
reg  ODK ;
reg  ODL ;
reg  ODM ;
reg  ODN ;
reg  ODO ;
reg  ODP ;
reg  OEA ;
reg  OEB ;
reg  OEC ;
reg  OED ;
reg  OEE ;
reg  OEF ;
reg  OEG ;
reg  OEH ;
reg  OEI ;
reg  OEJ ;
reg  OEK ;
reg  OEL ;
reg  OEM ;
reg  OEN ;
reg  OEO ;
reg  OEP ;
reg  OFA ;
reg  OFB ;
reg  OFC ;
reg  OFD ;
reg  OFE ;
reg  OFF ;
reg  OFG ;
reg  OFH ;
reg  OFI ;
reg  OFJ ;
reg  OFK ;
reg  OFL ;
reg  OFM ;
reg  OFN ;
reg  OFO ;
reg  OFP ;
reg  OGA ;
reg  OGB ;
reg  OGC ;
reg  OGD ;
reg  OGE ;
reg  OGF ;
reg  OGG ;
reg  OGH ;
reg  OGI ;
reg  OGJ ;
reg  OGK ;
reg  OGL ;
reg  OGM ;
reg  OGN ;
reg  OGO ;
reg  OGP ;
reg  OHA ;
reg  OHB ;
reg  OHC ;
reg  OHD ;
reg  OHE ;
reg  OHF ;
reg  OHG ;
reg  OHH ;
reg  OHI ;
reg  OHJ ;
reg  OHK ;
reg  OHL ;
reg  OHM ;
reg  OHN ;
reg  OHO ;
reg  OHP ;
reg  OIA ;
reg  OIB ;
reg  OIC ;
reg  OID ;
reg  OIE ;
reg  OIF ;
reg  OIG ;
reg  OIH ;
reg  oja ;
reg  ojb ;
reg  ojc ;
reg  ojd ;
reg  oje ;
reg  OJF ;
reg  OJG ;
reg  OJH ;
reg  OJI ;
reg  OJJ ;
reg  OJK ;
reg  ojl ;
reg  OKA ;
reg  OKB ;
reg  OKC ;
reg  OKD ;
reg  OKE ;
reg  OKF ;
reg  ola ;
reg  olb ;
reg  olc ;
reg  old ;
reg  olf ;
reg  oma ;
reg  omb ;
reg  omc ;
reg  omd ;
reg  omf ;
reg  ona ;
reg  onb ;
reg  onc ;
reg  ond ;
reg  one ;
reg  onf ;
reg  ORA ;
reg  ORB ;
reg  ORC ;
reg  ORD ;
reg  OSA ;
reg  OSB ;
reg  OSC ;
reg  OSD ;
reg  OSE ;
reg  OSF ;
reg  OSG ;
reg  OSH ;
reg  ota ;
reg  oua ;
reg  oub ;
reg  ouc ;
reg  QAA ;
reg  QAB ;
reg  QAC ;
reg  QAD ;
reg  QBA ;
reg  QBB ;
reg  qca ;
reg  qcb ;
reg  qcc ;
reg  qcd ;
reg  qce ;
reg  qda ;
reg  qdb ;
reg  qdc ;
reg  qdd ;
reg  qde ;
reg  qea ;
reg  qeb ;
reg  qec ;
reg  qed ;
reg  qee ;
reg  qef ;
reg  qeg ;
reg  qeh ;
reg  qei ;
reg  qej ;
reg  qek ;
reg  qfa ;
reg  qfb ;
reg  qfc ;
reg  qfd ;
reg  QGA ;
reg  qgb ;
reg  qgc ;
reg  qgd ;
reg  qge ;
reg  qha ;
reg  qhb ;
reg  qhc ;
reg  qhd ;
reg  qhe ;
reg  qhf ;
reg  qhg ;
reg  qhh ;
reg  qhi ;
reg  qhj ;
reg  qhk ;
reg  qhl ;
reg  qhm ;
reg  qhn ;
reg  qho ;
reg  qhp ;
reg  qhq ;
reg  qhr ;
reg  qhs ;
reg  QIA ;
reg  QIB ;
reg  qid ;
reg  QJA ;
reg  QJB ;
reg  qjd ;
reg  QKA ;
reg  QKB ;
reg  qkd ;
reg  QLA ;
reg  QLB ;
reg  QLD ;
reg  qle ;
reg  qma ;
reg  qmb ;
reg  qmc ;
reg  qna ;
reg  QNB ;
reg  qnc ;
reg  QND ;
reg  QNE ;
reg  QNF ;
reg  QOA ;
reg  QOB ;
reg  qod ;
reg  QOF ;
reg  QOG ;
reg  QOH ;
reg  qpa ;
reg  qpb ;
reg  qpc ;
reg  qpe ;
reg  qpf ;
reg  QQA ;
reg  QQB ;
reg  QRA ;
reg  QSA ;
reg  QSB ;
reg  qsd ;
reg  QTA ;
reg  QTB ;
reg  qtc ;
reg  QUA ;
reg  qub ;
reg  quc ;
reg  QVA ;
reg  qvb ;
reg  qvc ;
reg  qvd ;
reg  qve ;
reg  qvf ;
reg  qvg ;
reg  qvh ;
reg  qvi ;
reg  qvj ;
reg  qvk ;
reg  TGL ;
reg  TKA ;
reg  TKB ;
reg  TKC ;
reg  TKD ;
reg  txa ;
reg  txb ;
reg  txc ;
reg  txd ;
reg  txe ;
reg  txf ;
reg  txg ;
reg  txh ;
reg  vaa ;
reg  VAB ;
reg  VAC ;
reg  VAD ;
reg  VAE ;
reg  VAF ;
reg  VAG ;
reg  VAH ;
reg  VAI ;
reg  VAJ ;
reg  VAK ;
reg  VAL ;
reg  VAM ;
reg  VAN ;
reg  vba ;
reg  VBB ;
reg  VBC ;
reg  VBD ;
reg  VBE ;
reg  VBF ;
reg  VBG ;
reg  VBH ;
reg  VBI ;
reg  VBJ ;
reg  VBK ;
reg  VBL ;
reg  VBM ;
reg  VBN ;
reg  vca ;
reg  VCB ;
reg  VCC ;
reg  VCD ;
reg  VCE ;
reg  VCF ;
reg  VCG ;
reg  VCH ;
reg  VCI ;
reg  VCJ ;
reg  VCK ;
reg  VCL ;
reg  VCM ;
reg  VCN ;
reg  vda ;
reg  VDB ;
reg  VDC ;
reg  VDD ;
reg  VDE ;
reg  VDF ;
reg  VDG ;
reg  VDH ;
reg  VDI ;
reg  VDJ ;
reg  VDK ;
reg  VDL ;
reg  VDM ;
reg  VDN ;
reg  vea ;
reg  VEB ;
reg  VEC ;
reg  VED ;
reg  VEE ;
reg  VEF ;
reg  VEG ;
reg  VEH ;
reg  VEI ;
reg  VEJ ;
reg  VEK ;
reg  VEL ;
reg  VEM ;
reg  VEN ;
reg  vfa ;
reg  VFB ;
reg  VFC ;
reg  VFD ;
reg  VFE ;
reg  VFF ;
reg  VFG ;
reg  VFH ;
reg  VFI ;
reg  VFJ ;
reg  VFK ;
reg  VFL ;
reg  VFM ;
reg  VFN ;
reg  vga ;
reg  VGB ;
reg  VGC ;
reg  VGD ;
reg  VGE ;
reg  VGF ;
reg  VGG ;
reg  VGH ;
reg  VGI ;
reg  VGJ ;
reg  VGK ;
reg  VGL ;
reg  VGM ;
reg  VGN ;
reg  vha ;
reg  VHB ;
reg  VHC ;
reg  VHD ;
reg  VHE ;
reg  VHF ;
reg  VHG ;
reg  VHH ;
reg  VHI ;
reg  VHJ ;
reg  VHK ;
reg  VHL ;
reg  VHM ;
reg  VHN ;
wire  aaa ;
wire  aab ;
wire  aac ;
wire  aad ;
wire  aae ;
wire  aaf ;
wire  aag ;
wire  aah ;
wire  aai ;
wire  aaj ;
wire  aak ;
wire  aal ;
wire  aam ;
wire  aan ;
wire  aao ;
wire  aap ;
wire  aba ;
wire  abb ;
wire  abc ;
wire  abd ;
wire  abe ;
wire  abf ;
wire  abg ;
wire  abh ;
wire  abi ;
wire  abj ;
wire  abk ;
wire  abl ;
wire  abm ;
wire  abn ;
wire  abo ;
wire  abp ;
wire  baa ;
wire  bab ;
wire  bac ;
wire  bad ;
wire  bae ;
wire  baf ;
wire  BAI ;
wire  BAJ ;
wire  BAK ;
wire  BAL ;
wire  BAM ;
wire  BAN ;
wire  BBA ;
wire  BBB ;
wire  BBC ;
wire  BBD ;
wire  BBE ;
wire  BBF ;
wire  BBG ;
wire  bbh ;
wire  BBH ;
wire  BBI ;
wire  BBJ ;
wire  BBK ;
wire  BBL ;
wire  BBM ;
wire  BBN ;
wire  BBO ;
wire  bbp ;
wire  BBP ;
wire  BCA ;
wire  BCB ;
wire  BCC ;
wire  BCD ;
wire  BCE ;
wire  BCF ;
wire  BCG ;
wire  bch ;
wire  BCH ;
wire  BDA ;
wire  BDB ;
wire  BDC ;
wire  BDD ;
wire  BDE ;
wire  BDF ;
wire  BDG ;
wire  bdh ;
wire  BDH ;
wire  BDI ;
wire  BDJ ;
wire  BDK ;
wire  BDL ;
wire  BDM ;
wire  BDN ;
wire  BDO ;
wire  BDP ;
wire  BEA ;
wire  BEB ;
wire  BEC ;
wire  BED ;
wire  BEE ;
wire  BEF ;
wire  BEG ;
wire  BEH ;
wire  caa ;
wire  cab ;
wire  cac ;
wire  cad ;
wire  cae ;
wire  caf ;
wire  cba ;
wire  cbb ;
wire  cbc ;
wire  cbd ;
wire  cbe ;
wire  cbf ;
wire  cca ;
wire  ccb ;
wire  ccc ;
wire  ccd ;
wire  cce ;
wire  ccf ;
wire  cda ;
wire  cdb ;
wire  cdc ;
wire  cdd ;
wire  cde ;
wire  cdf ;
wire  cea ;
wire  ceb ;
wire  cec ;
wire  ced ;
wire  cee ;
wire  cef ;
wire  cfa ;
wire  cfb ;
wire  cfc ;
wire  cfd ;
wire  cfe ;
wire  cff ;
wire  daa ;
wire  DAA ;
wire  dab ;
wire  DAB ;
wire  dac ;
wire  DAC ;
wire  dad ;
wire  DAD ;
wire  dae ;
wire  DAE ;
wire  daf ;
wire  DAF ;
wire  dag ;
wire  DAG ;
wire  dah ;
wire  DAH ;
wire  dba ;
wire  DBA ;
wire  dbb ;
wire  DBB ;
wire  dbc ;
wire  DBC ;
wire  dbd ;
wire  DBD ;
wire  dbe ;
wire  DBE ;
wire  dbf ;
wire  DBF ;
wire  dbg ;
wire  DBG ;
wire  dbh ;
wire  DBH ;
wire  dca ;
wire  DCA ;
wire  dcb ;
wire  DCB ;
wire  dcc ;
wire  DCC ;
wire  dcd ;
wire  DCD ;
wire  dce ;
wire  DCE ;
wire  dcf ;
wire  DCF ;
wire  dcg ;
wire  DCG ;
wire  dch ;
wire  DCH ;
wire  dda ;
wire  DDA ;
wire  ddb ;
wire  DDB ;
wire  ddc ;
wire  DDC ;
wire  ddd ;
wire  DDD ;
wire  dde ;
wire  DDE ;
wire  ddf ;
wire  DDF ;
wire  ddg ;
wire  DDG ;
wire  ddh ;
wire  DDH ;
wire  dea ;
wire  DEA ;
wire  deb ;
wire  DEB ;
wire  dec ;
wire  DEC ;
wire  ded ;
wire  DED ;
wire  dee ;
wire  DEE ;
wire  def ;
wire  DEF ;
wire  deg ;
wire  DEG ;
wire  dfa ;
wire  DFA ;
wire  dfb ;
wire  DFB ;
wire  dfc ;
wire  DFC ;
wire  dfd ;
wire  DFD ;
wire  dfe ;
wire  DFE ;
wire  dff ;
wire  DFF ;
wire  dfg ;
wire  DFG ;
wire  dfh ;
wire  DFH ;
wire  EAA ;
wire  EAB ;
wire  EAC ;
wire  EAD ;
wire  EAE ;
wire  EAF ;
wire  EAG ;
wire  EAH ;
wire  EAI ;
wire  EAJ ;
wire  EAK ;
wire  EAL ;
wire  EAM ;
wire  EAN ;
wire  EAO ;
wire  EAP ;
wire  EBJ ;
wire  EBK ;
wire  EBL ;
wire  EBM ;
wire  EBN ;
wire  EBO ;
wire  EBP ;
wire  ECM ;
wire  ECN ;
wire  ECO ;
wire  ECP ;
wire  faa ;
wire  FAA ;
wire  fab ;
wire  FAB ;
wire  fac ;
wire  FAC ;
wire  fad ;
wire  FAD ;
wire  fae ;
wire  FAE ;
wire  faf ;
wire  FAF ;
wire  fag ;
wire  FAG ;
wire  fah ;
wire  FAH ;
wire  fai ;
wire  FAI ;
wire  faj ;
wire  FAJ ;
wire  fak ;
wire  FAK ;
wire  fal ;
wire  FAL ;
wire  fam ;
wire  FAM ;
wire  fan ;
wire  FAN ;
wire  fap ;
wire  FAP ;
wire  fba ;
wire  FBA ;
wire  fbb ;
wire  FBB ;
wire  fbc ;
wire  FBC ;
wire  fbd ;
wire  FBD ;
wire  fbe ;
wire  FBE ;
wire  fbf ;
wire  FBF ;
wire  fbh ;
wire  FBH ;
wire  fbi ;
wire  FBI ;
wire  fbj ;
wire  FBJ ;
wire  fbk ;
wire  FBK ;
wire  fbl ;
wire  FBL ;
wire  fbm ;
wire  FBM ;
wire  fbn ;
wire  FBN ;
wire  fbo ;
wire  FBO ;
wire  fbp ;
wire  FBP ;
wire  gaa ;
wire  gab ;
wire  gac ;
wire  gad ;
wire  gae ;
wire  gaf ;
wire  gag ;
wire  gah ;
wire  gai ;
wire  gaj ;
wire  gak ;
wire  GBA ;
wire  GBB ;
wire  GBC ;
wire  GBD ;
wire  GBE ;
wire  GBF ;
wire  GBG ;
wire  GBH ;
wire  GBK ;
wire  GBL ;
wire  GBN ;
wire  GBO ;
wire  GCA ;
wire  GCB ;
wire  GCC ;
wire  GCD ;
wire  GCE ;
wire  GCF ;
wire  GCH ;
wire  GCI ;
wire  GCJ ;
wire  GCK ;
wire  GCL ;
wire  GCM ;
wire  GCN ;
wire  GCO ;
wire  GCP ;
wire  GDA ;
wire  GDB ;
wire  GDC ;
wire  iaa ;
wire  iab ;
wire  iac ;
wire  iad ;
wire  iae ;
wire  iaf ;
wire  iag ;
wire  iah ;
wire  iai ;
wire  iaj ;
wire  iak ;
wire  ial ;
wire  iam ;
wire  ian ;
wire  iao ;
wire  iap ;
wire  iba ;
wire  ibb ;
wire  ibc ;
wire  ibd ;
wire  ibe ;
wire  ibf ;
wire  ibg ;
wire  ibh ;
wire  ibi ;
wire  ibj ;
wire  ibk ;
wire  ibl ;
wire  ibm ;
wire  ibn ;
wire  ibo ;
wire  ibp ;
wire  ica ;
wire  icb ;
wire  icc ;
wire  icd ;
wire  ice ;
wire  icf ;
wire  icg ;
wire  ich ;
wire  ici ;
wire  icj ;
wire  ick ;
wire  icl ;
wire  icm ;
wire  icn ;
wire  ico ;
wire  icp ;
wire  ida ;
wire  idb ;
wire  idc ;
wire  idd ;
wire  ide ;
wire  idf ;
wire  iea ;
wire  ieb ;
wire  ifa ;
wire  iga ;
wire  iha ;
wire  ihb ;
wire  ihf ;
wire  ija ;
wire  ika ;
wire  ikb ;
wire  ikc ;
wire  ikd ;
wire  ike ;
wire  ikf ;
wire  ikg ;
wire  ikh ;
wire  ila ;
wire  jaa ;
wire  JAA ;
wire  jab ;
wire  JAB ;
wire  jac ;
wire  JAC ;
wire  jba ;
wire  JBA ;
wire  jbb ;
wire  JBB ;
wire  jbc ;
wire  JBC ;
wire  jbd ;
wire  JBD ;
wire  jbe ;
wire  JBE ;
wire  jbf ;
wire  JBF ;
wire  jbg ;
wire  JBG ;
wire  jbh ;
wire  JBH ;
wire  jca ;
wire  JCA ;
wire  jcb ;
wire  JCB ;
wire  jcc ;
wire  JCC ;
wire  jcd ;
wire  JCD ;
wire  jcf ;
wire  JCF ;
wire  jcg ;
wire  JCG ;
wire  jch ;
wire  JCH ;
wire  jci ;
wire  JCI ;
wire  jcj ;
wire  JCJ ;
wire  jda ;
wire  JDA ;
wire  jdb ;
wire  JDB ;
wire  jdc ;
wire  JDC ;
wire  jea ;
wire  JEA ;
wire  jeb ;
wire  JEB ;
wire  JFA ;
wire  JFB ;
wire  JFC ;
wire  JFD ;
wire  JFE ;
wire  JFF ;
wire  JFG ;
wire  JFH ;
wire  jfi ;
wire  JGA ;
wire  JGB ;
wire  JGC ;
wire  JGD ;
wire  JGE ;
wire  JGF ;
wire  JGG ;
wire  JGH ;
wire  jgi ;
wire  laa ;
wire  lab ;
wire  lac ;
wire  lad ;
wire  lae ;
wire  laf ;
wire  lag ;
wire  lah ;
wire  lai ;
wire  laj ;
wire  lak ;
wire  lal ;
wire  lam ;
wire  lan ;
wire  lao ;
wire  lap ;
wire  LBA ;
wire  LBB ;
wire  LBC ;
wire  LBD ;
wire  LBE ;
wire  LBF ;
wire  LBG ;
wire  LBH ;
wire  LBI ;
wire  LBJ ;
wire  LBK ;
wire  LBL ;
wire  LBM ;
wire  LBN ;
wire  LBO ;
wire  LBP ;
wire  LCA ;
wire  LCB ;
wire  LCC ;
wire  LCD ;
wire  LCE ;
wire  LCF ;
wire  LCG ;
wire  LCH ;
wire  LCI ;
wire  LCJ ;
wire  LCK ;
wire  LCL ;
wire  LCM ;
wire  LCN ;
wire  LCO ;
wire  LCP ;
wire  LDA ;
wire  LDB ;
wire  LDC ;
wire  LDD ;
wire  LDE ;
wire  LDF ;
wire  LDG ;
wire  LDH ;
wire  LDI ;
wire  LDJ ;
wire  LDK ;
wire  LDL ;
wire  LDM ;
wire  LDN ;
wire  LDO ;
wire  LDP ;
wire  LEA ;
wire  LEB ;
wire  LEC ;
wire  LED ;
wire  LEE ;
wire  LEF ;
wire  LEG ;
wire  LEH ;
wire  LFA ;
wire  LFB ;
wire  LFC ;
wire  LFD ;
wire  LFE ;
wire  LFF ;
wire  LFG ;
wire  LFH ;
wire  LGA ;
wire  LGB ;
wire  LGC ;
wire  LGD ;
wire  LGE ;
wire  LGF ;
wire  LGG ;
wire  LGH ;
wire  maa ;
wire  mac ;
wire  mad ;
wire  mae ;
wire  maf ;
wire  mag ;
wire  mah ;
wire  mai ;
wire  maj ;
wire  mak ;
wire  mal ;
wire  mam ;
wire  man ;
wire  mao ;
wire  map ;
wire  mba ;
wire  mbb ;
wire  mbc ;
wire  naa ;
wire  nac ;
wire  nad ;
wire  nae ;
wire  naf ;
wire  nag ;
wire  nah ;
wire  nai ;
wire  naj ;
wire  nak ;
wire  nal ;
wire  nam ;
wire  nan ;
wire  nba ;
wire  nbb ;
wire  nbc ;
wire  nbd ;
wire  nbe ;
wire  nbf ;
wire  nbg ;
wire  nbh ;
wire  nbi ;
wire  nbj ;
wire  nbk ;
wire  nbl ;
wire  nbm ;
wire  nbn ;
wire  nbo ;
wire  nbp ;
wire  nca ;
wire  ncc ;
wire  ncd ;
wire  nce ;
wire  ncf ;
wire  ncg ;
wire  nch ;
wire  nci ;
wire  ncj ;
wire  nck ;
wire  ncl ;
wire  ncm ;
wire  ncn ;
wire  oaa ;
wire  oab ;
wire  oac ;
wire  oad ;
wire  oae ;
wire  oaf ;
wire  oag ;
wire  oah ;
wire  oai ;
wire  oaj ;
wire  oak ;
wire  oal ;
wire  oam ;
wire  oan ;
wire  oao ;
wire  oap ;
wire  oba ;
wire  obb ;
wire  obc ;
wire  obd ;
wire  obe ;
wire  obf ;
wire  obg ;
wire  obh ;
wire  obi ;
wire  obj ;
wire  obk ;
wire  obl ;
wire  obm ;
wire  obn ;
wire  obo ;
wire  obp ;
wire  oca ;
wire  ocb ;
wire  occ ;
wire  ocd ;
wire  oce ;
wire  ocf ;
wire  ocg ;
wire  och ;
wire  oci ;
wire  ocj ;
wire  ock ;
wire  ocl ;
wire  ocm ;
wire  ocn ;
wire  oco ;
wire  ocp ;
wire  oda ;
wire  odb ;
wire  odc ;
wire  odd ;
wire  ode ;
wire  odf ;
wire  odg ;
wire  odh ;
wire  odi ;
wire  odj ;
wire  odk ;
wire  odl ;
wire  odm ;
wire  odn ;
wire  odo ;
wire  odp ;
wire  oea ;
wire  oeb ;
wire  oec ;
wire  oed ;
wire  oee ;
wire  oef ;
wire  oeg ;
wire  oeh ;
wire  oei ;
wire  oej ;
wire  oek ;
wire  oel ;
wire  oem ;
wire  oen ;
wire  oeo ;
wire  oep ;
wire  ofa ;
wire  ofb ;
wire  ofc ;
wire  ofd ;
wire  ofe ;
wire  off ;
wire  ofg ;
wire  ofh ;
wire  ofi ;
wire  ofj ;
wire  ofk ;
wire  ofl ;
wire  ofm ;
wire  ofn ;
wire  ofo ;
wire  ofp ;
wire  oga ;
wire  ogb ;
wire  ogc ;
wire  ogd ;
wire  oge ;
wire  ogf ;
wire  ogg ;
wire  ogh ;
wire  ogi ;
wire  ogj ;
wire  ogk ;
wire  ogl ;
wire  ogm ;
wire  ogn ;
wire  ogo ;
wire  ogp ;
wire  oha ;
wire  ohb ;
wire  ohc ;
wire  ohd ;
wire  ohe ;
wire  ohf ;
wire  ohg ;
wire  ohh ;
wire  ohi ;
wire  ohj ;
wire  ohk ;
wire  ohl ;
wire  ohm ;
wire  ohn ;
wire  oho ;
wire  ohp ;
wire  oia ;
wire  oib ;
wire  oic ;
wire  oid ;
wire  oie ;
wire  oif ;
wire  oig ;
wire  oih ;
wire  OJA ;
wire  OJB ;
wire  OJC ;
wire  OJD ;
wire  OJE ;
wire  ojf ;
wire  ojg ;
wire  ojh ;
wire  oji ;
wire  ojj ;
wire  ojk ;
wire  OJL ;
wire  oka ;
wire  okb ;
wire  okc ;
wire  okd ;
wire  oke ;
wire  okf ;
wire  OLA ;
wire  OLB ;
wire  OLC ;
wire  OLD ;
wire  OLF ;
wire  OMA ;
wire  OMB ;
wire  OMC ;
wire  OMD ;
wire  OMF ;
wire  ONA ;
wire  ONB ;
wire  ONC ;
wire  OND ;
wire  ONE ;
wire  ONF ;
wire  ora ;
wire  orb ;
wire  orc ;
wire  ord ;
wire  osa ;
wire  osb ;
wire  osc ;
wire  osd ;
wire  ose ;
wire  osf ;
wire  osg ;
wire  osh ;
wire  OTA ;
wire  OUA ;
wire  OUB ;
wire  OUC ;
wire  qaa ;
wire  qab ;
wire  qac ;
wire  qad ;
wire  qba ;
wire  qbb ;
wire  QCA ;
wire  QCB ;
wire  QCC ;
wire  QCD ;
wire  QCE ;
wire  QDA ;
wire  QDB ;
wire  QDC ;
wire  QDD ;
wire  QDE ;
wire  QEA ;
wire  QEB ;
wire  QEC ;
wire  QED ;
wire  QEE ;
wire  QEF ;
wire  QEG ;
wire  QEH ;
wire  QEI ;
wire  QEJ ;
wire  QEK ;
wire  QFA ;
wire  QFB ;
wire  QFC ;
wire  QFD ;
wire  qga ;
wire  QGB ;
wire  QGC ;
wire  QGD ;
wire  QGE ;
wire  QHA ;
wire  QHB ;
wire  QHC ;
wire  QHD ;
wire  QHE ;
wire  QHF ;
wire  QHG ;
wire  QHH ;
wire  QHI ;
wire  QHJ ;
wire  QHK ;
wire  QHL ;
wire  QHM ;
wire  QHN ;
wire  QHO ;
wire  QHP ;
wire  QHQ ;
wire  QHR ;
wire  QHS ;
wire  qia ;
wire  qib ;
wire  QID ;
wire  qja ;
wire  qjb ;
wire  QJD ;
wire  qka ;
wire  qkb ;
wire  QKD ;
wire  qla ;
wire  qlb ;
wire  qld ;
wire  QLE ;
wire  QMA ;
wire  QMB ;
wire  QMC ;
wire  QNA ;
wire  qnb ;
wire  QNC ;
wire  qnd ;
wire  qne ;
wire  qnf ;
wire  qoa ;
wire  qob ;
wire  QOD ;
wire  qof ;
wire  qog ;
wire  qoh ;
wire  QPA ;
wire  QPB ;
wire  QPC ;
wire  QPE ;
wire  QPF ;
wire  qqa ;
wire  qqb ;
wire  qra ;
wire  qsa ;
wire  qsb ;
wire  QSD ;
wire  qta ;
wire  qtb ;
wire  QTC ;
wire  qua ;
wire  QUB ;
wire  QUC ;
wire  qva ;
wire  QVB ;
wire  QVC ;
wire  QVD ;
wire  QVE ;
wire  QVF ;
wire  QVG ;
wire  QVH ;
wire  QVI ;
wire  QVJ ;
wire  QVK ;
wire  taa ;
wire  TAA ;
wire  tab ;
wire  TAB ;
wire  tac ;
wire  TAC ;
wire  tad ;
wire  TAD ;
wire  tae ;
wire  TAE ;
wire  taf ;
wire  TAF ;
wire  tag ;
wire  TAG ;
wire  tah ;
wire  TAH ;
wire  tai ;
wire  TAI ;
wire  taj ;
wire  TAJ ;
wire  tak ;
wire  TAK ;
wire  tal ;
wire  TAL ;
wire  tam ;
wire  TAM ;
wire  tan ;
wire  TAN ;
wire  tao ;
wire  TAO ;
wire  tap ;
wire  TAP ;
wire  taq ;
wire  TAQ ;
wire  tar ;
wire  TAR ;
wire  tas ;
wire  TAS ;
wire  tat ;
wire  TAT ;
wire  tau ;
wire  TAU ;
wire  tav ;
wire  TAV ;
wire  taw ;
wire  TAW ;
wire  tax ;
wire  TAX ;
wire  tba ;
wire  TBA ;
wire  tbb ;
wire  TBB ;
wire  tbc ;
wire  TBC ;
wire  tbd ;
wire  TBD ;
wire  tbi ;
wire  TBI ;
wire  tbj ;
wire  TBJ ;
wire  tbk ;
wire  TBK ;
wire  tbl ;
wire  TBL ;
wire  tca ;
wire  TCA ;
wire  tcb ;
wire  TCB ;
wire  tda ;
wire  TDA ;
wire  tdb ;
wire  TDB ;
wire  tea ;
wire  TEA ;
wire  teb ;
wire  TEB ;
wire  tga ;
wire  TGA ;
wire  tgb ;
wire  TGB ;
wire  tgc ;
wire  TGC ;
wire  tgd ;
wire  TGD ;
wire  tge ;
wire  TGE ;
wire  tgf ;
wire  TGF ;
wire  tgg ;
wire  TGG ;
wire  tgh ;
wire  TGH ;
wire  tgi ;
wire  TGI ;
wire  tgj ;
wire  TGJ ;
wire  tgk ;
wire  TGK ;
wire  tgl ;
wire  tha ;
wire  THA ;
wire  thb ;
wire  THB ;
wire  thc ;
wire  THC ;
wire  thd ;
wire  THD ;
wire  the ;
wire  THE ;
wire  thf ;
wire  THF ;
wire  thg ;
wire  THG ;
wire  thh ;
wire  THH ;
wire  thi ;
wire  THI ;
wire  thj ;
wire  THJ ;
wire  thk ;
wire  THK ;
wire  thl ;
wire  THL ;
wire  thm ;
wire  THM ;
wire  thn ;
wire  THN ;
wire  tho ;
wire  THO ;
wire  thp ;
wire  THP ;
wire  thq ;
wire  THQ ;
wire  thr ;
wire  THR ;
wire  ths ;
wire  THS ;
wire  tht ;
wire  THT ;
wire  tka ;
wire  tkb ;
wire  tkc ;
wire  tkd ;
wire  TXA ;
wire  TXB ;
wire  TXC ;
wire  TXD ;
wire  TXE ;
wire  TXF ;
wire  TXG ;
wire  TXH ;
wire  VAA ;
wire  vab ;
wire  vac ;
wire  vad ;
wire  vae ;
wire  vaf ;
wire  vag ;
wire  vah ;
wire  vai ;
wire  vaj ;
wire  vak ;
wire  val ;
wire  vam ;
wire  van ;
wire  VBA ;
wire  vbb ;
wire  vbc ;
wire  vbd ;
wire  vbe ;
wire  vbf ;
wire  vbg ;
wire  vbh ;
wire  vbi ;
wire  vbj ;
wire  vbk ;
wire  vbl ;
wire  vbm ;
wire  vbn ;
wire  VCA ;
wire  vcb ;
wire  vcc ;
wire  vcd ;
wire  vce ;
wire  vcf ;
wire  vcg ;
wire  vch ;
wire  vci ;
wire  vcj ;
wire  vck ;
wire  vcl ;
wire  vcm ;
wire  vcn ;
wire  VDA ;
wire  vdb ;
wire  vdc ;
wire  vdd ;
wire  vde ;
wire  vdf ;
wire  vdg ;
wire  vdh ;
wire  vdi ;
wire  vdj ;
wire  vdk ;
wire  vdl ;
wire  vdm ;
wire  vdn ;
wire  VEA ;
wire  veb ;
wire  vec ;
wire  ved ;
wire  vee ;
wire  vef ;
wire  veg ;
wire  veh ;
wire  vei ;
wire  vej ;
wire  vek ;
wire  vel ;
wire  vem ;
wire  ven ;
wire  VFA ;
wire  vfb ;
wire  vfc ;
wire  vfd ;
wire  vfe ;
wire  vff ;
wire  vfg ;
wire  vfh ;
wire  vfi ;
wire  vfj ;
wire  vfk ;
wire  vfl ;
wire  vfm ;
wire  vfn ;
wire  VGA ;
wire  vgb ;
wire  vgc ;
wire  vgd ;
wire  vge ;
wire  vgf ;
wire  vgg ;
wire  vgh ;
wire  vgi ;
wire  vgj ;
wire  vgk ;
wire  vgl ;
wire  vgm ;
wire  vgn ;
wire  VHA ;
wire  vhb ;
wire  vhc ;
wire  vhd ;
wire  vhe ;
wire  vhf ;
wire  vhg ;
wire  vhh ;
wire  vhi ;
wire  vhj ;
wire  vhk ;
wire  vhl ;
wire  vhm ;
wire  vhn ;
wire  yya ;
wire  YYA ;
wire  yym ;
wire  YYM ;
wire  ZZI ;
wire  ZZO ;
assign ZZI = 1'b1;
assign ZZO = 1'b0;
assign VAA = ~vaa;  //complement 
assign vac = ~VAC;  //complement 
assign vae = ~VAE;  //complement 
assign vag = ~VAG;  //complement 
assign vah = ~VAH;  //complement 
assign vad = ~VAD;  //complement 
assign vaf = ~VAF;  //complement 
assign vai = ~VAI;  //complement 
assign vaj = ~VAJ;  //complement 
assign maa = ~MAA;  //complement 
assign mbc = ~MBC;  //complement 
assign naa = ~NAA;  //complement 
assign caa = ~CAA;  //complement 
assign cab = ~CAB;  //complement 
assign cac = ~CAC;  //complement 
assign daa = caa & ~( ZZI  ) | CAA & ( ZZI  );
assign DAA = ~daa ;
assign dab = cab & ~( caa & ZZI  ) | CAB & ( caa & ZZI  );
assign DAB = ~dab ;  //complement 
assign dac = cac & ~( cab & caa & ZZI  ) | CAC & ( cab & caa & ZZI  );
assign DAC = ~dac;  //complement;
assign DAG =  CAA & cab & cac & cad & cae & caf  ; 
assign dag = ~DAG;  //complement  
assign cad = ~CAD;  //complement 
assign cae = ~CAE;  //complement 
assign caf = ~CAF;  //complement 
assign dad = cad & ~( cac & cab & caa  ) | CAD & ( cac & cab & caa  );
assign DAD = ~dad ;
assign dae = cae & ~( cad & cac & cab & caa  ) | CAE & ( cad & cac & cab & caa  );
assign DAE = ~dae ;  //complement 
assign daf = caf & ~( cae & cad & cac & cab & caa  ) | CAF & ( cae & cad & cac & cab & caa  );
assign DAF = ~daf;  //complement;
assign dah =  caa & cab  |  CAC  |  CAD  |  CAE  |  CAF  ;
assign DAH = ~dah;  //complement 
assign nba = ~NBA;  //complement 
assign nbi = ~NBI;  //complement 
assign nca = ~NCA;  //complement 
assign vab = ~VAB;  //complement 
assign gaa = ~GAA;  //complement 
assign gai = ~GAI;  //complement 
assign FAA =  eap & eao & EAN & eam  ; 
assign faa = ~FAA;  //complement  
assign FBA =  eaj & eak  ; 
assign fba = ~FBA;  //complement 
assign vak = ~VAK;  //complement 
assign val = ~VAL;  //complement 
assign GBA = ~gba;  //complement 
assign GDA = ~gda;  //complement 
assign vam = ~VAM;  //complement 
assign van = ~VAN;  //complement 
assign GCA = ~gca;  //complement 
assign GCI = ~gci;  //complement 
assign FAI =  EBP & EBO & EBN & EBM  ; 
assign fai = ~FAI;  //complement  
assign FBI =  EBL & EBK  ; 
assign fbi = ~FBI;  //complement 
assign QHA = ~qha;  //complement 
assign qia = ~QIA;  //complement 
assign qib = ~QIB;  //complement 
assign QID = ~qid;  //complement 
assign oka = ~OKA;  //complement 
assign EAA = ~eaa;  //complement 
assign EAI = ~eai;  //complement 
assign laa = ~LAA;  //complement 
assign lai = ~LAI;  //complement 
assign oaa = ~OAA;  //complement 
assign oea = ~OEA;  //complement 
assign oei = ~OEI;  //complement 
assign LEA = ~lea;  //complement 
assign LEB = ~leb;  //complement 
assign LFA = ~lfa;  //complement 
assign LFB = ~lfb;  //complement 
assign LGA = ~lga;  //complement 
assign LGB = ~lgb;  //complement 
assign oai = ~OAI;  //complement 
assign oia = ~OIA;  //complement 
assign BAI = ~bai;  //complement 
assign LBA = ~lba;  //complement 
assign LCA = ~lca;  //complement 
assign LDA = ~lda;  //complement 
assign baa = ~BAA;  //complement 
assign LBI = ~lbi;  //complement 
assign LCI = ~lci;  //complement 
assign LDI = ~ldi;  //complement 
assign oba = ~OBA;  //complement 
assign ofa = ~OFA;  //complement 
assign ofi = ~OFI;  //complement 
assign THK = QDE; 
assign thk = ~THK; //complement 
assign THL = QDE; 
assign thl = ~THL;  //complement 
assign THM = QEF; 
assign thm = ~THM;  //complement 
assign THN = QEF; 
assign thn = ~THN;  //complement 
assign obi = ~OBI;  //complement 
assign OLA = ~ola;  //complement 
assign OMA = ~oma;  //complement 
assign ONA = ~ona;  //complement 
assign QGB = ~qgb;  //complement 
assign QGD = ~qgd;  //complement 
assign qta = ~QTA;  //complement 
assign qtb = ~QTB;  //complement 
assign oca = ~OCA;  //complement 
assign oci = ~OCI;  //complement 
assign aaa = ~AAA;  //complement 
assign aai = ~AAI;  //complement 
assign oga = ~OGA;  //complement 
assign ogi = ~OGI;  //complement 
assign BBA = ~bba;  //complement 
assign BBI = ~bbi;  //complement 
assign BCA = ~bca;  //complement 
assign BDA = ~bda;  //complement 
assign tbd = qge & qgd ; 
assign TBD = ~tbd ; //complement 
assign tbl = qge & qgd ; 
assign TBL = ~tbl ;  //complement 
assign osa = ~OSA;  //complement 
assign tbj = qga & qgb ; 
assign TBJ = ~tbj ; //complement 
assign tbb = qga & qgb ; 
assign TBB = ~tbb ;  //complement 
assign BDI = ~bdi;  //complement 
assign BEA = ~bea;  //complement 
assign oda = ~ODA;  //complement 
assign odi = ~ODI;  //complement 
assign aba = ~ABA;  //complement 
assign abi = ~ABI;  //complement 
assign oha = ~OHA;  //complement 
assign ohi = ~OHI;  //complement 
assign VBA = ~vba;  //complement 
assign vbc = ~VBC;  //complement 
assign vbe = ~VBE;  //complement 
assign vbg = ~VBG;  //complement 
assign vbh = ~VBH;  //complement 
assign vbd = ~VBD;  //complement 
assign vbf = ~VBF;  //complement 
assign vbi = ~VBI;  //complement 
assign vbj = ~VBJ;  //complement 
assign mac = ~MAC;  //complement 
assign mah = ~MAH;  //complement 
assign ncc = ~NCC;  //complement 
assign QSD = ~qsd;  //complement 
assign cba = ~CBA;  //complement 
assign cbb = ~CBB;  //complement 
assign cbc = ~CBC;  //complement 
assign dba = cba & ~( ZZI  ) | CBA & ( ZZI  );
assign DBA = ~dba ;
assign dbb = cbb & ~( cba & ZZI  ) | CBB & ( cba & ZZI  );
assign DBB = ~dbb ;  //complement 
assign dbc = cbc & ~( cbb & cba & ZZI  ) | CBC & ( cbb & cba & ZZI  );
assign DBC = ~dbc;  //complement;
assign DBG =  CBA & cbb & cbc & cbd & cbe & cbf  ; 
assign dbg = ~DBG;  //complement  
assign cbd = ~CBD;  //complement 
assign cbe = ~CBE;  //complement 
assign cbf = ~CBF;  //complement 
assign dbd = cbd & ~( cbc & cbb & cba  ) | CBD & ( cbc & cbb & cba  );
assign DBD = ~dbd ;
assign dbe = cbe & ~( cbd & cbc & cbb & cba  ) | CBE & ( cbd & cbc & cbb & cba  );
assign DBE = ~dbe ;  //complement 
assign dbf = cbf & ~( cbe & cbd & cbc & cbb & cba  ) | CBF & ( cbe & cbd & cbc & cbb & cba  );
assign DBF = ~dbf;  //complement;
assign dbh =  cba & cbb  |  CBC  |  CBD  |  CBE  |  CBF  ;
assign DBH = ~dbh;  //complement 
assign mai = ~MAI;  //complement 
assign maj = ~MAJ;  //complement 
assign mak = ~MAK;  //complement 
assign mal = ~MAL;  //complement 
assign nci = ~NCI;  //complement 
assign ncj = ~NCJ;  //complement 
assign nck = ~NCK;  //complement 
assign ncl = ~NCL;  //complement 
assign mam = ~MAM;  //complement 
assign ncm = ~NCM;  //complement 
assign ncn = ~NCN;  //complement 
assign man = ~MAN;  //complement 
assign nbb = ~NBB;  //complement 
assign nbj = ~NBJ;  //complement 
assign nch = ~NCH;  //complement 
assign vbb = ~VBB;  //complement 
assign lak = ~LAK;  //complement 
assign gab = ~GAB;  //complement 
assign gaj = ~GAJ;  //complement 
assign FAB =  EAP & eao & ean & EAM  ; 
assign fab = ~FAB;  //complement  
assign FBB =  EAL & EAK  ; 
assign fbb = ~FBB;  //complement 
assign vbk = ~VBK;  //complement 
assign vbl = ~VBL;  //complement 
assign GBB = ~gbb;  //complement 
assign jcg =  gcb & gcc  ; 
assign JCG = ~jcg;  //complement 
assign vbm = ~VBM;  //complement 
assign vbn = ~VBN;  //complement 
assign LDK = ~ldk;  //complement 
assign GCB = ~gcb;  //complement 
assign GCJ = ~gcj;  //complement 
assign FAJ =  EBP & EBO & EBN & ebm  ; 
assign faj = ~FAJ;  //complement  
assign FBJ =  EBL & ebk  ; 
assign fbj = ~FBJ;  //complement 
assign jcf =  YYA  |  gca  ; 
assign JCF = ~jcf;  //complement 
assign JCC =  GBK & YYM  |  GCA & YYA  ; 
assign jcc = ~JCC;  //complement 
assign jch =  YYM  |  gbk  ; 
assign JCH = ~jch;  //complement 
assign QHI = ~qhi;  //complement 
assign QHJ = ~qhj;  //complement 
assign QHK = ~qhk;  //complement 
assign QHM = ~qhm;  //complement 
assign QHG = ~qhg;  //complement 
assign QHH = ~qhh;  //complement 
assign jca =  gbh  ; 
assign JCA = ~jca;  //complement 
assign jcb =  gcj & gco  ; 
assign JCB = ~jcb;  //complement 
assign QHB = ~qhb;  //complement 
assign QHF = ~qhf;  //complement 
assign qja = ~QJA;  //complement 
assign qjb = ~QJB;  //complement 
assign QHO = ~qho;  //complement 
assign QHQ = ~qhq;  //complement 
assign QJD = ~qjd;  //complement 
assign QHL = ~qhl;  //complement 
assign QHN = ~qhn;  //complement 
assign EAC = ~eac;  //complement 
assign mao = ~MAO;  //complement 
assign map = ~MAP;  //complement 
assign EAB = ~eab;  //complement 
assign EAJ = ~eaj;  //complement 
assign EBJ = ~ebj;  //complement 
assign lab = ~LAB;  //complement 
assign laj = ~LAJ;  //complement 
assign oab = ~OAB;  //complement 
assign oeb = ~OEB;  //complement 
assign oej = ~OEJ;  //complement 
assign JAA = GAJ; 
assign jaa = ~JAA; //complement 
assign JAB = GAJ; 
assign jab = ~JAB;  //complement 
assign JAC = GAJ; 
assign jac = ~JAC;  //complement 
assign LFC = ~lfc;  //complement 
assign LFD = ~lfd;  //complement 
assign LGC = ~lgc;  //complement 
assign LGD = ~lgd;  //complement 
assign oaj = ~OAJ;  //complement 
assign oib = ~OIB;  //complement 
assign BAJ = ~baj;  //complement 
assign LBB = ~lbb;  //complement 
assign LCB = ~lcb;  //complement 
assign LDB = ~ldb;  //complement 
assign bab = ~BAB;  //complement 
assign LBJ = ~lbj;  //complement 
assign LCJ = ~lcj;  //complement 
assign LDJ = ~ldj;  //complement 
assign obb = ~OBB;  //complement 
assign ofb = ~OFB;  //complement 
assign ofj = ~OFJ;  //complement 
assign LEG = ~leg;  //complement 
assign LEH = ~leh;  //complement 
assign LEC = ~lec;  //complement 
assign obj = ~OBJ;  //complement 
assign LED = ~led;  //complement 
assign OLB = ~olb;  //complement 
assign OMB = ~omb;  //complement 
assign ONB = ~onb;  //complement 
assign QCA = ~qca;  //complement 
assign QFA = ~qfa;  //complement 
assign okb = ~OKB;  //complement 
assign ocb = ~OCB;  //complement 
assign ocj = ~OCJ;  //complement 
assign aab = ~AAB;  //complement 
assign aaj = ~AAJ;  //complement 
assign ogb = ~OGB;  //complement 
assign ogj = ~OGJ;  //complement 
assign tau =  qed & qeh & qfd  ; 
assign TAU = ~tau;  //complement 
assign tav =  qed & qeh & qfd  ; 
assign TAV = ~tav;  //complement 
assign BBB = ~bbb;  //complement 
assign BBJ = ~bbj;  //complement 
assign BCB = ~bcb;  //complement 
assign BDB = ~bdb;  //complement 
assign osb = ~OSB;  //complement 
assign tax =  qed & qeh & qfd  ; 
assign TAX = ~tax;  //complement 
assign taw =  qed & qeh & qfd  ; 
assign TAW = ~taw;  //complement 
assign QFB = ~qfb;  //complement 
assign QFC = ~qfc;  //complement 
assign QFD = ~qfd;  //complement 
assign BDJ = ~bdj;  //complement 
assign BEB = ~beb;  //complement 
assign odb = ~ODB;  //complement 
assign odj = ~ODJ;  //complement 
assign abb = ~ABB;  //complement 
assign abj = ~ABJ;  //complement 
assign ohb = ~OHB;  //complement 
assign ohj = ~OHJ;  //complement 
assign VCA = ~vca;  //complement 
assign vcc = ~VCC;  //complement 
assign vce = ~VCE;  //complement 
assign vcg = ~VCG;  //complement 
assign vch = ~VCH;  //complement 
assign vcd = ~VCD;  //complement 
assign vcf = ~VCF;  //complement 
assign vci = ~VCI;  //complement 
assign vcj = ~VCJ;  //complement 
assign mae = ~MAE;  //complement 
assign nac = ~NAC;  //complement 
assign nce = ~NCE;  //complement 
assign vcb = ~VCB;  //complement 
assign cca = ~CCA;  //complement 
assign ccb = ~CCB;  //complement 
assign ccc = ~CCC;  //complement 
assign dca = cca & ~( ZZI  ) | CCA & ( ZZI  );
assign DCA = ~dca ;
assign dcb = ccb & ~( cca & ZZI  ) | CCB & ( cca & ZZI  );
assign DCB = ~dcb ;  //complement 
assign dcc = ccc & ~( ccb & cca & ZZI  ) | CCC & ( ccb & cca & ZZI  );
assign DCC = ~dcc;  //complement;
assign DCG =  CCA & ccb & ccc & ccd & cce & ccf  ; 
assign dcg = ~DCG;  //complement  
assign ccd = ~CCD;  //complement 
assign cce = ~CCE;  //complement 
assign ccf = ~CCF;  //complement 
assign dcd = ccd & ~( ccc & ccb & cca  ) | CCD & ( ccc & ccb & cca  );
assign DCD = ~dcd ;
assign dce = cce & ~( ccd & ccc & ccb & cca  ) | CCE & ( ccd & ccc & ccb & cca  );
assign DCE = ~dce ;  //complement 
assign dcf = ccf & ~( cce & ccd & ccc & ccb & cca  ) | CCF & ( cce & ccd & ccc & ccb & cca  );
assign DCF = ~dcf;  //complement;
assign dch =  cca & ccb  |  CCC  |  CCD  |  CCE  |  CCF  ;
assign DCH = ~dch;  //complement 
assign nbc = ~NBC;  //complement 
assign nbk = ~NBK;  //complement 
assign gac = ~GAC;  //complement 
assign gak = ~GAK;  //complement 
assign FAC =  eap & ECO & ean & eam  ; 
assign fac = ~FAC;  //complement  
assign FBC =  eal & EAK & EAJ  ; 
assign fbc = ~FBC;  //complement 
assign vck = ~VCK;  //complement 
assign vcl = ~VCL;  //complement 
assign GBC = ~gbc;  //complement 
assign GBK = ~gbk;  //complement 
assign vcm = ~VCM;  //complement 
assign vcn = ~VCN;  //complement 
assign GCC = ~gcc;  //complement 
assign GCK = ~gck;  //complement 
assign FAK =  EBP & EBO & ebn & EBM  ; 
assign fak = ~FAK;  //complement  
assign FBK =  EBL & EBK  ; 
assign fbk = ~FBK;  //complement 
assign nag = ~NAG;  //complement 
assign nah = ~NAH;  //complement 
assign nai = ~NAI;  //complement 
assign naj = ~NAJ;  //complement 
assign nak = ~NAK;  //complement 
assign nal = ~NAL;  //complement 
assign nam = ~NAM;  //complement 
assign nan = ~NAN;  //complement 
assign QHP = ~qhp;  //complement 
assign QHC = ~qhc;  //complement 
assign qka = ~QKA;  //complement 
assign qkb = ~QKB;  //complement 
assign EAK = ~eak;  //complement 
assign EBK = ~ebk;  //complement 
assign lac = ~LAC;  //complement 
assign oac = ~OAC;  //complement 
assign oec = ~OEC;  //complement 
assign oek = ~OEK;  //complement 
assign LFE = ~lfe;  //complement 
assign LFF = ~lff;  //complement 
assign LGE = ~lge;  //complement 
assign LGF = ~lgf;  //complement 
assign LEE = ~lee;  //complement 
assign LEF = ~lef;  //complement 
assign LFG = ~lfg;  //complement 
assign LGG = ~lgg;  //complement 
assign oak = ~OAK;  //complement 
assign oic = ~OIC;  //complement 
assign BAK = ~bak;  //complement 
assign LBC = ~lbc;  //complement 
assign LCC = ~lcc;  //complement 
assign LDC = ~ldc;  //complement 
assign bac = ~BAC;  //complement 
assign LBK = ~lbk;  //complement 
assign LCK = ~lck;  //complement 
assign obc = ~OBC;  //complement 
assign ofc = ~OFC;  //complement 
assign ofk = ~OFK;  //complement 
assign QEB = ~qeb;  //complement 
assign QED = ~qed;  //complement 
assign QEK = ~qek;  //complement 
assign TAI = QEB; 
assign tai = ~TAI; //complement 
assign TAJ = QEB; 
assign taj = ~TAJ;  //complement 
assign TAQ = QED; 
assign taq = ~TAQ;  //complement 
assign TAR = QED; 
assign tar = ~TAR;  //complement 
assign obk = ~OBK;  //complement 
assign OLC = ~olc;  //complement 
assign OMC = ~omc;  //complement 
assign ONC = ~onc;  //complement 
assign QEA = ~qea;  //complement 
assign QEC = ~qec;  //complement 
assign THI = QEK; 
assign thi = ~THI; //complement 
assign THJ = QEK; 
assign thj = ~THJ;  //complement 
assign occ = ~OCC;  //complement 
assign ock = ~OCK;  //complement 
assign aac = ~AAC;  //complement 
assign aak = ~AAK;  //complement 
assign ogc = ~OGC;  //complement 
assign ogk = ~OGK;  //complement 
assign BBC = ~bbc;  //complement 
assign BBK = ~bbk;  //complement 
assign BCC = ~bcc;  //complement 
assign BDC = ~bdc;  //complement 
assign osc = ~OSC;  //complement 
assign BDK = ~bdk;  //complement 
assign BEC = ~bec;  //complement 
assign odc = ~ODC;  //complement 
assign odk = ~ODK;  //complement 
assign abc = ~ABC;  //complement 
assign abk = ~ABK;  //complement 
assign ohc = ~OHC;  //complement 
assign ohk = ~OHK;  //complement 
assign VDA = ~vda;  //complement 
assign vdc = ~VDC;  //complement 
assign vde = ~VDE;  //complement 
assign vdg = ~VDG;  //complement 
assign vdh = ~VDH;  //complement 
assign yya =  ZZO  ; 
assign YYA = ~yya;  //complement 
assign yym =  ZZO  ; 
assign YYM = ~yym;  //complement 
assign vdd = ~VDD;  //complement 
assign vdf = ~VDF;  //complement 
assign vdi = ~VDI;  //complement 
assign vdj = ~VDJ;  //complement 
assign jci =  yym  |  gbo  ; 
assign JCI = ~jci;  //complement 
assign jcj =  YYM  |  gbo  ; 
assign JCJ = ~jcj;  //complement 
assign cda = ~CDA;  //complement 
assign cdb = ~CDB;  //complement 
assign cdc = ~CDC;  //complement 
assign dda = cda & ~( ZZI  ) | CDA & ( ZZI  );
assign DDA = ~dda ;
assign ddb = cdb & ~( cda & ZZI  ) | CDB & ( cda & ZZI  );
assign DDB = ~ddb ;  //complement 
assign ddc = cdc & ~( cdb & cda & ZZI  ) | CDC & ( cdb & cda & ZZI  );
assign DDC = ~ddc;  //complement;
assign DDG =  CDA & cdb & cdc & cdd & cde & cdf  ; 
assign ddg = ~DDG;  //complement  
assign cdd = ~CDD;  //complement 
assign cde = ~CDE;  //complement 
assign cdf = ~CDF;  //complement 
assign ddd = cdd & ~( cdc & cdb & cda  ) | CDD & ( cdc & cdb & cda  );
assign DDD = ~ddd ;
assign dde = cde & ~( cdd & cdc & cdb & cda  ) | CDE & ( cdd & cdc & cdb & cda  );
assign DDE = ~dde ;  //complement 
assign ddf = cdf & ~( cde & cdd & cdc & cdb & cda  ) | CDF & ( cde & cdd & cdc & cdb & cda  );
assign DDF = ~ddf;  //complement;
assign ddh =  cda & cdb  |  CDC  |  CDD  |  CDE  |  CDF  ;
assign DDH = ~ddh;  //complement 
assign nbd = ~NBD;  //complement 
assign nbl = ~NBL;  //complement 
assign vdb = ~VDB;  //complement 
assign gad = ~GAD;  //complement 
assign FAD =  EAP & eao & EAN & EAM  ; 
assign fad = ~FAD;  //complement  
assign FBD =  eal & EAK & eaj  ; 
assign fbd = ~FBD;  //complement 
assign vdk = ~VDK;  //complement 
assign vdl = ~VDL;  //complement 
assign GBD = ~gbd;  //complement 
assign GBL = ~gbl;  //complement 
assign jcd =  gcl & gcd & gcb  ; 
assign JCD = ~jcd;  //complement 
assign vdm = ~VDM;  //complement 
assign vdn = ~VDN;  //complement 
assign GCD = ~gcd;  //complement 
assign GCL = ~gcl;  //complement 
assign FAL =  EBP & EBO & ebn & ebm  ; 
assign fal = ~FAL;  //complement  
assign FAM =  ebp & ebo & EBN & EBM  ; 
assign fam = ~FAM;  //complement 
assign mad = ~MAD;  //complement 
assign maf = ~MAF;  //complement 
assign nad = ~NAD;  //complement 
assign naf = ~NAF;  //complement 
assign ncd = ~NCD;  //complement 
assign ncf = ~NCF;  //complement 
assign QHR = ~qhr;  //complement 
assign QHS = ~qhs;  //complement 
assign QHD = ~qhd;  //complement 
assign qla = ~QLA;  //complement 
assign qlb = ~QLB;  //complement 
assign QKD = ~qkd;  //complement 
assign QLE = ~qle;  //complement 
assign FBL =  EBL  ; 
assign fbl = ~FBL;  //complement  
assign EAD = ~ead;  //complement 
assign EAL = ~eal;  //complement 
assign EBL = ~ebl;  //complement 
assign lad = ~LAD;  //complement 
assign lal = ~LAL;  //complement 
assign oad = ~OAD;  //complement 
assign oed = ~OED;  //complement 
assign oel = ~OEL;  //complement 
assign LFH = ~lfh;  //complement 
assign LGH = ~lgh;  //complement 
assign tae = qdd; 
assign TAE = ~tae; //complement 
assign taf = qdd; 
assign TAF = ~taf;  //complement 
assign TAK = QDE; 
assign tak = ~TAK;  //complement 
assign TAL = QDE; 
assign tal = ~TAL;  //complement 
assign oal = ~OAL;  //complement 
assign oid = ~OID;  //complement 
assign QDE = ~qde;  //complement 
assign BAL = ~bal;  //complement 
assign LBD = ~lbd;  //complement 
assign LCD = ~lcd;  //complement 
assign LDD = ~ldd;  //complement 
assign bad = ~BAD;  //complement 
assign LBL = ~lbl;  //complement 
assign LCL = ~lcl;  //complement 
assign LDL = ~ldl;  //complement 
assign obd = ~OBD;  //complement 
assign ofd = ~OFD;  //complement 
assign ofl = ~OFL;  //complement 
assign OUA = ~oua;  //complement 
assign OUC = ~ouc;  //complement 
assign TBA = QGC; 
assign tba = ~TBA; //complement 
assign tbc = qgc; 
assign TBC = ~tbc;  //complement 
assign TBI = QGC; 
assign tbi = ~TBI;  //complement 
assign tbk = qgc; 
assign TBK = ~tbk;  //complement 
assign obl = ~OBL;  //complement 
assign OLD = ~old;  //complement 
assign OMD = ~omd;  //complement 
assign OND = ~ond;  //complement 
assign QDA = ~qda;  //complement 
assign QGC = ~qgc;  //complement 
assign QDB = ~qdb;  //complement 
assign QDC = ~qdc;  //complement 
assign QDD = ~qdd;  //complement 
assign ocd = ~OCD;  //complement 
assign ocl = ~OCL;  //complement 
assign aad = ~AAD;  //complement 
assign aal = ~AAL;  //complement 
assign ogd = ~OGD;  //complement 
assign ogl = ~OGL;  //complement 
assign TAG = QDD; 
assign tag = ~TAG; //complement 
assign TAH = QDD; 
assign tah = ~TAH;  //complement 
assign osd = ~OSD;  //complement 
assign BDL = ~bdl;  //complement 
assign BED = ~bed;  //complement 
assign BBD = ~bbd;  //complement 
assign BBL = ~bbl;  //complement 
assign BCD = ~bcd;  //complement 
assign BDD = ~bdd;  //complement 
assign odd = ~ODD;  //complement 
assign odl = ~ODL;  //complement 
assign abd = ~ABD;  //complement 
assign abl = ~ABL;  //complement 
assign ohd = ~OHD;  //complement 
assign ohl = ~OHL;  //complement 
assign VEA = ~vea;  //complement 
assign vec = ~VEC;  //complement 
assign vee = ~VEE;  //complement 
assign veg = ~VEG;  //complement 
assign veh = ~VEH;  //complement 
assign ved = ~VED;  //complement 
assign vef = ~VEF;  //complement 
assign vei = ~VEI;  //complement 
assign vej = ~VEJ;  //complement 
assign nae = ~NAE;  //complement 
assign ncg = ~NCG;  //complement 
assign JGA = ~mbc & ~mbb & ~mba  ; 
assign JGB = ~mbc & ~mbb &  mba  ; 
assign JGC = ~mbc &  mbb & ~mba  ; 
assign JGD = ~mbc &  mbb &  mba  ; 
assign JGE =  mbc & ~mbb & ~mba  ; 
assign JGF =  mbc & ~mbb &  mba ; 
assign JGG =  mbc &  mbb & ~mba  ; 
assign JGH =  mbc &  mbb &  mba ; 
assign jgi = ZZI ; 
assign cea = ~CEA;  //complement 
assign ceb = ~CEB;  //complement 
assign cec = ~CEC;  //complement 
assign dea = cea & ~( ZZI  ) | CEA & ( ZZI  );
assign DEA = ~dea ;
assign deb = ceb & ~( cea & ZZI  ) | CEB & ( cea & ZZI  );
assign DEB = ~deb ;  //complement 
assign dec = cec & ~( ceb & cea & ZZI  ) | CEC & ( ceb & cea & ZZI  );
assign DEC = ~dec;  //complement;
assign DEG =  CEA & ceb & cec & ced & cee & cef  ; 
assign deg = ~DEG;  //complement  
assign ced = ~CED;  //complement 
assign cee = ~CEE;  //complement 
assign cef = ~CEF;  //complement 
assign ded = ced & ~( cec & ceb & cea  ) | CED & ( cec & ceb & cea  );
assign DED = ~ded ;
assign dee = cee & ~( ced & cec & ceb & cea  ) | CEE & ( ced & cec & ceb & cea  );
assign DEE = ~dee ;  //complement 
assign def = cef & ~( cee & ced & cec & ceb & cea  ) | CEF & ( cee & ced & cec & ceb & cea  );
assign DEF = ~def;  //complement;
assign okc = ~OKC;  //complement 
assign nbe = ~NBE;  //complement 
assign nbm = ~NBM;  //complement 
assign veb = ~VEB;  //complement 
assign gae = ~GAE;  //complement 
assign FAE =  EAP & ECO & ean & EAM  ; 
assign fae = ~FAE;  //complement  
assign FBE =  eal & EAK  ; 
assign fbe = ~FBE;  //complement 
assign vek = ~VEK;  //complement 
assign vel = ~VEL;  //complement 
assign GBE = ~gbe;  //complement 
assign JDB =  GCM & GCI  ; 
assign jdb = ~JDB;  //complement 
assign vem = ~VEM;  //complement 
assign ven = ~VEN;  //complement 
assign GCE = ~gce;  //complement 
assign GCM = ~gcm;  //complement 
assign FAN =  EBP & ebo & EBN & EBM  ; 
assign fan = ~FAN;  //complement  
assign FBM =  ebl  ; 
assign fbm = ~FBM;  //complement 
assign THO = QEF; 
assign tho = ~THO; //complement 
assign THP = QEF; 
assign thp = ~THP;  //complement 
assign THQ = QED; 
assign thq = ~THQ;  //complement 
assign THR = QED; 
assign thr = ~THR;  //complement 
assign mag = ~MAG;  //complement 
assign QHE = ~qhe;  //complement 
assign qsa = ~QSA;  //complement 
assign qsb = ~QSB;  //complement 
assign oke = ~OKE;  //complement 
assign EAE = ~eae;  //complement 
assign EAM = ~eam;  //complement 
assign EBM = ~ebm;  //complement 
assign ECM = ~ecm;  //complement 
assign lae = ~LAE;  //complement 
assign lam = ~LAM;  //complement 
assign oae = ~OAE;  //complement 
assign oee = ~OEE;  //complement 
assign oem = ~OEM;  //complement 
assign OLF = ~olf;  //complement 
assign OMF = ~omf;  //complement 
assign JFA = ~gai & ~gah & ~gag  ; 
assign JFB = ~gai & ~gah &  gag  ; 
assign JFC = ~gai &  gah & ~gag  ; 
assign JFD = ~gai &  gah &  gag  ; 
assign JFE =  gai & ~gah & ~gag  ; 
assign JFF =  gai & ~gah &  gag ; 
assign JFG =  gai &  gah & ~gag  ; 
assign JFH =  gai &  gah &  gag ; 
assign jfi = ZZI ; 
assign oam = ~OAM;  //complement 
assign oie = ~OIE;  //complement 
assign BAM = ~bam;  //complement 
assign LBE = ~lbe;  //complement 
assign LCE = ~lce;  //complement 
assign LDE = ~lde;  //complement 
assign bae = ~BAE;  //complement 
assign LBM = ~lbm;  //complement 
assign LCM = ~lcm;  //complement 
assign LDM = ~ldm;  //complement 
assign obe = ~OBE;  //complement 
assign ofe = ~OFE;  //complement 
assign ofm = ~OFM;  //complement 
assign QEF = ~qef;  //complement 
assign QEH = ~qeh;  //complement 
assign qqb = ~QQB;  //complement 
assign ONE = ~one;  //complement 
assign TAM = QEF; 
assign tam = ~TAM; //complement 
assign TAN = QEF; 
assign tan = ~TAN;  //complement 
assign TAO = QEF; 
assign tao = ~TAO;  //complement 
assign TAP = QEF; 
assign tap = ~TAP;  //complement 
assign obm = ~OBM;  //complement 
assign orc = ~ORC;  //complement 
assign ord = ~ORD;  //complement 
assign QEE = ~qee;  //complement 
assign QEG = ~qeg;  //complement 
assign OUB = ~oub;  //complement 
assign oce = ~OCE;  //complement 
assign ocm = ~OCM;  //complement 
assign aae = ~AAE;  //complement 
assign aam = ~AAM;  //complement 
assign oge = ~OGE;  //complement 
assign ogm = ~OGM;  //complement 
assign BDM = ~bdm;  //complement 
assign BEE = ~bee;  //complement 
assign BBE = ~bbe;  //complement 
assign BBM = ~bbm;  //complement 
assign BCE = ~bce;  //complement 
assign BDE = ~bde;  //complement 
assign ose = ~OSE;  //complement 
assign ode = ~ODE;  //complement 
assign odm = ~ODM;  //complement 
assign abe = ~ABE;  //complement 
assign abm = ~ABM;  //complement 
assign ohe = ~OHE;  //complement 
assign ohm = ~OHM;  //complement 
assign VFA = ~vfa;  //complement 
assign vfc = ~VFC;  //complement 
assign vfe = ~VFE;  //complement 
assign vfg = ~VFG;  //complement 
assign vfh = ~VFH;  //complement 
assign vfd = ~VFD;  //complement 
assign vff = ~VFF;  //complement 
assign vfi = ~VFI;  //complement 
assign vfj = ~VFJ;  //complement 
assign cfa = ~CFA;  //complement 
assign cfb = ~CFB;  //complement 
assign cfc = ~CFC;  //complement 
assign dfa = cfa & ~( ZZI  ) | CFA & ( ZZI  );
assign DFA = ~dfa ;
assign dfb = cfb & ~( cfa & ZZI  ) | CFB & ( cfa & ZZI  );
assign DFB = ~dfb ;  //complement 
assign dfc = cfc & ~( cfb & cfa & ZZI  ) | CFC & ( cfb & cfa & ZZI  );
assign DFC = ~dfc;  //complement;
assign DFG =  CFA & cfb & cfc & cfd & cfe & cff  ; 
assign dfg = ~DFG;  //complement  
assign cfd = ~CFD;  //complement 
assign cfe = ~CFE;  //complement 
assign cff = ~CFF;  //complement 
assign dfd = cfd & ~( cfc & cfb & cfa  ) | CFD & ( cfc & cfb & cfa  );
assign DFD = ~dfd ;
assign dfe = cfe & ~( cfd & cfc & cfb & cfa  ) | CFE & ( cfd & cfc & cfb & cfa  );
assign DFE = ~dfe ;  //complement 
assign dff = cff & ~( cfe & cfd & cfc & cfb & cfa  ) | CFF & ( cfe & cfd & cfc & cfb & cfa  );
assign DFF = ~dff;  //complement;
assign dfh =  cfa & cfb  |  CFC  |  CFD  |  CFE  |  CFF  ;
assign DFH = ~dfh;  //complement 
assign nbf = ~NBF;  //complement 
assign nbn = ~NBN;  //complement 
assign vfb = ~VFB;  //complement 
assign vgb = ~VGB;  //complement 
assign gaf = ~GAF;  //complement 
assign FBF =  eal & eak & EAJ  ; 
assign fbf = ~FBF;  //complement  
assign vfk = ~VFK;  //complement 
assign vfl = ~VFL;  //complement 
assign GBF = ~gbf;  //complement 
assign GBN = ~gbn;  //complement 
assign GDB = ~gdb;  //complement 
assign GDC = ~gdc;  //complement 
assign vfm = ~VFM;  //complement 
assign vfn = ~VFN;  //complement 
assign GCF = ~gcf;  //complement 
assign GCN = ~gcn;  //complement 
assign FAP =  ebp & EBO & ebn & ebm  ; 
assign fap = ~FAP;  //complement  
assign FBN =  ebl & EBK  ; 
assign fbn = ~FBN;  //complement 
assign QMA = ~qma;  //complement 
assign QMB = ~qmb;  //complement 
assign QMC = ~qmc;  //complement 
assign QPA = ~qpa;  //complement 
assign QPB = ~qpb;  //complement 
assign QOD = ~qod;  //complement 
assign qog = ~QOG;  //complement 
assign qoh = ~QOH;  //complement 
assign QTC = ~qtc;  //complement 
assign okf = ~OKF;  //complement 
assign EAF = ~eaf;  //complement 
assign EAN = ~ean;  //complement 
assign EBN = ~ebn;  //complement 
assign ECN = ~ecn;  //complement 
assign laf = ~LAF;  //complement 
assign lan = ~LAN;  //complement 
assign oaf = ~OAF;  //complement 
assign oef = ~OEF;  //complement 
assign oen = ~OEN;  //complement 
assign qof = ~QOF;  //complement 
assign JEA =  GCN & QRA & QAA  ; 
assign jea = ~JEA;  //complement 
assign JEB =  GCN & QRA & QAA  ; 
assign jeb = ~JEB;  //complement 
assign oan = ~OAN;  //complement 
assign oif = ~OIF;  //complement 
assign BAN = ~ban;  //complement 
assign LBF = ~lbf;  //complement 
assign LCF = ~lcf;  //complement 
assign LDF = ~ldf;  //complement 
assign baf = ~BAF;  //complement 
assign LBN = ~lbn;  //complement 
assign LDN = ~ldn;  //complement 
assign obf = ~OBF;  //complement 
assign off = ~OFF;  //complement 
assign ofn = ~OFN;  //complement 
assign qga = ~QGA;  //complement 
assign qoa = ~QOA;  //complement 
assign qob = ~QOB;  //complement 
assign obn = ~OBN;  //complement 
assign OJA = ~oja;  //complement 
assign OJB = ~ojb;  //complement 
assign OJL = ~ojl;  //complement 
assign ONF = ~onf;  //complement 
assign QEI = ~qei;  //complement 
assign QGE = ~qge;  //complement 
assign ora = ~ORA;  //complement 
assign orb = ~ORB;  //complement 
assign ocf = ~OCF;  //complement 
assign ocn = ~OCN;  //complement 
assign aaf = ~AAF;  //complement 
assign aan = ~AAN;  //complement 
assign ogf = ~OGF;  //complement 
assign ogn = ~OGN;  //complement 
assign LCN = ~lcn;  //complement 
assign QEJ = ~qej;  //complement 
assign qqa = ~QQA;  //complement 
assign TAS = QEJ; 
assign tas = ~TAS; //complement 
assign TAT = QEJ; 
assign tat = ~TAT;  //complement 
assign osf = ~OSF;  //complement 
assign BDN = ~bdn;  //complement 
assign BEF = ~bef;  //complement 
assign BBF = ~bbf;  //complement 
assign BBN = ~bbn;  //complement 
assign BCF = ~bcf;  //complement 
assign BDF = ~bdf;  //complement 
assign odf = ~ODF;  //complement 
assign odn = ~ODN;  //complement 
assign abf = ~ABF;  //complement 
assign abn = ~ABN;  //complement 
assign ohf = ~OHF;  //complement 
assign ohn = ~OHN;  //complement 
assign VGA = ~vga;  //complement 
assign vgc = ~VGC;  //complement 
assign vge = ~VGE;  //complement 
assign vgg = ~VGG;  //complement 
assign vgh = ~VGH;  //complement 
assign vgd = ~VGD;  //complement 
assign vgf = ~VGF;  //complement 
assign vgi = ~VGI;  //complement 
assign vgj = ~VGJ;  //complement 
assign mba = ~MBA;  //complement 
assign nbg = ~NBG;  //complement 
assign nbo = ~NBO;  //complement 
assign gag = ~GAG;  //complement 
assign FAF =  ecp & ECO & ecn & ECM  ; 
assign faf = ~FAF;  //complement  
assign FAG =  EAP & EAO & EAN & eam  ; 
assign fag = ~FAG;  //complement 
assign vgk = ~VGK;  //complement 
assign vgl = ~VGL;  //complement 
assign GBG = ~gbg;  //complement 
assign GBO = ~gbo;  //complement 
assign GCH = ~gch;  //complement 
assign GCP = ~gcp;  //complement 
assign vgm = ~VGM;  //complement 
assign vgn = ~VGN;  //complement 
assign GCO = ~gco;  //complement 
assign FBO =  ebl & ebk  ; 
assign fbo = ~FBO;  //complement 
assign jda =  gcf & gch & gcm  ; 
assign JDA = ~jda;  //complement 
assign QPC = ~qpc;  //complement 
assign TGK = QBB; 
assign tgk = ~TGK; //complement 
assign qld = ~QLD;  //complement 
assign qua = ~QUA;  //complement 
assign qva = ~QVA;  //complement 
assign EAG = ~eag;  //complement 
assign EAO = ~eao;  //complement 
assign EBO = ~ebo;  //complement 
assign ECO = ~eco;  //complement 
assign lag = ~LAG;  //complement 
assign lao = ~LAO;  //complement 
assign oag = ~OAG;  //complement 
assign oeg = ~OEG;  //complement 
assign oeo = ~OEO;  //complement 
assign the = qdd; 
assign THE = ~the; //complement 
assign thf = qdd; 
assign THF = ~thf;  //complement 
assign THG = QDD; 
assign thg = ~THG;  //complement 
assign THH = QDD; 
assign thh = ~THH;  //complement 
assign ojj = ~OJJ;  //complement 
assign ojk = ~OJK;  //complement 
assign oao = ~OAO;  //complement 
assign oig = ~OIG;  //complement 
assign LBG = ~lbg;  //complement 
assign LCG = ~lcg;  //complement 
assign LDG = ~ldg;  //complement 
assign LBO = ~lbo;  //complement 
assign LCO = ~lco;  //complement 
assign LDO = ~ldo;  //complement 
assign obg = ~OBG;  //complement 
assign ofg = ~OFG;  //complement 
assign ofo = ~OFO;  //complement 
assign TGA = QBA; 
assign tga = ~TGA; //complement 
assign TGB = QBA; 
assign tgb = ~TGB;  //complement 
assign TGC = QBA; 
assign tgc = ~TGC;  //complement 
assign TGD = QBA; 
assign tgd = ~TGD;  //complement 
assign TGE = QBA; 
assign tge = ~TGE; //complement 
assign TGF = QBA; 
assign tgf = ~TGF;  //complement 
assign obo = ~OBO;  //complement 
assign ojf = ~OJF;  //complement 
assign ojg = ~OJG;  //complement 
assign ojh = ~OJH;  //complement 
assign oji = ~OJI;  //complement 
assign TGG = QBB; 
assign tgg = ~TGG; //complement 
assign TGH = QBB; 
assign tgh = ~TGH;  //complement 
assign TGI = QBB; 
assign tgi = ~TGI;  //complement 
assign TGJ = QBB; 
assign tgj = ~TGJ;  //complement 
assign qba = ~QBA;  //complement 
assign qbb = ~QBB;  //complement 
assign tgl = ~TGL;  //complement 
assign ocg = ~OCG;  //complement 
assign oco = ~OCO;  //complement 
assign aag = ~AAG;  //complement 
assign aao = ~AAO;  //complement 
assign ogg = ~OGG;  //complement 
assign ogo = ~OGO;  //complement 
assign okd = ~OKD;  //complement 
assign BBG = ~bbg;  //complement 
assign BBO = ~bbo;  //complement 
assign BCG = ~bcg;  //complement 
assign BDG = ~bdg;  //complement 
assign osg = ~OSG;  //complement 
assign BDO = ~bdo;  //complement 
assign BEG = ~beg;  //complement 
assign odg = ~ODG;  //complement 
assign odo = ~ODO;  //complement 
assign abg = ~ABG;  //complement 
assign abo = ~ABO;  //complement 
assign ohg = ~OHG;  //complement 
assign oho = ~OHO;  //complement 
assign THS = QEJ; 
assign ths = ~THS; //complement 
assign THT = QEJ; 
assign tht = ~THT;  //complement 
assign VHA = ~vha;  //complement 
assign vhc = ~VHC;  //complement 
assign vhe = ~VHE;  //complement 
assign vhg = ~VHG;  //complement 
assign vhh = ~VHH;  //complement 
assign vhd = ~VHD;  //complement 
assign vhf = ~VHF;  //complement 
assign vhi = ~VHI;  //complement 
assign vhj = ~VHJ;  //complement 
assign mbb = ~MBB;  //complement 
assign nbh = ~NBH;  //complement 
assign nbp = ~NBP;  //complement 
assign vhb = ~VHB;  //complement 
assign gah = ~GAH;  //complement 
assign FAH =  eap & EAO & EAN & EAM  ; 
assign fah = ~FAH;  //complement  
assign FBH =  EAL & eak & eaj  ; 
assign fbh = ~FBH;  //complement 
assign vhk = ~VHK;  //complement 
assign vhl = ~VHL;  //complement 
assign GBH = ~gbh;  //complement 
assign jdc =  gco & gcf & gch  ; 
assign JDC = ~jdc;  //complement 
assign vhm = ~VHM;  //complement 
assign vhn = ~VHN;  //complement 
assign FBP =  EBJ  ; 
assign fbp = ~FBP;  //complement  
assign QVB = ~qvb;  //complement 
assign QVD = ~qvd;  //complement 
assign QVF = ~qvf;  //complement 
assign QVH = ~qvh;  //complement 
assign QPE = ~qpe;  //complement 
assign QPF = ~qpf;  //complement 
assign TCA = QAD & GDA ; 
assign tca = ~TCA ; //complement 
assign TCB = QAD & GDA ; 
assign tcb = ~TCB ;  //complement 
assign QVC = ~qvc;  //complement 
assign QVE = ~qve;  //complement 
assign QVG = ~qvg;  //complement 
assign QVI = ~qvi;  //complement 
assign QVJ = ~qvj;  //complement 
assign QVK = ~qvk;  //complement 
assign bbh = aap; 
assign BBH = ~bbh; //complement 
assign bbp = abh; 
assign BBP = ~bbp;  //complement 
assign bch = abp; 
assign BCH = ~bch;  //complement 
assign bdh = bbp; 
assign BDH = ~bdh;  //complement 
assign TXE = ~txe;  //complement 
assign TXF = ~txf;  //complement 
assign TXG = ~txg;  //complement 
assign TXH = ~txh;  //complement 
assign EAH = ~eah;  //complement 
assign EAP = ~eap;  //complement 
assign EBP = ~ebp;  //complement 
assign ECP = ~ecp;  //complement 
assign lah = ~LAH;  //complement 
assign lap = ~LAP;  //complement 
assign oah = ~OAH;  //complement 
assign oeh = ~OEH;  //complement 
assign oep = ~OEP;  //complement 
assign tka = ~TKA;  //complement 
assign tkb = ~TKB;  //complement 
assign tkc = ~TKC;  //complement 
assign tkd = ~TKD;  //complement 
assign oih = ~OIH;  //complement 
assign oap = ~OAP;  //complement 
assign OJC = ~ojc;  //complement 
assign OJD = ~ojd;  //complement 
assign OJE = ~oje;  //complement 
assign QCE = ~qce;  //complement 
assign TDA = QAD & qra ; 
assign tda = ~TDA ; //complement 
assign TDB = QAD & qra ; 
assign tdb = ~TDB ;  //complement 
assign TEA = QAD & QRA ; 
assign tea = ~TEA ;  //complement 
assign TEB = QAD & QRA; 
assign teb = ~TEB; 
assign LBP = ~lbp;  //complement 
assign LCP = ~lcp;  //complement 
assign LDP = ~ldp;  //complement 
assign qra = ~QRA;  //complement 
assign obh = ~OBH;  //complement 
assign ofh = ~OFH;  //complement 
assign ofp = ~OFP;  //complement 
assign LBH = ~lbh;  //complement 
assign LCH = ~lch;  //complement 
assign LDH = ~ldh;  //complement 
assign qnb = ~QNB;  //complement 
assign qnd = ~QND;  //complement 
assign qne = ~QNE;  //complement 
assign qnf = ~QNF;  //complement 
assign obp = ~OBP;  //complement 
assign OTA = ~ota;  //complement 
assign QNA = ~qna;  //complement 
assign QNC = ~qnc;  //complement 
assign qaa = ~QAA;  //complement 
assign qab = ~QAB;  //complement 
assign qac = ~QAC;  //complement 
assign qad = ~QAD;  //complement 
assign och = ~OCH;  //complement 
assign ocp = ~OCP;  //complement 
assign aah = ~AAH;  //complement 
assign aap = ~AAP;  //complement 
assign ogh = ~OGH;  //complement 
assign ogp = ~OGP;  //complement 
assign taa = qcd; 
assign TAA = ~taa; //complement 
assign tab = qcd; 
assign TAB = ~tab;  //complement 
assign tac = qcd; 
assign TAC = ~tac;  //complement 
assign tad = qcd; 
assign TAD = ~tad;  //complement 
assign jbe = abp & QCE ; 
assign JBE = ~jbe ; //complement 
assign jbf = abp & QCE ; 
assign JBF = ~jbf ;  //complement 
assign jbg = abp & QCE ; 
assign JBG = ~jbg ;  //complement 
assign jbh = abp & QCE; 
assign JBH = ~jbh; 
assign THA = QCE; 
assign tha = ~THA; //complement 
assign THB = QCE; 
assign thb = ~THB;  //complement 
assign THC = QCE; 
assign thc = ~THC;  //complement 
assign THD = QCE; 
assign thd = ~THD;  //complement 
assign QCB = ~qcb;  //complement 
assign QCC = ~qcc;  //complement 
assign QCD = ~qcd;  //complement 
assign jba = abp & QCD ; 
assign JBA = ~jba ; //complement 
assign jbb = abp & QCD ; 
assign JBB = ~jbb ;  //complement 
assign jbc = abp & QCD ; 
assign JBC = ~jbc ;  //complement 
assign jbd = abp & QCD; 
assign JBD = ~jbd; 
assign odh = ~ODH;  //complement 
assign odp = ~ODP;  //complement 
assign abh = ~ABH;  //complement 
assign abp = ~ABP;  //complement 
assign ohh = ~OHH;  //complement 
assign ohp = ~OHP;  //complement 
assign TXA = ~txa;  //complement 
assign TXB = ~txb;  //complement 
assign TXC = ~txc;  //complement 
assign TXD = ~txd;  //complement 
assign BDP = ~bdp;  //complement 
assign BEH = ~beh;  //complement 
assign QUB = ~qub;  //complement 
assign QUC = ~quc;  //complement 
assign osh = ~OSH;  //complement 
assign iaa = ~IAA; //complement 
assign iab = ~IAB; //complement 
assign iac = ~IAC; //complement 
assign iad = ~IAD; //complement 
assign iae = ~IAE; //complement 
assign iaf = ~IAF; //complement 
assign iag = ~IAG; //complement 
assign iah = ~IAH; //complement 
assign iai = ~IAI; //complement 
assign iaj = ~IAJ; //complement 
assign iak = ~IAK; //complement 
assign ial = ~IAL; //complement 
assign iam = ~IAM; //complement 
assign ian = ~IAN; //complement 
assign iao = ~IAO; //complement 
assign iap = ~IAP; //complement 
assign iba = ~IBA; //complement 
assign ibb = ~IBB; //complement 
assign ibc = ~IBC; //complement 
assign ibd = ~IBD; //complement 
assign ibe = ~IBE; //complement 
assign ibf = ~IBF; //complement 
assign ibg = ~IBG; //complement 
assign ibh = ~IBH; //complement 
assign ibi = ~IBI; //complement 
assign ibj = ~IBJ; //complement 
assign ibk = ~IBK; //complement 
assign ibl = ~IBL; //complement 
assign ibm = ~IBM; //complement 
assign ibn = ~IBN; //complement 
assign ibo = ~IBO; //complement 
assign ibp = ~IBP; //complement 
assign ica = ~ICA; //complement 
assign icb = ~ICB; //complement 
assign icc = ~ICC; //complement 
assign icd = ~ICD; //complement 
assign ice = ~ICE; //complement 
assign icf = ~ICF; //complement 
assign icg = ~ICG; //complement 
assign ich = ~ICH; //complement 
assign ici = ~ICI; //complement 
assign icj = ~ICJ; //complement 
assign ick = ~ICK; //complement 
assign icl = ~ICL; //complement 
assign icm = ~ICM; //complement 
assign icn = ~ICN; //complement 
assign ico = ~ICO; //complement 
assign icp = ~ICP; //complement 
assign ida = ~IDA; //complement 
assign idb = ~IDB; //complement 
assign idc = ~IDC; //complement 
assign idd = ~IDD; //complement 
assign ide = ~IDE; //complement 
assign idf = ~IDF; //complement 
assign iea = ~IEA; //complement 
assign ieb = ~IEB; //complement 
assign ifa = ~IFA; //complement 
assign iga = ~IGA; //complement 
assign iha = ~IHA; //complement 
assign ihb = ~IHB; //complement 
assign ihf = ~IHF; //complement 
assign ija = ~IJA; //complement 
assign ika = ~IKA; //complement 
assign ikb = ~IKB; //complement 
assign ikc = ~IKC; //complement 
assign ikd = ~IKD; //complement 
assign ike = ~IKE; //complement 
assign ikf = ~IKF; //complement 
assign ikg = ~IKG; //complement 
assign ikh = ~IKH; //complement 
assign ila = ~ILA; //complement 
always@(posedge IZZ )
   begin 
 vaa <=  naa  |  nba  ; 
 VAC <=  NAC & NBA  |  VAB  ; 
 VAE <=  NAE & NBA  |  VAD  ; 
 VAG <=  NAG & NBA  |  VAF  ; 
 VAH <=  NAH & NBA  |  VAG  ; 
 VAD <=  NAD & NBA  |  VAC  ; 
 VAF <=  NAF & NBA  |  VAE  ; 
 VAI <=  NAI & NBA  |  VAH  ; 
 VAJ <=  NAJ & NBA  |  VAI  ; 
 MAA <= QHA ; 
 MBC <= GAI ; 
 NAA <= MAA ; 
 CAA <= DAA & QIB |  BAA & qib ; 
 CAB <= DAB & QIB |  BAB & qib ; 
 CAC <= DAC & QIB |  BAC & qib ; 
 CAD <= DAD & QIB |  BAD & qib ; 
 CAE <= DAE & QIB |  BAE & qib ; 
 CAF <= DAF & QIB |  BAF & qib ; 
 NBA <= JGA ; 
 NBI <= JGA ; 
 NCA <= MAA ; 
 VAB <= VAA ; 
 GAA <=  EAA & TGG  |  GAA & tgg  ; 
 GAI <=  EAI & TGG  |  GAI & tgg  ; 
 VAK <=  NAK & NBI  |  VAJ  ; 
 VAL <=  NAL & NBI  |  VAK  ; 
 gba <=  faa & TGB  |  fbi & TGC  |  gba & tgh  ; 
 gda <=  faa & fab & TGI  |  fbi & TGL  |  gda & tgl  ; 
 VAM <=  NAM & NBI  |  VAL  ; 
 VAN <=  NAN & NBI  |  VAM  ; 
 gca <=  fai & TGD  |  FBI & TGE  |  gca & tgi  ; 
 gci <=  ZZO & TGD  |  fbp & TGE  |  gci & tgi  ; 
 qha <=  jci  |  tda  ; 
 QIA <=  QIA & dag  |  GCN & QAB  ; 
 QIB <=  QIA & dag  |  GCN & QAB  ; 
 qid <=  dah  |  qia  ; 
 OKA <=  DAH & qid & QIA  |  QTB  ; 
 eaa <= ica ; 
 eai <= ici ; 
 LAA <=  ICA & tca  |  GAA & TCA  ; 
 LAI <=  ICI & tca  |  JAB & TCA  ; 
 OAA <=  AAA & TAA  |  ICA & TAE  |  LBA & TAI  |  LAA & TAM  ; 
 OEA <=  ICA & TBA  |  LAA & TBB  |  LGA & TKA  ; 
 OEI <=  ICI & TBA  |  LAI & TBB  |  LFA & TKA  ; 
 lea <= ika ; 
 leb <= ikb ; 
 lfa <= lea ; 
 lfb <= leb ; 
 lga <= lfa ; 
 lgb <= lfb ; 
 OAI <=  AAI & TAB  |  ICI & TAF  |  LBI & TAJ  |  LAI & TAN  ; 
 OIA <=  VAN  |  NBI & MAO  |  JFA & JEA  ; 
 bai <= ida ; 
 lba <= laa ; 
 lca <= lba ; 
 lda <= lca ; 
 BAA <= IDA ; 
 lbi <= lai ; 
 lci <= lbi ; 
 ldi <= lci ; 
 OBA <=  ABA & TAC  |  LAA & TAK  |  IBA & TAO  |  TAQ  ; 
 OFA <=  LAA & TBC  |  LEA & TKC  |  TBD  ; 
 OFI <=  LAI & TBC  |  IKA & TKC  |  TBD  ; 
 OBI <=  ABI & TAD  |  LAI & TAL  |  LBI & TAP  |  TAR  ; 
 ola <= qia ; 
 oma <= qia ; 
 ona <= baa ; 
 qgb <=  gba  |  qaa  ; 
 qgd <=  gba  |  qaa  |  gaj  ; 
 QTA <= IHA ; 
 QTB <= IHA ; 
 OCA <=  LCA & TAG  |  LAA & TAS  |  JBE & TAW  ; 
 OCI <=  LCI & TAG  |  LAI & TAS  |  JBG & TAW  ; 
 AAA <= IAA ; 
 AAI <= IAI ; 
 OGA <= IAA ; 
 OGI <= IAI ; 
 bba <= aai ; 
 bbi <= aba ; 
 bca <= abi ; 
 bda <= bbi ; 
 OSA <=  TXA & AAA  |  TXB & BBA  |  TXC & BDA  |  TXD & BEA  ; 
 bdi <= bca ; 
 bea <= bdi ; 
 ODA <=  LDA & TAH  |  LBA & TAT  |  JBA & TAX  ; 
 ODI <=  LDI & TAH  |  LBI & TAT  |  JBC & TAX  ; 
 ABA <= IBA ; 
 ABI <= IBI ; 
 OHA <= IBA ; 
 OHI <= IBI ; 
 vba <=  naa  |  nbb  ; 
 VBC <=  NAC & NBB  |  VBB  ; 
 VBE <=  NAE & NBB  |  VBD  ; 
 VBG <=  NAG & NBB  |  VBF  ; 
 VBH <=  NAH & NBB  |  VBG  ; 
 VBD <=  NAD & NBB  |  VBC  ; 
 VBF <=  NAF & NBB  |  VBE  ; 
 VBI <=  NAI & NBB  |  VBH  ; 
 VBJ <=  NAJ & NBB  |  VBI  ; 
 MAC <= QHB ; 
 MAH <= QHF ; 
 NCC <= MAC ; 
 qsd <=  dfh  |  qsd  ; 
 CBA <= DBA & QJB |  BAA & qjb ; 
 CBB <= DBB & QJB |  BAB & qjb ; 
 CBC <= DBC & QJB |  BAC & qjb ; 
 CBD <= DBD & QJB |  BAD & qjb ; 
 CBE <= DBE & QJB |  BAE & qjb ; 
 CBF <= DBF & QJB |  BAF & qjb ; 
 MAI <= QHG ; 
 MAJ <= QHH ; 
 MAK <= QHI ; 
 MAL <= QHJ ; 
 NCI <= MAI ; 
 NCJ <= MAJ ; 
 NCK <= MAK ; 
 NCL <= MAL ; 
 MAM <=  QHK  |  QHL  ; 
 NCM <= MAM ; 
 NCN <=  MAN  |  QHO  ; 
 MAN <=  QHM  |  QHN  ; 
 NBB <= JGB ; 
 NBJ <= JGB ; 
 NCH <= MAH ; 
 VBB <= VBA ; 
 LAK <=  ICK & tca  |  JAB & TCA  ; 
 GAB <=  EAB & TGG  |  GAB & tgg  ; 
 GAJ <=  EAJ & TGG  |  GAJ & tgg  ; 
 VBK <=  NAK & NBJ  |  VBJ  ; 
 VBL <=  NAL & NBJ  |  VBK  ; 
 gbb <=  fad & TGB  |  fba & TGC  |  gbb & tgh  ; 
 VBM <=  NAM & NBJ  |  VBL  ; 
 VBN <=  NAN & NBJ  |  VBM  ; 
 ldk <= lck ; 
 gcb <=  faj & TGD  |  fbm & TGE  |  gcb & tgi  ; 
 gcj <=  fak & TGD  |  fbm & TGE  |  gcj & tgi  ; 
 qhi <=  jcb  |  tdb  ; 
 qhj <=  jcg  |  tdb  ; 
 qhk <=  jca  |  tdb  ; 
 qhm <=  gcd  |  tdb  ; 
 qhg <=  jcf  |  tea  ; 
 qhh <=  jch  |  tea  ; 
 qhb <=  jci  |  tea  ; 
 qhf <=  jch  |  tda  ; 
 QJA <=  QJA & dbg  |  JCD & QAB  ; 
 QJB <=  QJA & dbg  |  JCD & QAB  ; 
 qho <=  jca  |  teb  ; 
 qhq <=  gcd  |  teb  ; 
 qjd <=  dbh  |  qia  ; 
 qhl <=  jcb  |  tdb  ; 
 qhn <=  jcg  |  tdb  ; 
 eac <= icc ; 
 MAO <=  QHP  |  QHQ  ; 
 MAP <=  QHP  |  QHQ  ; 
 eab <= icb ; 
 eaj <= icj ; 
 ebj <= icj ; 
 LAB <=  ICB & tca  |  GAB & TCA  ; 
 LAJ <=  ICJ & tca  |  JAB & TCA  ; 
 OAB <=  AAB & TAA  |  ICB & TAE  |  LBB & TAI  |  LAB & TAM  ; 
 OEB <=  ICB & TBA  |  LAB & TBB  |  LGB & TKA  ; 
 OEJ <=  ICJ & TBA  |  LAJ & TBB  |  LFB & TKA  ; 
 lfc <= lec ; 
 lfd <= led ; 
 lgc <= lfc ; 
 lgd <= lfd ; 
 OAJ <=  AAJ & TAB  |  ICJ & TAF  |  LBJ & TAJ  |  LAJ & TAN  ; 
 OIB <=  VBN  |  NBJ & MAO  |  JFB & JEA  ; 
 baj <= idb ; 
 lbb <= lab ; 
 lcb <= lbb ; 
 ldb <= lcb ; 
 BAB <= IDB ; 
 lbj <= laj ; 
 lcj <= lbj ; 
 ldj <= lcj ; 
 OBB <=  ABB & TAC  |  LAB & TAK  |  IBB & TAO  |  TAQ  ; 
 OFB <=  LAB & TBC  |  LEB & TKC  |  TBD  ; 
 OFJ <=  LAJ & TBC  |  IKB & TKC  |  TBD  ; 
 leg <= ikg ; 
 leh <= ikh ; 
 lec <= ikc ; 
 OBJ <=  ABJ & TAD  |  LAJ & TAL  |  LBJ & TAP  |  TAR  ; 
 led <= ikd ; 
 olb <= qja ; 
 omb <= qja ; 
 onb <= bab ; 
 qca <=  gbb  |  qaa  ; 
 qfa <=  gbb  |  qaa  |  gaj  ; 
 OKB <=  DBH & qjd & QJA  |  IJA  |  QTB  ; 
 OCB <=  LCB & TAG  |  LAB & TAS  |  JBE & TAW  ; 
 OCJ <=  LCJ & TAG  |  LAJ & TAS  |  JBG & TAW  ; 
 AAB <= IAB ; 
 AAJ <= IAJ ; 
 OGB <= IAB ; 
 OGJ <= IAJ ; 
 bbb <= aaj ; 
 bbj <= abb ; 
 bcb <= abj ; 
 bdb <= bbj ; 
 OSB <=  TXA & AAB  |  TXB & BBB  |  TXC & BDB  |  TXD & BEB  ; 
 qfb <= qfa ; 
 qfc <= qfb ; 
 qfd <= qfc ; 
 bdj <= bcb ; 
 beb <= bdj ; 
 ODB <=  LDB & TAH  |  LBB & TAT  |  JBA & TAX  ; 
 ODJ <=  LDJ & TAH  |  LBJ & TAT  |  JBC & TAX  ; 
 ABB <= IBB ; 
 ABJ <= IBJ ; 
 OHB <= IBB ; 
 OHJ <= IBJ ; 
 vca <=  naa  |  nbc  ; 
 VCC <=  NAC & NBC  |  VCB  ; 
 VCE <=  NAE & NBC  |  VCD  ; 
 VCG <=  NAG & NBC  |  VCF  ; 
 VCH <=  NAH & NBC  |  VCG  ; 
 VCD <=  NAD & NBC  |  VCC  ; 
 VCF <=  NAF & NBC  |  VCE  ; 
 VCI <=  NAI & NBC  |  VCH  ; 
 VCJ <=  NAJ & NBC  |  VCI  ; 
 MAE <= QHC ; 
 NAC <= MAC ; 
 NCE <= MAE ; 
 VCB <= VCA ; 
 CCA <= DCA & QKB |  BAA & qkb ; 
 CCB <= DCB & QKB |  BAB & qkb ; 
 CCC <= DCC & QKB |  BAC & qkb ; 
 CCD <= DCD & QKB |  BAD & qkb ; 
 CCE <= DCE & QKB |  BAE & qkb ; 
 CCF <= DCF & QKB |  BAF & qkb ; 
 NBC <= JGC ; 
 NBK <= JGC ; 
 GAC <=  EAC & TGG  |  GAC & tgg  ; 
 GAK <=  EAK & TGG  |  GAK & tgg  ; 
 VCK <=  NAK & NBK  |  VCJ  ; 
 VCL <=  NAL & NBK  |  VCK  ; 
 gbc <=  fab & TGB  |  fbb & TGC  |  gbc & tgh  ; 
 gbk <=  fae & TGB  |  fbl & TGC  |  gbk & tgh  ; 
 VCM <=  NAM & NBK  |  VCL  ; 
 VCN <=  NAN & NBK  |  VCM  ; 
 gcc <=  fai & TGD  |  fbk & TGE  |  gcc & tgi  ; 
 gck <=  fan & TGD  |  fbn & TGE  |  gck & tgi  ; 
 NAG <= MAG ; 
 NAH <= MAH ; 
 NAI <= MAI ; 
 NAJ <= MAJ ; 
 NAK <= MAK ; 
 NAL <= MAL ; 
 NAM <= MAM ; 
 NAN <=  MAN  |  QHO  ; 
 qhp <=  gcn  |  tdb  ; 
 qhc <=  jcc  |  tda  ; 
 QKA <=  QKA & dcg  |  GCA & QAB  ; 
 QKB <=  QKA & dcg  |  GCA & QAB  ; 
 eak <= ick ; 
 ebk <= ick ; 
 LAC <=  ICC & tca  |  GAC & TCA  ; 
 OAC <=  AAC & TAA  |  ICC & TAE  |  LBC & TAI  |  LAC & TAM  ; 
 OEC <=  ICC & TBA  |  LAC & TBB  |  LGC & TKA  ; 
 OEK <=  ICK & TBA  |  LAK & TBB  |  LFC & TKA  ; 
 lfe <= lee ; 
 lff <= lef ; 
 lge <= lfe ; 
 lgf <= lff ; 
 lee <= ike ; 
 lef <= ikf ; 
 lfg <= leg ; 
 lgg <= lfg ; 
 OAK <=  AAK & TAB  |  ICK & TAF  |  LBK & TAJ  |  LAK & TAN  ; 
 OIC <=  VCN  |  NBK & MAO  |  JFC & JEA  ; 
 bak <= idc ; 
 lbc <= lac ; 
 lcc <= lbc ; 
 ldc <= lcc ; 
 BAC <= IDC ; 
 lbk <= lak ; 
 lck <= lbk ; 
 OBC <=  ABC & TAC  |  LAC & TAK  |  LBC & TAO  |  TAQ  ; 
 OFC <=  LAC & TBC  |  LEC & TKC  |  TBD  ; 
 OFK <=  LAK & TBC  |  IKC & TKC  |  TBD  ; 
 qeb <= qea ; 
 qed <= qec ; 
 qek <= qea ; 
 OBK <=  ABK & TAD  |  LAK & TAL  |  LBK & TAP  |  TAR  ; 
 olc <= qka ; 
 omc <= qka ; 
 onc <= bac ; 
 qea <=  gbc  |  qaa  ; 
 qec <=  gbc  |  qaa  |  gaj  ; 
 OCC <=  LCC & TAG  |  LAC & TAS  |  JBE & TAW  ; 
 OCK <=  LCK & TAG  |  LAK & TAS  |  JBG & TAW  ; 
 AAC <= IAC ; 
 AAK <= IAK ; 
 OGC <= IAC ; 
 OGK <= IAK ; 
 bbc <= aak ; 
 bbk <= abc ; 
 bcc <= abk ; 
 bdc <= bbk ; 
 OSC <=  TXA & AAC  |  TXB & BBC  |  TXC & BDC  |  TXD & BEC  ; 
 bdk <= bcc ; 
 bec <= bdk ; 
 ODC <=  LDC & TAH  |  LBC & TAT  |  JBA & TAX  ; 
 ODK <=  LDK & TAH  |  LBK & TAT  |  JBC & TAX  ; 
 ABC <= IBC ; 
 ABK <= IBK ; 
 OHC <= IBC ; 
 OHK <= IBK ; 
 vda <=  naa  |  nbd  ; 
 VDC <=  NAC & NBA  |  VDB  ; 
 VDE <=  NAE & NBA  |  VDD  ; 
 VDG <=  NAG & NBA  |  VDF  ; 
 VDH <=  NAH & NBA  |  VDG  ; 
 VDD <=  NAD & NBA  |  VDC  ; 
 VDF <=  NAF & NBA  |  VDE  ; 
 VDI <=  NAI & NBA  |  VDH  ; 
 VDJ <=  NAJ & NBA  |  VDI  ; 
 CDA <= DDA & QLB |  BAI & qlb ; 
 CDB <= DDB & QLB |  BAJ & qlb ; 
 CDC <= DDC & QLB |  BAK & qlb ; 
 CDD <= DDD & QLB |  BAL & qlb ; 
 CDE <= DDE & QLB |  BAM & qlb ; 
 CDF <= DDF & QLB |  BAN & qlb ; 
 NBD <= JGD ; 
 NBL <= JGD ; 
 VDB <= VDA ; 
 GAD <=  EAD & TGG  |  GAD & tgg  ; 
 VDK <=  NAK & NBL  |  VDJ  ; 
 VDL <=  NAL & NBL  |  VDK  ; 
 gbd <=  faf & TGB  |  fbc & TGC  |  gbd & tgh  ; 
 gbl <=  fac & TGB  |  fbe & TGC  |  gbl & tgh  ; 
 VDM <=  NAM & NBL  |  VDL  ; 
 VDN <=  NAN & NBL  |  VDM  ; 
 gcd <=  fal & TGD  |  fbk & TGE  |  gcd & tgi  ; 
 gcl <=  fam & TGD  |  fbm & TGE  |  gcl & tgi  ; 
 MAD <= QHR ; 
 MAF <= QHS ; 
 NAD <= MAD ; 
 NAF <= MAF ; 
 NCD <= MAD ; 
 NCF <= MAF ; 
 qhr <=  jcj  |  tdb  ; 
 qhs <=  jcj  |  teb  ; 
 qhd <=  jcf  |  tda  ; 
 QLA <=  QLA & ddg  |  GBK & QAB  |  QMC  ; 
 QLB <=  QLA & ddg  |  GBK & QAB  |  QMC  ; 
 qkd <=  dch  |  qka  ; 
 qle <=  ddh  |  qla  ; 
 ead <= icd ; 
 eal <= icl ; 
 ebl <= icl ; 
 LAD <=  ICD & tca  |  GAD & TCA  ; 
 LAL <=  ICL & tca  |  JAB & TCA  ; 
 OAD <=  AAD & TAA  |  ICD & TAE  |  LBD & TAI  |  LAD & TAM  ; 
 OED <=  ICD & TBA  |  LAD & TBB  |  LGD & TKA  ; 
 OEL <=  ICL & TBA  |  LAL & TBB  |  LFD & TKA  ; 
 lfh <= leh ; 
 lgh <= lfh ; 
 OAL <=  AAL & TAB  |  ICL & TAF  |  LBL & TAJ  |  LAL & TAN  ; 
 OID <=  VDN  |  NBL & MAO  |  JFD & JEA  ; 
 qde <=  qdc  ; 
 bal <= idd ; 
 lbd <= lad ; 
 lcd <= lbd ; 
 ldd <= lcd ; 
 BAD <= IDD ; 
 lbl <= lal ; 
 lcl <= lbl ; 
 ldl <= lcl ; 
 OBD <=  ABD & TAC  |  LAD & TAK  |  LBD & TAO  |  TAQ  ; 
 OFD <=  LAD & TBC  |  LED & TKC  |  TBD  ; 
 OFL <=  LAL & TBC  |  IKD & TKC  |  TBD  ; 
 oua <=  gad  ; 
 ouc <=  gak  |  qad  ; 
 OBL <=  ABL & TAD  |  LAL & TAL  |  LBL & TAP  |  TAR  ; 
 old <= qla ; 
 omd <= qla ; 
 ond <= bad ; 
 qda <=  gbd  |  qaa  ; 
 qgc <=  gbl  |  qaa  ; 
 qdb <= qda ; 
 qdc <= qdb ; 
 qdd <= qdc ; 
 OCD <=  LCD & TAG  |  LAD & TAS  |  JBE & TAW  ; 
 OCL <=  LCL & TAG  |  LAL & TAS  |  JBG & TAW  ; 
 AAD <= IAD ; 
 AAL <= IAL ; 
 OGD <= IAD ; 
 OGL <= IAL ; 
 OSD <=  TXA & AAD  |  TXB & BBD  |  TXC & BDD  |  TXD & BED  ; 
 bdl <= bcd ; 
 bed <= bdl ; 
 bbd <= aal ; 
 bbl <= abd ; 
 bcd <= abl ; 
 bdd <= bbl ; 
 ODD <=  LDD & TAH  |  LBD & TAT  |  JBA & TAX  ; 
 ODL <=  LDL & TAH  |  LBL & TAT  |  JBC & TAX  ; 
 ABD <= IBD ; 
 ABL <= IBL ; 
 OHD <= IBD ; 
 OHL <= IBL ; 
 vea <=  nca  |  nbe  ; 
 VEC <=  NCC & NBE  |  VEB  ; 
 VEE <=  NCE & NBE  |  VED  ; 
 VEG <=  NCG & NBE  |  VEF  ; 
 VEH <=  NCH & NBE  |  VEG  ; 
 VED <=  NCD & NBE  |  VEC  ; 
 VEF <=  NCF & NBE  |  VEE  ; 
 VEI <=  NCI & NBE  |  VEH  ; 
 VEJ <=  NCJ & NBE  |  VEI  ; 
 NAE <= MAE ; 
 NCG <= MAG ; 
 CEA <= DEA & QOB |  BAI & qob ; 
 CEB <= DEB & QOB |  BAJ & qob ; 
 CEC <= DEC & QOB |  BAK & qob ; 
 CED <= DED & QOB |  BAL & qob ; 
 CEE <= DEE & QOB |  BAM & qob ; 
 CEF <= DEF & QOB |  BAN & qob ; 
 OKC <=  DCH & qkd & QKA  |  QTB  ; 
 NBE <= JGE ; 
 NBM <= JGE ; 
 VEB <= VEA ; 
 GAE <=  EAE & TGA  |  GAE & tga  ; 
 VEK <=  NCK & NBM  |  VEJ  ; 
 VEL <=  NCL & NBM  |  VEK  ; 
 gbe <=  faf & TGJ  |  fba & TGK  |  gbe & tgb  ; 
 VEM <=  NCM & NBM  |  VEL  ; 
 VEN <=  NCN & NBM  |  VEM  ; 
 gce <=  fap & TGF  |  TGH & fbj  |  gce & tgd  ; 
 gcm <=  fah & TGF  |  TGH & fbj  |  gcm & tgd  ; 
 MAG <=  QHD  |  QHE  ; 
 qhe <=  jcc  |  tea  ; 
 QSA <=  QSA & dfg  |  JCB & QAC  ; 
 QSB <=  QSA & dfg  |  JCB & QAC  ; 
 OKE <=  DEG & QOA  |  JDC & QAC  |  QTA  ; 
 eae <= ice ; 
 eam <= icm ; 
 ebm <= icm ; 
 ecm <= icm ; 
 LAE <=  ICE & tcb  |  GAE & TCB  ; 
 LAM <=  ICM & tcb  |  JAC & TCB  ; 
 OAE <=  AAE & THA  |  ICE & THE  |  LBE & THI  |  LAE & THM  ; 
 OEE <=  ICE & TBI  |  LAE & TBJ  |  LGE & TKB  ; 
 OEM <=  ICM & TBI  |  LAM & TBJ  |  LFE & TKB  ; 
 olf <= qsa ; 
 omf <= qsa ; 
 OAM <=  AAM & THB  |  ICM & THF  |  LBM & THJ  |  LAM & THN  ; 
 OIE <=  VEN  |  NBM & MAP  |  JFE & JEB  ; 
 bam <= ide ; 
 lbe <= lae ; 
 lce <= lbe ; 
 lde <= lce ; 
 BAE <= IDE ; 
 lbm <= lam ; 
 lcm <= lbm ; 
 ldm <= lcm ; 
 OBE <=  ABE & THC  |  LAE & THK  |  LBE & THO  |  THQ  ; 
 OFE <=  LAE & TBK  |  LEE & TKD  |  TBL  ; 
 OFM <=  LAM & TBK  |  IKE & TKD  |  TBL  ; 
 qef <= qee ; 
 qeh <= qeg ; 
 QQB <= QPF ; 
 one <= bae ; 
 OBM <=  ABM & THD  |  LAM & THL  |  LBM & THP  |  THR  ; 
 ORC <=  QPE  |  QQB  ; 
 ORD <=  QOD  ; 
 qee <=  gbe  |  qaa  ; 
 qeg <=  gbe  |  qaa  |  gaj  ; 
 oub <=  gaj  |  qad  ; 
 OCE <=  LCE & THG  |  LAE & THS  |  JBF & TAU  ; 
 OCM <=  LCM & THG  |  LAM & THS  |  JBH & TAU  ; 
 AAE <= IAE ; 
 AAM <= IAM ; 
 OGE <= IAE ; 
 OGM <= IAM ; 
 bdm <= bce ; 
 bee <= bdm ; 
 bbe <= aam ; 
 bbm <= abe ; 
 bce <= abm ; 
 bde <= bbm ; 
 OSE <=  TXE & AAE  |  TXF & BBE  |  TXG & BDE  |  TXH & BEE  ; 
 ODE <=  LDE & THH  |  LBE & THT  |  JBB & TAV  ; 
 ODM <=  LDM & THH  |  LBM & THT  |  JBD & TAV  ; 
 ABE <= IBE ; 
 ABM <= IBM ; 
 OHE <= IBE ; 
 OHM <= IBM ; 
 vfa <=  nca  |  nbf  ; 
 VFC <=  NCC & NBF  |  VFB  ; 
 VFE <=  NCE & NBF  |  VFD  ; 
 VFG <=  NCG & NBF  |  VFF  ; 
 VFH <=  NCH & NBF  |  VFG  ; 
 VFD <=  NCD & NBF  |  VFC  ; 
 VFF <=  NCF & NBF  |  VFE  ; 
 VFI <=  NCI & NBF  |  VFH  ; 
 VFJ <=  NCJ & NBF  |  VFI  ; 
 CFA <= DFA & QSB |  BAI & qsb ; 
 CFB <= DFB & QSB |  BAJ & qsb ; 
 CFC <= DFC & QSB |  BAK & qsb ; 
 CFD <= DFD & QSB |  BAL & qsb ; 
 CFE <= DFE & QSB |  BAM & qsb ; 
 CFF <= DFF & QSB |  BAN & qsb ; 
 NBF <= JGF ; 
 NBN <= JGF ; 
 VFB <= VFA ; 
 VGB <= VGA ; 
 GAF <=  EAF & TGA  |  GAF & tga  ; 
 VFK <=  NCK & NBN  |  VFJ  ; 
 VFL <=  NCL & NBN  |  VFK  ; 
 gbf <=  faf & TGJ  |  fbd & TGK  |  gbf & tgb  ; 
 gbn <=  fac & TGJ  |  fbf & TGK  |  gbn & tgb  ; 
 gdb <=  fan & TGI  |  fbh & TGL  |  gbd & tgl  ; 
 gdc <=  fan & TGI  |  fbi & TGL  |  gdc & tgl  ; 
 VFM <=  NCM & NBN  |  VFL  ; 
 VFN <=  NCN & NBN  |  VFM  ; 
 gcf <=  fap & TGF  |  fbk & TGH  |  gcf & tgd  ; 
 gcn <=  fal & TGF  |  FBK & TGH  |  gcn & tgd  ; 
 qma <= qha ; 
 qmb <= qma ; 
 qmc <= qmb ; 
 qpa <=  jda  |  qac  ; 
 qpb <=  gcp  |  gci  |  qac  ; 
 qod <= qob ; 
 QOG <= QOF ; 
 QOH <= QOG ; 
 qtc <= qta ; 
 OKF <=  DFH & qsd & QSA  |  QTA  ; 
 eaf <= icf ; 
 ean <= icn ; 
 ebn <= icn ; 
 ecn <= icn ; 
 LAF <=  ICF & tcb  |  GAF & TCB  ; 
 LAN <=  ICN & tcb  |  JAC & TCB  ; 
 OAF <=  AAF & THA  |  ICF & THE  |  LBF & THI  |  LAF & THM  ; 
 OEF <=  ICF & TBI  |  LAF & TBJ  |  LGF & TKB  ; 
 OEN <=  ICN & TBI  |  LAN & TBJ  |  LFF & TKB  ; 
 QOF <=  QOF & deg & qtc  |  JDB & QAA  ; 
 OAN <=  AAN & THB  |  ICN & THF  |  LBN & THJ  |  LAN & THN  ; 
 OIF <=  VFN  |  NBN & MAP  |  JFF & JEB  ; 
 ban <= idf ; 
 lbf <= laf ; 
 lcf <= lbf ; 
 ldf <= lcf ; 
 BAF <= IDF ; 
 lbn <= lan ; 
 ldn <= lcn ; 
 OBF <=  ABF & THC  |  LAF & THK  |  LBF & THO  |  THQ  ; 
 OFF <=  LAF & TBK  |  LEF & TKD  |  TBL  ; 
 OFN <=  LAN & TBK  |  IKF & TKD  |  TBL  ; 
 QGA <=  GBG & QAA  ; 
 QOA <=  QOA & deg  |  GCM & QAA  ; 
 QOB <=  QOA & deg  |  GCM & QAA  ; 
 OBN <=  ABN & THD  |  LAN & THL  |  LBN & THP  |  THR  ; 
 oja <= qnc ; 
 ojb <= qnd ; 
 ojl <= qnc ; 
 onf <= baf ; 
 qei <=  gbe  |  qaa  ; 
 qge <=  gbn  |  qaa  ; 
 ORA <=  QPA  ; 
 ORB <=  QPB  |  QQA  |  QOH  ; 
 OCF <=  LCF & THG  |  LAF & THS  |  JBF & TAU  ; 
 OCN <=  LCN & THG  |  LAN & THS  |  JBH & TAU  ; 
 AAF <= IAF ; 
 AAN <= IAN ; 
 OGF <= IAF ; 
 OGN <= IAN ; 
 lcn <= lbn ; 
 qej <= qei ; 
 QQA <= QPC ; 
 OSF <=  TXE & AAF  |  TXF & BBF  |  TXG & BDF  |  TXH & BEF  ; 
 bdn <= bcf ; 
 bef <= bdn ; 
 bbf <= aan ; 
 bbn <= abf ; 
 bcf <= abn ; 
 bdf <= bbn ; 
 ODF <=  LDF & THH  |  LBF & THT  |  JBB & TAV  ; 
 ODN <=  LDN & THH  |  LBN & THT  |  JBD & TAV  ; 
 ABF <= IBF ; 
 ABN <= IBN ; 
 OHF <= IBF ; 
 OHN <= IBN ; 
 vga <=  nca  |  nbg  ; 
 VGC <=  NCC & NBF  |  VGB  ; 
 VGE <=  NCE & NBF  |  VGD  ; 
 VGG <=  NCG & NBF  |  VGF  ; 
 VGH <=  NCH & NBF  |  VGG  ; 
 VGD <=  NCD & NBF  |  VGC  ; 
 VGF <=  NCF & NBF  |  VGE  ; 
 VGI <=  NCI & NBF  |  VGH  ; 
 VGJ <=  NCJ & NBF  |  VGI  ; 
 MBA <= GAG ; 
 NBG <= JGG ; 
 NBO <= JGG ; 
 GAG <=  EAG & TGA  |  GAG & tga  ; 
 VGK <=  NCK & NBN  |  VGJ  ; 
 VGL <=  NCL & NBN  |  VGK  ; 
 gbg <=  fac & TGJ  |  fbo & TGK  |  gbg & tgb  ; 
 gbo <=  fag & TGJ  |  fbb & TGK  |  gbo & tgb  ; 
 gch <=  faf & TGF  |  fbk & TGI  |  gch & tgd  ; 
 gcp <=  faf & TGF  |  fbj & TGI  |  gcp & tgd  ; 
 VGM <=  NCM & NBO  |  VGL  ; 
 VGN <=  NCN & NBO  |  VGM  ; 
 gco <=  faj & TGF  |  TGH & fbj  |  gco & tgd  ; 
 qpc <=  gch  |  gci  |  qac  ; 
 QLD <= QAC & GCK ; 
 QUA <= QAC & GDB ; 
 QVA <= QAC & GDC ; 
 eag <= icg ; 
 eao <= ico ; 
 ebo <= ico ; 
 eco <= ico ; 
 LAG <=  ICG & tcb  |  JAA & TCB  ; 
 LAO <=  ICO & tcb  |  JAC & TCB  ; 
 OAG <=  AAG & THA  |  ICG & THE  |  LBG & THI  |  LAG & THM  ; 
 OEG <=  ICG & TBI  |  LAG & TBJ  |  LGG & TKB  ; 
 OEO <=  ICO & TBI  |  LAO & TBJ  |  LFG & TKB  ; 
 OJJ <= QNF ; 
 OJK <= QNF ; 
 OAO <=  AAO & THB  |  ICO & THF  |  LBO & THJ  |  LAO & THN  ; 
 OIG <=  VGN  |  NBO & MAP  |  JFG & JEB  ; 
 lbg <= lag ; 
 lcg <= lbg ; 
 ldg <= lcg ; 
 lbo <= lao ; 
 lco <= lbo ; 
 ldo <= lco ; 
 OBG <=  ABG & THC  |  LAG & THK  |  LBG & THO  |  THQ  ; 
 OFG <=  LAG & TBK  |  LEG & TKD  |  TBL  ; 
 OFO <=  LAO & TBK  |  IKG & TKD  |  TBL  ; 
 OBO <=  ABO & THD  |  LAO & THL  |  LBO & THP  |  THR  ; 
 OJF <= QNF ; 
 OJG <= QNF ; 
 OJH <= QNF ; 
 OJI <= QNF ; 
 QBA <= IFA ; 
 QBB <= IFA ; 
 TGL <= QBB ; 
 OCG <=  LCG & THG  |  LAG & THS  |  JBF & TAU  ; 
 OCO <=  LCO & THG  |  LAO & THS  |  JBH & TAU  ; 
 AAG <= IAG ; 
 AAO <= IAO ; 
 OGG <= IAG ; 
 OGO <= IAO ; 
 OKD <=  DDH & qle & QLA  |  QLD  |  QTA  ; 
 bbg <= aao ; 
 bbo <= abg ; 
 bcg <= abo ; 
 bdg <= bbo ; 
 OSG <=  TXE & AAG  |  TXF & BBG  |  TXG & BDG  |  TXH & BEG  ; 
 bdo <= bcg ; 
 beg <= bdo ; 
 ODG <=  LDG & THH  |  LBG & THT  |  JBB & TAV  ; 
 ODO <=  LDO & THH  |  LBO & THT  |  JBD & TAV  ; 
 ABG <= IBG ; 
 ABO <= IBO ; 
 OHG <= IBG ; 
 OHO <= IBO ; 
 vha <=  nca  |  nbh  ; 
 VHC <=  NCC & NBH  |  VHB  ; 
 VHE <=  NCE & NBH  |  VHD  ; 
 VHG <=  NCG & NBH  |  VHF  ; 
 VHH <=  NCH & NBH  |  VHG  ; 
 VHD <=  NCD & NBH  |  VHC  ; 
 VHF <=  NCF & NBH  |  VHE  ; 
 VHI <=  NCI & NBH  |  VHH  ; 
 VHJ <=  NCJ & NBH  |  VHI  ; 
 MBB <= GAH ; 
 NBH <= JGH ; 
 NBP <= JGH ; 
 VHB <= VHA ; 
 GAH <=  EAH & TGA  |  GAH & tga  ; 
 VHK <=  NCK & NBH  |  VHJ  ; 
 VHL <=  NCL & NBH  |  VHK  ; 
 gbh <=  fah & TGJ  |  fbh & TGK  |  gbh & tgb  ; 
 VHM <=  NCM & NBH  |  VHL  ; 
 VHN <=  NCN & NBH  |  VHM  ; 
 qvb <= qva ; 
 qvd <= qvc ; 
 qvf <= qve ; 
 qvh <= qvg ; 
 qpe <=  gce  |  gci  |  qac  ; 
 qpf <=  gcf  |  gci  |  qac  ; 
 qvc <= qvb ; 
 qve <= qvd ; 
 qvg <= qvf ; 
 qvi <= qvh ; 
 qvj <= qvi ; 
 qvk <= qvj ; 
 txe <= quc ; 
 txf <= txa ; 
 txg <= txb ; 
 txh <= txc ; 
 eah <= ich ; 
 eap <= icp ; 
 ebp <= icp ; 
 ecp <= icp ; 
 LAH <=  ICH & tcb  |  JAA & TCB  ; 
 LAP <=  ICP & tcb  |  JAC & TCB  ; 
 OAH <=  AAH & THA  |  ICH & THE  |  LBH & THI  |  LAH & THM  ; 
 OEH <=  ICH & TBI  |  LAH & TBJ  |  LGH & TKB  ; 
 OEP <=  ICP & TBI  |  LAP & TBJ  |  LFH & TKB  ; 
 TKA <= qvk ; 
 TKB <= qvk ; 
 TKC <= qvk ; 
 TKD <= qvk ; 
 OIH <=  VHN  |  NBP & MAP  |  JFH & JEB  ; 
 OAP <=  AAP & THB  |  ICP & THF  |  LBP & THJ  |  LAP & THN  ; 
 ojc <= qne ; 
 ojd <= qnf ; 
 oje <= qnc ; 
 qce <= qcc ; 
 lbp <= lap ; 
 lcp <= lbp ; 
 ldp <= lcp ; 
 QRA <= ILA ; 
 OBH <=  ABH & THC  |  LAH & THK  |  LBH & THO  |  THQ  ; 
 OFH <=  LAH & TBK  |  LEH & TKD  |  TBL  ; 
 OFP <=  LAP & TBK  |  IKH & TKD  |  TBL  ; 
 lbh <= lah ; 
 lch <= lbh ; 
 ldh <= lch ; 
 QNB <= QNA ; 
 QND <= QNC ; 
 QNE <= QND ; 
 QNF <= QNE ; 
 OBP <=  ABP & THD  |  LAP & THL  |  LBP & THP  |  THR  ; 
 ota <=  ZZO & qnc  |  gdb & gdc  |  qad  ; 
 qna <=  iga & qnc  ; 
 qnc <=  QNC & IGA  |  QNB & qnc  |  QNA & qnc  ; 
 QAA <= IEB & IEA ; 
 QAB <= IEB & IEA ; 
 QAC <= IEB & IEA ; 
 QAD <= IEB & IEA ; 
 OCH <=  LCH & THG  |  LAH & THS  |  JBF & TAU  ; 
 OCP <=  LCP & THG  |  LAP & THS  |  JBH & TAU  ; 
 AAH <= IAH ; 
 AAP <= IAP ; 
 OGH <= IAH ; 
 OGP <= IAP ; 
 qcb <= qca ; 
 qcc <= qcb ; 
 qcd <= qcc ; 
 ODH <=  LDH & THH  |  LBH & THT  |  JBB & TAV  ; 
 ODP <=  LDP & THH  |  LBP & THT  |  JBD & TAV  ; 
 ABH <= IBH ; 
 ABP <= IBP ; 
 OHH <= IBH ; 
 OHP <= IBP ; 
 txa <= quc ; 
 txb <= txa ; 
 txc <= txb ; 
 txd <= txc ; 
 bdp <= bch ; 
 beh <= bdp ; 
 qub <= qua ; 
 quc <= qub ; 
 OSH <=  TXE & AAH  |  TXF & BBH  |  TXG & BDH  |  TXH & BEH  ; 
end
endmodule;
